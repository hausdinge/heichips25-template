VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO delay_line
  CLASS BLOCK ;
  FOREIGN delay_line ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 60.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 15.380 0.000 17.580 60.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 16.280 60.000 18.480 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 46.280 60.000 48.480 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 21.580 0.000 23.780 60.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 22.480 60.000 24.680 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 59.600 34.280 60.000 ;
    END
  END clk
  PIN clk_delayed
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.700 0.400 40.100 ;
    END
  END clk_delayed
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2.200 0.000 2.600 0.400 ;
    END
  END reset
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 28.120 59.600 28.520 60.000 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.140 0.400 32.540 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.300 0.400 31.700 ;
    END
  END sel[2]
  PIN trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 34.840 59.600 35.240 60.000 ;
    END
  END trim[0]
  PIN trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.600 23.740 60.000 24.140 ;
    END
  END trim[1]
  PIN trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END trim[2]
  PIN trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.860 0.400 18.260 ;
    END
  END trim[3]
  PIN trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 36.760 59.600 37.160 60.000 ;
    END
  END trim[4]
  PIN trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.600 33.820 60.000 34.220 ;
    END
  END trim[5]
  PIN trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 35.800 0.000 36.200 0.400 ;
    END
  END trim[6]
  PIN trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 12.760 0.000 13.160 0.400 ;
    END
  END trim[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 57.120 53.070 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 57.120 53.140 ;
      LAYER Metal2 ;
        RECT 3.255 59.390 27.910 59.600 ;
        RECT 28.730 59.390 33.670 59.600 ;
        RECT 34.490 59.390 34.630 59.600 ;
        RECT 35.450 59.390 36.550 59.600 ;
        RECT 37.370 59.390 58.185 59.600 ;
        RECT 3.255 0.610 58.185 59.390 ;
        RECT 3.255 0.100 12.550 0.610 ;
        RECT 13.370 0.100 25.030 0.610 ;
        RECT 25.850 0.100 35.590 0.610 ;
        RECT 36.410 0.100 58.185 0.610 ;
      LAYER Metal3 ;
        RECT 0.400 40.310 59.600 56.380 ;
        RECT 0.610 39.490 59.600 40.310 ;
        RECT 0.400 34.430 59.600 39.490 ;
        RECT 0.400 33.610 59.390 34.430 ;
        RECT 0.400 32.750 59.600 33.610 ;
        RECT 0.610 31.930 59.600 32.750 ;
        RECT 0.400 31.910 59.600 31.930 ;
        RECT 0.610 31.090 59.600 31.910 ;
        RECT 0.400 24.350 59.600 31.090 ;
        RECT 0.400 23.530 59.390 24.350 ;
        RECT 0.400 18.470 59.600 23.530 ;
        RECT 0.610 17.650 59.600 18.470 ;
        RECT 0.400 0.320 59.600 17.650 ;
      LAYER Metal4 ;
        RECT 14.295 42.690 15.170 50.965 ;
        RECT 17.790 42.690 21.370 50.965 ;
        RECT 23.990 42.690 51.465 50.965 ;
      LAYER Metal5 ;
        RECT 14.255 43.160 51.505 43.360 ;
  END
END delay_line
END LIBRARY

