* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for delay_line abstract view
.subckt delay_line VDD VSS clk clk_delayed delay[0] delay[1] delay[2] delay[3]
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for adc abstract view
.subckt adc VDD VSS analog_in[0] analog_in[1] analog_in[2] analog_in[3] analog_in[4]
+ analog_in[5] analog_in[6] analog_in[7] clk data_out[0] data_out[1] data_out[2] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] ready start
.ends

* Black-box entry subcircuit for multimode_dll abstract view
.subckt multimode_dll VDD VSS bias clk0_out clk0_phase_sel[0] clk0_phase_sel[1] clk0_phase_sel[2]
+ clk0_phase_sel[3] clk0_phase_sel[4] clk1_out clk1_phase_sel[0] clk1_phase_sel[1]
+ clk1_phase_sel[2] clk1_phase_sel[3] clk1_phase_sel[4] clk2_out clk2_phase_sel[0]
+ clk2_phase_sel[1] clk2_phase_sel[2] clk2_phase_sel[3] clk2_phase_sel[4] dco enable
+ ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14] ext_trim[15]
+ ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20] ext_trim[21]
+ ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3] ext_trim[4]
+ ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] f_clk0_divider[0] f_clk0_divider[1]
+ f_clk0_divider[2] f_clk0_divider[3] f_clk0_divider[4] f_clk1_divider[0] f_clk1_divider[1]
+ f_clk1_divider[2] f_clk1_divider[3] f_clk1_divider[4] f_clk2_divider[0] f_clk2_divider[1]
+ f_clk2_divider[2] f_clk2_divider[3] f_clk2_divider[4] f_osc_multiply_factor[0] f_osc_multiply_factor[1]
+ f_osc_multiply_factor[2] f_osc_multiply_factor[3] f_osc_multiply_factor[4] mode_xor[0]
+ mode_xor[1] mode_xor[2] osc osc_out resetb stable
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_11_807 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_27_940 VPWR VGND sg13g2_decap_8
XFILLER_46_759 VPWR VGND sg13g2_decap_8
XFILLER_45_203 VPWR VGND sg13g2_decap_8
X_294_ net29 VGND VPWR _054_ data\[47\] clknet_4_3_0_clk_regs sg13g2_dfrbpq_1
XFILLER_6_800 VPWR VGND sg13g2_decap_8
XFILLER_42_95 VPWR VGND sg13g2_fill_1
XFILLER_49_564 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_decap_8
XFILLER_45_792 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_46_556 VPWR VGND sg13g2_decap_8
XFILLER_42_740 VPWR VGND sg13g2_decap_8
X_277_ net30 VGND VPWR _037_ data\[30\] clknet_4_2_0_clk_regs sg13g2_dfrbpq_1
XFILLER_38_4 VPWR VGND sg13g2_fill_1
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_0_839 VPWR VGND sg13g2_decap_8
XFILLER_43_559 VPWR VGND sg13g2_decap_8
X_200_ data\[39\] data\[40\] net17 _047_ VPWR VGND sg13g2_mux2_1
X_131_ clk_delayed net5 _095_ VPWR VGND net4 sg13g2_nand3b_1
XFILLER_2_165 VPWR VGND sg13g2_decap_4
XFILLER_3_655 VPWR VGND sg13g2_decap_8
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_46_353 VPWR VGND sg13g2_decap_8
XFILLER_30_765 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_38_821 VPWR VGND sg13g2_decap_8
XFILLER_0_636 VPWR VGND sg13g2_decap_8
XFILLER_29_821 VPWR VGND sg13g2_decap_8
XFILLER_12_765 VPWR VGND sg13g2_decap_8
XFILLER_3_430 VPWR VGND sg13g2_fill_2
XFILLER_3_496 VPWR VGND sg13g2_fill_2
XFILLER_47_651 VPWR VGND sg13g2_decap_8
XFILLER_46_150 VPWR VGND sg13g2_decap_8
XFILLER_26_835 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_29_52 VPWR VGND sg13g2_decap_4
XFILLER_32_849 VPWR VGND sg13g2_decap_8
XFILLER_44_665 VPWR VGND sg13g2_decap_8
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_43_186 VPWR VGND sg13g2_decap_8
XFILLER_4_772 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_fill_2
XFILLER_2_709 VPWR VGND sg13g2_decap_8
Xheichips25_template_43 VPWR VGND uio_oe[1] sg13g2_tielo
Xheichips25_template_54 VPWR VGND uo_out[4] sg13g2_tielo
Xoutput7 net7 uio_out[1] VPWR VGND sg13g2_buf_1
XFILLER_49_746 VPWR VGND sg13g2_decap_8
XFILLER_0_263 VPWR VGND sg13g2_decap_8
XFILLER_1_797 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_44_484 VPWR VGND sg13g2_decap_8
XFILLER_9_842 VPWR VGND sg13g2_decap_4
XFILLER_46_738 VPWR VGND sg13g2_decap_8
XFILLER_27_996 VPWR VGND sg13g2_decap_8
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_6_845 VPWR VGND sg13g2_fill_2
X_293_ net31 VGND VPWR _053_ data\[46\] clknet_4_1_0_clk_regs sg13g2_dfrbpq_1
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_1_583 VPWR VGND sg13g2_decap_8
XFILLER_45_771 VPWR VGND sg13g2_decap_8
XFILLER_49_543 VPWR VGND sg13g2_decap_8
XFILLER_44_292 VPWR VGND sg13g2_fill_2
XFILLER_36_793 VPWR VGND sg13g2_decap_8
XFILLER_3_837 VPWR VGND sg13g2_decap_8
XFILLER_46_535 VPWR VGND sg13g2_decap_8
XFILLER_42_796 VPWR VGND sg13g2_decap_8
XFILLER_27_793 VPWR VGND sg13g2_decap_8
X_276_ net34 VGND VPWR _036_ data\[29\] clknet_4_9_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_340 VPWR VGND sg13g2_decap_8
XFILLER_18_793 VPWR VGND sg13g2_decap_8
XFILLER_0_818 VPWR VGND sg13g2_decap_4
X_130_ VPWR net12 _094_ VGND sg13g2_inv_1
XFILLER_3_634 VPWR VGND sg13g2_decap_8
XFILLER_47_833 VPWR VGND sg13g2_decap_8
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_46_332 VPWR VGND sg13g2_decap_8
XFILLER_42_582 VPWR VGND sg13g2_decap_8
X_259_ net37 VGND VPWR _019_ data\[12\] clknet_4_7_0_clk_regs sg13g2_dfrbpq_1
XFILLER_38_800 VPWR VGND sg13g2_decap_8
XFILLER_29_800 VPWR VGND sg13g2_decap_8
XFILLER_0_615 VPWR VGND sg13g2_decap_8
XFILLER_35_814 VPWR VGND sg13g2_decap_8
XFILLER_47_630 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_26_814 VPWR VGND sg13g2_decap_8
XFILLER_41_828 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_32_828 VPWR VGND sg13g2_decap_8
XFILLER_44_644 VPWR VGND sg13g2_decap_8
XFILLER_17_847 VPWR VGND sg13g2_fill_1
XFILLER_25_880 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_8
XFILLER_23_828 VPWR VGND sg13g2_decap_8
Xheichips25_template_44 VPWR VGND uio_oe[2] sg13g2_tielo
Xheichips25_template_55 VPWR VGND uo_out[5] sg13g2_tielo
XFILLER_15_55 VPWR VGND sg13g2_fill_1
XFILLER_15_44 VPWR VGND sg13g2_decap_8
XFILLER_49_725 VPWR VGND sg13g2_decap_8
Xoutput10 net10 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput8 net8 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_776 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_9_821 VPWR VGND sg13g2_decap_8
XFILLER_48_791 VPWR VGND sg13g2_decap_8
XFILLER_2_507 VPWR VGND sg13g2_fill_2
XFILLER_46_717 VPWR VGND sg13g2_decap_8
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_27_975 VPWR VGND sg13g2_decap_8
XFILLER_42_42 VPWR VGND sg13g2_decap_8
X_292_ net33 VGND VPWR _052_ data\[45\] clknet_4_6_0_clk_regs sg13g2_dfrbpq_1
XFILLER_10_842 VPWR VGND sg13g2_decap_4
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_45_750 VPWR VGND sg13g2_decap_8
XFILLER_49_599 VPWR VGND sg13g2_decap_8
XFILLER_44_271 VPWR VGND sg13g2_decap_8
XFILLER_36_772 VPWR VGND sg13g2_decap_8
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_27_772 VPWR VGND sg13g2_decap_8
XFILLER_46_514 VPWR VGND sg13g2_decap_8
XFILLER_37_20 VPWR VGND sg13g2_fill_1
XFILLER_42_775 VPWR VGND sg13g2_decap_8
X_275_ net34 VGND VPWR _035_ data\[28\] clknet_4_9_0_clk_regs sg13g2_dfrbpq_1
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_33_786 VPWR VGND sg13g2_decap_8
XFILLER_18_772 VPWR VGND sg13g2_decap_8
XFILLER_24_786 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_3_613 VPWR VGND sg13g2_decap_8
XFILLER_47_812 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_46_311 VPWR VGND sg13g2_decap_8
XFILLER_42_561 VPWR VGND sg13g2_decap_8
XFILLER_15_786 VPWR VGND sg13g2_decap_8
XFILLER_15_797 VPWR VGND sg13g2_fill_1
XFILLER_46_388 VPWR VGND sg13g2_decap_8
X_189_ data\[28\] data\[29\] net19 _036_ VPWR VGND sg13g2_mux2_1
X_258_ net36 VGND VPWR _018_ data\[11\] clknet_4_7_0_clk_regs sg13g2_dfrbpq_1
XFILLER_38_856 VPWR VGND sg13g2_decap_4
Xclkbuf_4_9_0_clk_regs clknet_0_clk_regs clknet_4_9_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_49_193 VPWR VGND sg13g2_decap_8
XFILLER_29_856 VPWR VGND sg13g2_decap_4
XFILLER_48_609 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_44_826 VPWR VGND sg13g2_decap_8
XFILLER_43_303 VPWR VGND sg13g2_decap_4
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_3_432 VPWR VGND sg13g2_fill_1
XFILLER_3_498 VPWR VGND sg13g2_fill_1
XFILLER_47_686 VPWR VGND sg13g2_decap_8
XFILLER_46_185 VPWR VGND sg13g2_decap_8
XFILLER_7_793 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_4
XFILLER_41_807 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_0_402 VPWR VGND sg13g2_fill_2
XFILLER_44_623 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_0_479 VPWR VGND sg13g2_fill_2
XFILLER_17_826 VPWR VGND sg13g2_decap_8
XFILLER_40_851 VPWR VGND sg13g2_decap_8
XFILLER_32_807 VPWR VGND sg13g2_decap_8
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_43_133 VPWR VGND sg13g2_decap_4
XFILLER_43_166 VPWR VGND sg13g2_fill_2
XFILLER_6_25 VPWR VGND sg13g2_decap_4
XFILLER_3_284 VPWR VGND sg13g2_decap_4
XFILLER_23_807 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
Xheichips25_template_45 VPWR VGND uio_oe[3] sg13g2_tielo
Xheichips25_template_56 VPWR VGND uo_out[6] sg13g2_tielo
XFILLER_14_807 VPWR VGND sg13g2_decap_8
XFILLER_31_55 VPWR VGND sg13g2_fill_1
XFILLER_49_704 VPWR VGND sg13g2_decap_8
XFILLER_0_221 VPWR VGND sg13g2_decap_8
Xoutput11 net11 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_0_298 VPWR VGND sg13g2_fill_1
XFILLER_44_464 VPWR VGND sg13g2_fill_2
XFILLER_9_800 VPWR VGND sg13g2_decap_8
XFILLER_48_770 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_decap_8
XFILLER_27_954 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_10_821 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_42_76 VPWR VGND sg13g2_decap_8
X_291_ net33 VGND VPWR _051_ data\[44\] clknet_4_6_0_clk_regs sg13g2_dfrbpq_1
Xclkbuf_4_11_0_clk_regs clknet_0_clk_regs clknet_4_11_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_6_814 VPWR VGND sg13g2_decap_8
XFILLER_6_847 VPWR VGND sg13g2_fill_1
XFILLER_49_578 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_44_250 VPWR VGND sg13g2_decap_8
XFILLER_44_294 VPWR VGND sg13g2_fill_1
XFILLER_42_209 VPWR VGND sg13g2_decap_4
XFILLER_42_754 VPWR VGND sg13g2_decap_8
X_274_ net34 VGND VPWR _034_ data\[27\] clknet_4_8_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_33_765 VPWR VGND sg13g2_decap_8
XFILLER_24_765 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_3_669 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_46_367 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_decap_4
XFILLER_15_765 VPWR VGND sg13g2_decap_8
X_326_ net32 VGND VPWR _086_ u_shift_reg.locked clknet_4_1_0_clk_regs sg13g2_dfrbpq_1
XFILLER_30_779 VPWR VGND sg13g2_decap_8
X_188_ data\[27\] data\[28\] net19 _035_ VPWR VGND sg13g2_mux2_1
X_257_ net36 VGND VPWR _017_ data\[10\] clknet_4_11_0_clk_regs sg13g2_dfrbpq_1
XFILLER_38_835 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_44_805 VPWR VGND sg13g2_decap_8
XFILLER_29_835 VPWR VGND sg13g2_decap_8
XFILLER_34_44 VPWR VGND sg13g2_decap_8
XFILLER_34_55 VPWR VGND sg13g2_fill_1
XFILLER_12_779 VPWR VGND sg13g2_decap_8
XFILLER_3_466 VPWR VGND sg13g2_decap_4
XFILLER_47_665 VPWR VGND sg13g2_decap_8
XFILLER_46_164 VPWR VGND sg13g2_decap_8
XFILLER_43_860 VPWR VGND sg13g2_fill_2
X_309_ net28 VGND VPWR _069_ data\[62\] clknet_4_3_0_clk_regs sg13g2_dfrbpq_1
XFILLER_7_772 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_26_849 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_20_24 VPWR VGND sg13g2_decap_4
XFILLER_44_602 VPWR VGND sg13g2_decap_8
XFILLER_17_805 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_44_679 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_3_263 VPWR VGND sg13g2_decap_8
XFILLER_4_786 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
Xheichips25_template_46 VPWR VGND uio_oe[4] sg13g2_tielo
Xheichips25_template_57 VPWR VGND uo_out[7] sg13g2_tielo
Xoutput12 net12 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_277 VPWR VGND sg13g2_decap_8
XFILLER_1_723 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_44_443 VPWR VGND sg13g2_decap_8
XFILLER_44_498 VPWR VGND sg13g2_decap_8
XFILLER_2_509 VPWR VGND sg13g2_fill_1
XFILLER_27_933 VPWR VGND sg13g2_decap_8
XFILLER_39_793 VPWR VGND sg13g2_decap_8
XFILLER_10_800 VPWR VGND sg13g2_decap_8
X_290_ net33 VGND VPWR _050_ data\[43\] clknet_4_5_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_1_597 VPWR VGND sg13g2_decap_8
XFILLER_45_785 VPWR VGND sg13g2_decap_8
XFILLER_46_549 VPWR VGND sg13g2_decap_8
XFILLER_42_733 VPWR VGND sg13g2_decap_8
XFILLER_42_711 VPWR VGND sg13g2_fill_2
XFILLER_42_700 VPWR VGND sg13g2_decap_8
X_273_ net35 VGND VPWR _033_ data\[26\] clknet_4_8_0_clk_regs sg13g2_dfrbpq_1
XFILLER_1_383 VPWR VGND sg13g2_fill_2
XFILLER_45_582 VPWR VGND sg13g2_decap_8
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_2_158 VPWR VGND sg13g2_decap_8
XFILLER_3_648 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_46_346 VPWR VGND sg13g2_decap_8
X_325_ net41 VGND VPWR _085_ data\[78\] clknet_4_15_0_clk_regs sg13g2_dfrbpq_1
XFILLER_42_596 VPWR VGND sg13g2_decap_8
X_187_ data\[26\] data\[27\] net19 _034_ VPWR VGND sg13g2_mux2_1
X_256_ net39 VGND VPWR _016_ data\[9\] clknet_4_10_0_clk_regs sg13g2_dfrbpq_1
XFILLER_38_814 VPWR VGND sg13g2_decap_8
XFILLER_2_681 VPWR VGND sg13g2_decap_8
XFILLER_49_151 VPWR VGND sg13g2_decap_8
XFILLER_0_629 VPWR VGND sg13g2_decap_8
Xu_delay_line VPWR VGND clknet_1_1__leaf_clk clk_delayed data\[75\] data\[76\] data\[77\]
+ data\[78\] delay_line
XFILLER_29_814 VPWR VGND sg13g2_decap_8
XFILLER_34_23 VPWR VGND sg13g2_decap_4
XFILLER_3_423 VPWR VGND sg13g2_decap_8
Xclkload0 VPWR clkload0/Y clknet_4_1_0_clk_regs VGND sg13g2_inv_1
XFILLER_3_489 VPWR VGND sg13g2_decap_8
XFILLER_35_828 VPWR VGND sg13g2_decap_8
XFILLER_47_644 VPWR VGND sg13g2_decap_8
XFILLER_46_143 VPWR VGND sg13g2_decap_8
X_308_ net29 VGND VPWR _068_ data\[61\] clknet_4_2_0_clk_regs sg13g2_dfrbpq_1
X_239_ _103_ net2 u_shift_reg.locked _086_ VPWR VGND sg13g2_a21o_1
XFILLER_26_828 VPWR VGND sg13g2_decap_8
XFILLER_0_404 VPWR VGND sg13g2_fill_1
XFILLER_29_34 VPWR VGND sg13g2_fill_2
XFILLER_29_45 VPWR VGND sg13g2_decap_8
XFILLER_44_658 VPWR VGND sg13g2_decap_8
XFILLER_45_77 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_fill_1
XFILLER_25_894 VPWR VGND sg13g2_decap_8
XFILLER_43_179 VPWR VGND sg13g2_decap_8
XFILLER_4_765 VPWR VGND sg13g2_decap_8
XFILLER_47_441 VPWR VGND sg13g2_decap_8
Xheichips25_template_47 VPWR VGND uio_oe[5] sg13g2_tielo
XFILLER_22_842 VPWR VGND sg13g2_decap_4
Xoutput13 net13 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_702 VPWR VGND sg13g2_decap_8
XFILLER_49_739 VPWR VGND sg13g2_decap_8
XFILLER_0_256 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_13_842 VPWR VGND sg13g2_decap_4
XFILLER_44_422 VPWR VGND sg13g2_decap_8
XFILLER_44_477 VPWR VGND sg13g2_decap_8
XFILLER_9_846 VPWR VGND sg13g2_fill_2
XFILLER_9_835 VPWR VGND sg13g2_decap_8
XFILLER_0_790 VPWR VGND sg13g2_decap_8
XFILLER_27_912 VPWR VGND sg13g2_decap_8
XFILLER_39_772 VPWR VGND sg13g2_decap_8
XFILLER_27_989 VPWR VGND sg13g2_decap_8
XFILLER_6_838 VPWR VGND sg13g2_decap_8
XFILLER_27_1010 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_1_576 VPWR VGND sg13g2_decap_8
XFILLER_45_764 VPWR VGND sg13g2_decap_8
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_44_285 VPWR VGND sg13g2_decap_8
XFILLER_36_786 VPWR VGND sg13g2_decap_8
XFILLER_46_528 VPWR VGND sg13g2_decap_8
XFILLER_42_789 VPWR VGND sg13g2_decap_8
XFILLER_27_786 VPWR VGND sg13g2_decap_8
X_272_ net35 VGND VPWR _032_ data\[25\] clknet_4_8_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_45_561 VPWR VGND sg13g2_decap_8
XFILLER_18_786 VPWR VGND sg13g2_decap_8
XFILLER_3_627 VPWR VGND sg13g2_decap_8
XFILLER_2_137 VPWR VGND sg13g2_decap_8
XFILLER_47_826 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_46_325 VPWR VGND sg13g2_decap_8
X_324_ net41 VGND VPWR _084_ data\[77\] clknet_4_15_0_clk_regs sg13g2_dfrbpq_1
XFILLER_42_575 VPWR VGND sg13g2_decap_8
X_255_ net39 VGND VPWR _015_ data\[8\] clknet_4_11_0_clk_regs sg13g2_dfrbpq_1
X_186_ data\[25\] data\[26\] net20 _033_ VPWR VGND sg13g2_mux2_1
XFILLER_2_660 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_49_130 VPWR VGND sg13g2_decap_8
XFILLER_0_608 VPWR VGND sg13g2_decap_8
XFILLER_34_13 VPWR VGND sg13g2_decap_4
Xclkload1 VPWR clkload1/Y clknet_4_3_0_clk_regs VGND sg13g2_inv_1
XFILLER_47_623 VPWR VGND sg13g2_decap_8
XFILLER_35_807 VPWR VGND sg13g2_decap_8
XFILLER_46_199 VPWR VGND sg13g2_decap_8
X_238_ data\[77\] data\[78\] net27 _085_ VPWR VGND sg13g2_mux2_1
X_307_ net30 VGND VPWR _067_ data\[60\] clknet_4_2_0_clk_regs sg13g2_dfrbpq_1
X_169_ data\[8\] data\[9\] net25 _016_ VPWR VGND sg13g2_mux2_1
XFILLER_26_807 VPWR VGND sg13g2_decap_8
XFILLER_34_851 VPWR VGND sg13g2_decap_8
XFILLER_0_449 VPWR VGND sg13g2_decap_4
XFILLER_40_821 VPWR VGND sg13g2_decap_8
XFILLER_44_637 VPWR VGND sg13g2_decap_8
XFILLER_25_873 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
Xclkbuf_4_8_0_clk_regs clknet_0_clk_regs clknet_4_8_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_3_298 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_31_821 VPWR VGND sg13g2_fill_2
XFILLER_43_692 VPWR VGND sg13g2_decap_8
Xheichips25_template_48 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_22_821 VPWR VGND sg13g2_decap_8
XFILLER_31_25 VPWR VGND sg13g2_fill_1
XFILLER_1_769 VPWR VGND sg13g2_decap_8
XFILLER_49_718 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_44_401 VPWR VGND sg13g2_decap_8
XFILLER_9_814 VPWR VGND sg13g2_decap_8
XFILLER_13_821 VPWR VGND sg13g2_decap_4
XFILLER_48_784 VPWR VGND sg13g2_decap_8
XFILLER_47_294 VPWR VGND sg13g2_decap_8
XFILLER_27_968 VPWR VGND sg13g2_decap_8
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_10_846 VPWR VGND sg13g2_fill_2
XFILLER_10_835 VPWR VGND sg13g2_decap_8
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_45_743 VPWR VGND sg13g2_decap_8
XFILLER_44_264 VPWR VGND sg13g2_decap_8
XFILLER_48_581 VPWR VGND sg13g2_decap_8
XFILLER_36_765 VPWR VGND sg13g2_decap_8
XFILLER_3_809 VPWR VGND sg13g2_decap_8
XFILLER_27_765 VPWR VGND sg13g2_decap_8
XFILLER_46_507 VPWR VGND sg13g2_decap_8
XFILLER_42_768 VPWR VGND sg13g2_decap_8
X_271_ net35 VGND VPWR _031_ data\[24\] clknet_4_10_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_fill_1
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_33_779 VPWR VGND sg13g2_decap_8
XFILLER_45_540 VPWR VGND sg13g2_decap_8
XFILLER_18_765 VPWR VGND sg13g2_decap_8
Xclkbuf_4_10_0_clk_regs clknet_0_clk_regs clknet_4_10_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_24_779 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_3_606 VPWR VGND sg13g2_decap_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_46_304 VPWR VGND sg13g2_decap_8
XFILLER_15_779 VPWR VGND sg13g2_decap_8
X_323_ net41 VGND VPWR _083_ data\[76\] clknet_4_15_0_clk_regs sg13g2_dfrbpq_1
X_254_ net39 VGND VPWR _014_ data\[7\] clknet_4_11_0_clk_regs sg13g2_dfrbpq_1
X_185_ data\[24\] data\[25\] net20 _032_ VPWR VGND sg13g2_mux2_1
XFILLER_38_849 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_4
XFILLER_49_186 VPWR VGND sg13g2_decap_8
XFILLER_44_819 VPWR VGND sg13g2_decap_8
XFILLER_37_860 VPWR VGND sg13g2_fill_2
XFILLER_29_849 VPWR VGND sg13g2_decap_8
XFILLER_20_793 VPWR VGND sg13g2_decap_8
Xclkload2 VPWR clkload2/Y clknet_4_5_0_clk_regs VGND sg13g2_inv_1
XFILLER_28_860 VPWR VGND sg13g2_fill_2
XFILLER_47_679 VPWR VGND sg13g2_decap_8
XFILLER_47_602 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
X_306_ net30 VGND VPWR _066_ data\[59\] clknet_4_2_0_clk_regs sg13g2_dfrbpq_1
XFILLER_46_178 VPWR VGND sg13g2_decap_8
X_237_ data\[76\] data\[77\] net27 _084_ VPWR VGND sg13g2_mux2_1
XFILLER_7_786 VPWR VGND sg13g2_decap_8
XFILLER_11_793 VPWR VGND sg13g2_decap_8
X_168_ data\[7\] data\[8\] net25 _015_ VPWR VGND sg13g2_mux2_1
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_17_819 VPWR VGND sg13g2_decap_8
XFILLER_29_36 VPWR VGND sg13g2_fill_1
XFILLER_40_800 VPWR VGND sg13g2_decap_8
XFILLER_44_616 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_43_137 VPWR VGND sg13g2_fill_2
XFILLER_3_200 VPWR VGND sg13g2_fill_2
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_3_277 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_31_855 VPWR VGND sg13g2_decap_8
XFILLER_31_800 VPWR VGND sg13g2_decap_8
XFILLER_43_671 VPWR VGND sg13g2_decap_8
XFILLER_42_170 VPWR VGND sg13g2_fill_2
Xheichips25_template_49 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_22_800 VPWR VGND sg13g2_decap_8
XFILLER_31_48 VPWR VGND sg13g2_decap_8
XFILLER_0_214 VPWR VGND sg13g2_decap_8
XFILLER_1_737 VPWR VGND sg13g2_decap_8
XFILLER_44_457 VPWR VGND sg13g2_decap_8
XFILLER_13_800 VPWR VGND sg13g2_decap_8
XFILLER_48_763 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_27_947 VPWR VGND sg13g2_decap_8
XFILLER_10_814 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_6_807 VPWR VGND sg13g2_decap_8
XFILLER_45_799 VPWR VGND sg13g2_decap_8
XFILLER_45_722 VPWR VGND sg13g2_decap_8
XFILLER_44_243 VPWR VGND sg13g2_decap_8
XFILLER_48_560 VPWR VGND sg13g2_decap_8
XFILLER_42_747 VPWR VGND sg13g2_decap_8
X_270_ net35 VGND VPWR _030_ data\[23\] clknet_4_10_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_45_596 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_8
X_322_ net41 VGND VPWR _082_ data\[75\] clknet_4_15_0_clk_regs sg13g2_dfrbpq_1
X_253_ net39 VGND VPWR _013_ data\[6\] clknet_4_11_0_clk_regs sg13g2_dfrbpq_1
X_184_ data\[23\] data\[24\] net20 _031_ VPWR VGND sg13g2_mux2_1
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_2_695 VPWR VGND sg13g2_decap_8
XFILLER_46_861 VPWR VGND sg13g2_fill_1
XFILLER_46_850 VPWR VGND sg13g2_decap_8
XFILLER_38_828 VPWR VGND sg13g2_decap_8
XFILLER_49_165 VPWR VGND sg13g2_decap_8
XFILLER_45_382 VPWR VGND sg13g2_decap_8
XFILLER_29_828 VPWR VGND sg13g2_decap_8
XFILLER_20_772 VPWR VGND sg13g2_decap_8
Xclkload3 VPWR clkload3/Y clknet_4_7_0_clk_regs VGND sg13g2_inv_1
XFILLER_47_658 VPWR VGND sg13g2_decap_8
XFILLER_46_157 VPWR VGND sg13g2_decap_8
XFILLER_43_853 VPWR VGND sg13g2_decap_8
X_305_ net36 VGND VPWR _065_ data\[58\] clknet_4_6_0_clk_regs sg13g2_dfrbpq_1
X_236_ data\[75\] data\[76\] net27 _083_ VPWR VGND sg13g2_mux2_1
X_167_ data\[6\] data\[7\] net25 _014_ VPWR VGND sg13g2_mux2_1
XFILLER_7_765 VPWR VGND sg13g2_decap_8
XFILLER_11_772 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_20_28 VPWR VGND sg13g2_fill_1
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_3_212 VPWR VGND sg13g2_fill_2
XFILLER_3_256 VPWR VGND sg13g2_decap_8
XFILLER_10_50 VPWR VGND sg13g2_decap_4
XFILLER_4_779 VPWR VGND sg13g2_decap_8
XFILLER_43_650 VPWR VGND sg13g2_decap_8
XFILLER_16_820 VPWR VGND sg13g2_fill_1
XFILLER_47_455 VPWR VGND sg13g2_decap_8
X_219_ data\[58\] data\[59\] net16 _066_ VPWR VGND sg13g2_mux2_1
XFILLER_18_0 VPWR VGND sg13g2_fill_2
XFILLER_1_716 VPWR VGND sg13g2_decap_8
XFILLER_44_436 VPWR VGND sg13g2_decap_8
XFILLER_48_742 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clknet_0_clk delaynet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_27_926 VPWR VGND sg13g2_decap_8
XFILLER_39_786 VPWR VGND sg13g2_decap_8
XFILLER_26_49 VPWR VGND sg13g2_decap_8
XFILLER_27_1024 VPWR VGND sg13g2_decap_4
XFILLER_45_701 VPWR VGND sg13g2_decap_8
XFILLER_45_778 VPWR VGND sg13g2_decap_8
XFILLER_42_726 VPWR VGND sg13g2_decap_8
XFILLER_2_800 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_45_575 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_46_339 VPWR VGND sg13g2_decap_8
XFILLER_42_589 VPWR VGND sg13g2_decap_8
Xfanout40 net41 net40 VPWR VGND sg13g2_buf_1
X_321_ net41 VGND VPWR _081_ data\[74\] clknet_4_15_0_clk_regs sg13g2_dfrbpq_1
X_252_ net39 VGND VPWR _012_ data\[5\] clknet_4_11_0_clk_regs sg13g2_dfrbpq_1
X_183_ data\[22\] data\[23\] net20 _030_ VPWR VGND sg13g2_mux2_1
XFILLER_38_807 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_2_674 VPWR VGND sg13g2_decap_8
XFILLER_49_144 VPWR VGND sg13g2_decap_8
XFILLER_45_361 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_29_807 VPWR VGND sg13g2_decap_8
Xclkload4 VPWR clkload4/Y clknet_4_9_0_clk_regs VGND sg13g2_inv_1
XFILLER_3_416 VPWR VGND sg13g2_decap_8
XFILLER_43_832 VPWR VGND sg13g2_decap_8
XFILLER_47_637 VPWR VGND sg13g2_decap_8
XFILLER_46_136 VPWR VGND sg13g2_decap_8
X_235_ data\[74\] data\[75\] net27 _082_ VPWR VGND sg13g2_mux2_1
X_304_ net36 VGND VPWR _064_ data\[57\] clknet_4_6_0_clk_regs sg13g2_dfrbpq_1
X_166_ data\[5\] data\[6\] net25 _013_ VPWR VGND sg13g2_mux2_1
XFILLER_41_7 VPWR VGND sg13g2_decap_4
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_2_471 VPWR VGND sg13g2_decap_8
XFILLER_34_821 VPWR VGND sg13g2_decap_8
XFILLER_29_27 VPWR VGND sg13g2_decap_8
XFILLER_25_821 VPWR VGND sg13g2_decap_8
XFILLER_40_835 VPWR VGND sg13g2_decap_4
XFILLER_25_887 VPWR VGND sg13g2_decap_8
Xclkbuf_regs_0_clk clk_regs clk VPWR VGND sg13g2_buf_16
XFILLER_47_434 VPWR VGND sg13g2_decap_8
X_149_ VPWR _002_ _109_ VGND sg13g2_inv_1
X_218_ data\[57\] data\[58\] net21 _065_ VPWR VGND sg13g2_mux2_1
XFILLER_22_846 VPWR VGND sg13g2_fill_2
XFILLER_22_835 VPWR VGND sg13g2_decap_8
XFILLER_13_835 VPWR VGND sg13g2_decap_8
XFILLER_44_415 VPWR VGND sg13g2_decap_8
XFILLER_9_828 VPWR VGND sg13g2_decap_8
XFILLER_13_846 VPWR VGND sg13g2_fill_2
XFILLER_48_798 VPWR VGND sg13g2_decap_8
XFILLER_48_721 VPWR VGND sg13g2_decap_8
XFILLER_0_783 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_30_0 VPWR VGND sg13g2_fill_2
XFILLER_27_905 VPWR VGND sg13g2_decap_8
XFILLER_39_765 VPWR VGND sg13g2_decap_8
Xclkbuf_4_7_0_clk_regs clknet_0_clk_regs clknet_4_7_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_27_1003 VPWR VGND sg13g2_decap_8
XFILLER_1_569 VPWR VGND sg13g2_decap_8
XFILLER_49_529 VPWR VGND sg13g2_decap_8
XFILLER_26_982 VPWR VGND sg13g2_decap_8
XFILLER_45_757 VPWR VGND sg13g2_decap_8
XFILLER_44_278 VPWR VGND sg13g2_decap_8
XFILLER_5_842 VPWR VGND sg13g2_decap_4
XFILLER_0_580 VPWR VGND sg13g2_decap_8
XFILLER_36_779 VPWR VGND sg13g2_decap_8
XFILLER_48_595 VPWR VGND sg13g2_decap_8
XFILLER_37_27 VPWR VGND sg13g2_fill_1
XFILLER_37_38 VPWR VGND sg13g2_fill_2
XFILLER_27_779 VPWR VGND sg13g2_decap_8
XFILLER_1_355 VPWR VGND sg13g2_fill_1
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_45_554 VPWR VGND sg13g2_decap_8
XFILLER_18_779 VPWR VGND sg13g2_decap_8
XFILLER_41_793 VPWR VGND sg13g2_decap_8
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_4_53 VPWR VGND sg13g2_fill_2
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_32_793 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
XFILLER_46_318 VPWR VGND sg13g2_decap_8
Xfanout41 net42 net41 VPWR VGND sg13g2_buf_1
XFILLER_42_568 VPWR VGND sg13g2_decap_8
Xfanout30 net42 net30 VPWR VGND sg13g2_buf_1
X_182_ data\[21\] data\[22\] net24 _029_ VPWR VGND sg13g2_mux2_1
X_320_ net40 VGND VPWR _080_ data\[73\] clknet_4_14_0_clk_regs sg13g2_dfrbpq_1
XFILLER_23_793 VPWR VGND sg13g2_decap_8
X_251_ net36 VGND VPWR _011_ data\[4\] clknet_4_7_0_clk_regs sg13g2_dfrbpq_1
XFILLER_2_653 VPWR VGND sg13g2_decap_8
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_45_340 VPWR VGND sg13g2_decap_4
XFILLER_14_793 VPWR VGND sg13g2_decap_8
XFILLER_49_690 VPWR VGND sg13g2_decap_8
Xclkload5 VPWR clkload5/Y clknet_4_11_0_clk_regs VGND sg13g2_inv_1
XFILLER_34_17 VPWR VGND sg13g2_fill_1
XFILLER_47_616 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_43_811 VPWR VGND sg13g2_decap_8
X_234_ data\[73\] data\[74\] net27 _081_ VPWR VGND sg13g2_mux2_1
X_303_ net33 VGND VPWR _063_ data\[56\] clknet_4_6_0_clk_regs sg13g2_dfrbpq_1
X_165_ data\[4\] data\[5\] net21 _012_ VPWR VGND sg13g2_mux2_1
XFILLER_34_800 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_46_682 VPWR VGND sg13g2_decap_8
XFILLER_25_800 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_8
XFILLER_40_858 VPWR VGND sg13g2_decap_4
XFILLER_40_814 VPWR VGND sg13g2_decap_8
XFILLER_3_214 VPWR VGND sg13g2_fill_1
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_31_814 VPWR VGND sg13g2_decap_8
XFILLER_43_685 VPWR VGND sg13g2_decap_8
X_148_ _108_ VPWR _109_ VGND u_shift_reg.bit_count\[2\] _106_ sg13g2_o21ai_1
X_217_ data\[56\] data\[57\] net18 _064_ VPWR VGND sg13g2_mux2_1
XFILLER_2_291 VPWR VGND sg13g2_fill_2
XFILLER_3_781 VPWR VGND sg13g2_decap_8
XFILLER_32_4 VPWR VGND sg13g2_decap_8
XFILLER_22_814 VPWR VGND sg13g2_decap_8
XFILLER_31_18 VPWR VGND sg13g2_decap_8
XFILLER_0_228 VPWR VGND sg13g2_fill_1
XFILLER_9_807 VPWR VGND sg13g2_decap_8
XFILLER_13_814 VPWR VGND sg13g2_decap_8
XFILLER_48_700 VPWR VGND sg13g2_decap_8
XFILLER_0_762 VPWR VGND sg13g2_decap_8
XFILLER_48_777 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_23_0 VPWR VGND sg13g2_fill_2
XFILLER_26_18 VPWR VGND sg13g2_decap_4
XFILLER_10_828 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_45_736 VPWR VGND sg13g2_decap_8
XFILLER_26_961 VPWR VGND sg13g2_decap_8
XFILLER_44_257 VPWR VGND sg13g2_decap_8
XFILLER_5_821 VPWR VGND sg13g2_decap_4
XFILLER_44_791 VPWR VGND sg13g2_decap_8
XFILLER_48_574 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_45_533 VPWR VGND sg13g2_decap_8
XFILLER_41_772 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_32_772 VPWR VGND sg13g2_decap_8
XFILLER_17_791 VPWR VGND sg13g2_decap_8
XFILLER_2_109 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
Xfanout20 net22 net20 VPWR VGND sg13g2_buf_1
X_181_ data\[20\] data\[21\] net24 _028_ VPWR VGND sg13g2_mux2_1
XFILLER_23_772 VPWR VGND sg13g2_decap_8
Xfanout31 net32 net31 VPWR VGND sg13g2_buf_1
Xfanout42 net1 net42 VPWR VGND sg13g2_buf_1
X_250_ net36 VGND VPWR _010_ data\[3\] clknet_4_7_0_clk_regs sg13g2_dfrbpq_1
XFILLER_2_632 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_1_186 VPWR VGND sg13g2_fill_1
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_14_772 VPWR VGND sg13g2_decap_8
XFILLER_45_396 VPWR VGND sg13g2_decap_8
XFILLER_37_842 VPWR VGND sg13g2_decap_8
Xclkload6 VPWR clkload6/Y clknet_4_13_0_clk_regs VGND sg13g2_inv_1
XFILLER_20_786 VPWR VGND sg13g2_decap_8
XFILLER_28_842 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_decap_8
X_302_ net33 VGND VPWR _062_ data\[55\] clknet_4_4_0_clk_regs sg13g2_dfrbpq_1
XFILLER_42_333 VPWR VGND sg13g2_decap_4
X_233_ data\[72\] data\[73\] net26 _080_ VPWR VGND sg13g2_mux2_1
XFILLER_7_779 VPWR VGND sg13g2_decap_8
XFILLER_11_786 VPWR VGND sg13g2_decap_8
X_164_ data\[3\] data\[4\] net21 _011_ VPWR VGND sg13g2_mux2_1
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_46_661 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_45_182 VPWR VGND sg13g2_decap_8
XFILLER_44_609 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
Xheichips25_template VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_31_848 VPWR VGND sg13g2_decap_8
XFILLER_43_664 VPWR VGND sg13g2_decap_8
XFILLER_42_130 VPWR VGND sg13g2_decap_4
XFILLER_42_163 VPWR VGND sg13g2_decap_8
X_147_ u_shift_reg.bit_count\[1\] u_shift_reg.bit_count\[2\] u_shift_reg.bit_count\[0\]
+ _108_ VPWR VGND _097_ sg13g2_nand4_1
X_216_ data\[55\] data\[56\] net18 _063_ VPWR VGND sg13g2_mux2_1
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_3_760 VPWR VGND sg13g2_decap_8
XFILLER_0_207 VPWR VGND sg13g2_decap_8
XFILLER_21_41 VPWR VGND sg13g2_decap_8
XFILLER_0_741 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_10_807 VPWR VGND sg13g2_decap_8
XFILLER_26_940 VPWR VGND sg13g2_decap_8
XFILLER_45_715 VPWR VGND sg13g2_decap_8
XFILLER_44_236 VPWR VGND sg13g2_decap_8
XFILLER_5_800 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_44_770 VPWR VGND sg13g2_decap_8
XFILLER_42_707 VPWR VGND sg13g2_decap_4
XFILLER_37_18 VPWR VGND sg13g2_fill_2
XFILLER_2_814 VPWR VGND sg13g2_decap_8
XFILLER_45_501 VPWR VGND sg13g2_decap_8
XFILLER_45_589 VPWR VGND sg13g2_decap_8
XFILLER_4_55 VPWR VGND sg13g2_fill_1
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_49_851 VPWR VGND sg13g2_decap_8
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
Xfanout21 net22 net21 VPWR VGND sg13g2_buf_1
XFILLER_13_42 VPWR VGND sg13g2_decap_8
XFILLER_13_31 VPWR VGND sg13g2_fill_1
XFILLER_13_20 VPWR VGND sg13g2_decap_8
X_180_ data\[19\] data\[20\] net24 _027_ VPWR VGND sg13g2_mux2_1
Xfanout32 net33 net32 VPWR VGND sg13g2_buf_1
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_2_611 VPWR VGND sg13g2_decap_8
XFILLER_2_688 VPWR VGND sg13g2_decap_8
XFILLER_46_843 VPWR VGND sg13g2_decap_8
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_45_375 VPWR VGND sg13g2_decap_8
XFILLER_37_821 VPWR VGND sg13g2_decap_8
Xclkload7 VPWR clkload7/Y clknet_4_14_0_clk_regs VGND sg13g2_inv_1
XFILLER_20_765 VPWR VGND sg13g2_decap_8
XFILLER_28_821 VPWR VGND sg13g2_decap_8
X_232_ data\[71\] data\[72\] net26 _079_ VPWR VGND sg13g2_mux2_1
X_301_ net31 VGND VPWR _061_ data\[54\] clknet_4_1_0_clk_regs sg13g2_dfrbpq_1
XFILLER_11_765 VPWR VGND sg13g2_decap_8
X_163_ data\[2\] data\[3\] net21 _010_ VPWR VGND sg13g2_mux2_1
XFILLER_49_60 VPWR VGND sg13g2_decap_8
XFILLER_34_835 VPWR VGND sg13g2_decap_4
XFILLER_46_640 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_46_0 VPWR VGND sg13g2_decap_8
XFILLER_25_835 VPWR VGND sg13g2_fill_1
XFILLER_10_54 VPWR VGND sg13g2_fill_2
XFILLER_43_643 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
X_215_ data\[54\] data\[55\] net17 _062_ VPWR VGND sg13g2_mux2_1
X_146_ _106_ _107_ _001_ VPWR VGND sg13g2_nor2_1
XFILLER_30_860 VPWR VGND sg13g2_fill_2
XFILLER_1_709 VPWR VGND sg13g2_decap_8
XFILLER_44_429 VPWR VGND sg13g2_decap_8
XFILLER_48_735 VPWR VGND sg13g2_decap_8
XFILLER_0_720 VPWR VGND sg13g2_decap_8
XFILLER_0_797 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_8_842 VPWR VGND sg13g2_decap_4
X_129_ _094_ _090_ clk1_out _089_ adc_data\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_27_919 VPWR VGND sg13g2_decap_8
XFILLER_39_779 VPWR VGND sg13g2_decap_8
XFILLER_27_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_26_996 VPWR VGND sg13g2_decap_8
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_0_594 VPWR VGND sg13g2_decap_8
XFILLER_35_793 VPWR VGND sg13g2_decap_8
XFILLER_27_52 VPWR VGND sg13g2_decap_4
XFILLER_26_793 VPWR VGND sg13g2_decap_8
XFILLER_45_568 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
Xclkbuf_4_6_0_clk_regs clknet_0_clk_regs clknet_4_6_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_49_830 VPWR VGND sg13g2_decap_8
Xfanout33 net42 net33 VPWR VGND sg13g2_buf_1
Xfanout22 net23 net22 VPWR VGND sg13g2_buf_1
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_2_667 VPWR VGND sg13g2_decap_8
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_46_822 VPWR VGND sg13g2_decap_8
XFILLER_45_354 VPWR VGND sg13g2_decap_8
XFILLER_37_800 VPWR VGND sg13g2_decap_8
Xclkload8 VPWR clkload8/Y clknet_4_15_0_clk_regs VGND sg13g2_inv_1
XFILLER_3_409 VPWR VGND sg13g2_decap_8
XFILLER_43_825 VPWR VGND sg13g2_decap_8
XFILLER_28_800 VPWR VGND sg13g2_decap_8
XFILLER_24_31 VPWR VGND sg13g2_decap_8
X_300_ net31 VGND VPWR _060_ data\[53\] clknet_4_1_0_clk_regs sg13g2_dfrbpq_1
X_231_ data\[70\] data\[71\] net26 _078_ VPWR VGND sg13g2_mux2_1
X_162_ data\[1\] data\[2\] net21 _009_ VPWR VGND sg13g2_mux2_1
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_19_800 VPWR VGND sg13g2_decap_8
XFILLER_34_858 VPWR VGND sg13g2_decap_4
XFILLER_34_814 VPWR VGND sg13g2_decap_8
XFILLER_46_696 VPWR VGND sg13g2_decap_8
XFILLER_45_140 VPWR VGND sg13g2_decap_8
XFILLER_39_0 VPWR VGND sg13g2_decap_4
XFILLER_25_814 VPWR VGND sg13g2_decap_8
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
XFILLER_40_839 VPWR VGND sg13g2_fill_2
XFILLER_40_828 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_43_622 VPWR VGND sg13g2_decap_8
XFILLER_43_699 VPWR VGND sg13g2_decap_8
X_214_ data\[53\] data\[54\] net17 _061_ VPWR VGND sg13g2_mux2_1
X_145_ VGND VPWR u_shift_reg.bit_count\[0\] _097_ _107_ u_shift_reg.bit_count\[1\]
+ sg13g2_a21oi_1
XFILLER_3_795 VPWR VGND sg13g2_decap_8
XFILLER_22_828 VPWR VGND sg13g2_decap_8
XFILLER_46_493 VPWR VGND sg13g2_decap_8
XFILLER_44_408 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_0_776 VPWR VGND sg13g2_decap_8
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
X_128_ VPWR net11 _093_ VGND sg13g2_inv_1
XFILLER_8_821 VPWR VGND sg13g2_decap_8
XFILLER_3_592 VPWR VGND sg13g2_decap_8
XFILLER_47_791 VPWR VGND sg13g2_decap_8
XFILLER_46_290 VPWR VGND sg13g2_decap_8
XFILLER_26_975 VPWR VGND sg13g2_decap_8
XFILLER_5_846 VPWR VGND sg13g2_fill_2
XFILLER_5_835 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_0_573 VPWR VGND sg13g2_decap_8
XFILLER_48_588 VPWR VGND sg13g2_decap_8
XFILLER_35_772 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_45_547 VPWR VGND sg13g2_decap_8
XFILLER_41_786 VPWR VGND sg13g2_decap_8
XFILLER_26_772 VPWR VGND sg13g2_decap_8
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_17_772 VPWR VGND sg13g2_decap_8
XFILLER_32_786 VPWR VGND sg13g2_decap_8
Xfanout34 net37 net34 VPWR VGND sg13g2_buf_1
XFILLER_23_786 VPWR VGND sg13g2_decap_8
Xfanout23 _098_ net23 VPWR VGND sg13g2_buf_1
XFILLER_46_801 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_fill_2
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_2_646 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_14_786 VPWR VGND sg13g2_decap_8
XFILLER_37_856 VPWR VGND sg13g2_decap_4
XFILLER_49_683 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_47_609 VPWR VGND sg13g2_decap_8
XFILLER_43_804 VPWR VGND sg13g2_decap_8
XFILLER_28_856 VPWR VGND sg13g2_decap_4
XFILLER_46_119 VPWR VGND sg13g2_fill_1
X_230_ data\[69\] data\[70\] net26 _077_ VPWR VGND sg13g2_mux2_1
X_161_ data\[0\] data\[1\] net21 _008_ VPWR VGND sg13g2_mux2_1
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_46_675 VPWR VGND sg13g2_decap_8
XFILLER_45_196 VPWR VGND sg13g2_decap_8
XFILLER_6_793 VPWR VGND sg13g2_decap_8
XFILLER_49_480 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
XFILLER_40_807 VPWR VGND sg13g2_decap_8
XFILLER_19_54 VPWR VGND sg13g2_fill_2
XFILLER_19_32 VPWR VGND sg13g2_decap_4
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_31_807 VPWR VGND sg13g2_decap_8
XFILLER_43_678 VPWR VGND sg13g2_decap_8
XFILLER_43_601 VPWR VGND sg13g2_decap_8
X_213_ data\[52\] data\[53\] net15 _060_ VPWR VGND sg13g2_mux2_1
X_144_ _106_ u_shift_reg.bit_count\[0\] u_shift_reg.bit_count\[1\] _097_ VPWR VGND
+ sg13g2_and3_1
XFILLER_3_774 VPWR VGND sg13g2_decap_8
XFILLER_46_472 VPWR VGND sg13g2_decap_8
XFILLER_22_807 VPWR VGND sg13g2_decap_8
XFILLER_13_807 VPWR VGND sg13g2_decap_8
XFILLER_21_55 VPWR VGND sg13g2_fill_1
XFILLER_0_755 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_8_800 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_127_ _093_ _090_ clk2_out _089_ adc_data\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_560 VPWR VGND sg13g2_fill_1
XFILLER_3_571 VPWR VGND sg13g2_decap_8
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_45_729 VPWR VGND sg13g2_decap_8
XFILLER_26_954 VPWR VGND sg13g2_decap_8
XFILLER_5_814 VPWR VGND sg13g2_decap_8
XFILLER_0_552 VPWR VGND sg13g2_decap_8
XFILLER_44_784 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_decap_8
XFILLER_43_272 VPWR VGND sg13g2_decap_4
XFILLER_1_316 VPWR VGND sg13g2_fill_2
XFILLER_45_526 VPWR VGND sg13g2_decap_8
XFILLER_45_515 VPWR VGND sg13g2_fill_1
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_41_765 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_32_765 VPWR VGND sg13g2_decap_8
XFILLER_44_581 VPWR VGND sg13g2_decap_8
Xfanout35 net37 net35 VPWR VGND sg13g2_buf_1
Xfanout24 net25 net24 VPWR VGND sg13g2_buf_1
XFILLER_23_765 VPWR VGND sg13g2_decap_8
XFILLER_2_625 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_46_857 VPWR VGND sg13g2_decap_4
XFILLER_14_765 VPWR VGND sg13g2_decap_8
XFILLER_45_389 VPWR VGND sg13g2_decap_8
XFILLER_37_835 VPWR VGND sg13g2_decap_8
XFILLER_49_662 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_20_779 VPWR VGND sg13g2_decap_8
XFILLER_28_835 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_fill_2
XFILLER_42_326 VPWR VGND sg13g2_decap_8
XFILLER_42_337 VPWR VGND sg13g2_fill_1
XFILLER_24_55 VPWR VGND sg13g2_fill_1
XFILLER_11_779 VPWR VGND sg13g2_decap_8
X_160_ data\[0\] net3 _097_ _007_ VPWR VGND sg13g2_mux2_1
XFILLER_2_433 VPWR VGND sg13g2_fill_1
XFILLER_46_654 VPWR VGND sg13g2_decap_8
XFILLER_49_74 VPWR VGND sg13g2_decap_8
XFILLER_45_175 VPWR VGND sg13g2_decap_8
XFILLER_6_772 VPWR VGND sg13g2_decap_8
X_289_ net32 VGND VPWR _049_ data\[42\] clknet_4_5_0_clk_regs sg13g2_dfrbpq_1
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
XFILLER_33_860 VPWR VGND sg13g2_fill_2
XFILLER_43_657 VPWR VGND sg13g2_decap_8
X_212_ data\[51\] data\[52\] net14 _059_ VPWR VGND sg13g2_mux2_1
XFILLER_35_21 VPWR VGND sg13g2_fill_1
XFILLER_42_123 VPWR VGND sg13g2_decap_8
XFILLER_42_134 VPWR VGND sg13g2_fill_2
X_143_ u_shift_reg.bit_count\[0\] u_shift_reg.bit_count\[1\] _105_ VPWR VGND sg13g2_and2_1
XFILLER_2_230 VPWR VGND sg13g2_decap_4
XFILLER_3_753 VPWR VGND sg13g2_decap_8
XFILLER_46_451 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_8
XFILLER_21_12 VPWR VGND sg13g2_fill_2
XFILLER_0_734 VPWR VGND sg13g2_decap_8
XFILLER_48_749 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_43_454 VPWR VGND sg13g2_decap_8
X_126_ VPWR net10 _092_ VGND sg13g2_inv_1
XFILLER_16_4 VPWR VGND sg13g2_decap_4
XFILLER_26_933 VPWR VGND sg13g2_decap_8
XFILLER_38_793 VPWR VGND sg13g2_decap_8
XFILLER_45_708 VPWR VGND sg13g2_decap_8
XFILLER_16_23 VPWR VGND sg13g2_decap_4
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_44_763 VPWR VGND sg13g2_decap_8
XFILLER_29_793 VPWR VGND sg13g2_decap_8
XFILLER_2_807 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_49_844 VPWR VGND sg13g2_decap_8
XFILLER_0_361 VPWR VGND sg13g2_fill_1
XFILLER_0_372 VPWR VGND sg13g2_decap_8
XFILLER_0_383 VPWR VGND sg13g2_fill_2
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_44_560 VPWR VGND sg13g2_decap_8
Xfanout14 net15 net14 VPWR VGND sg13g2_buf_1
XFILLER_13_13 VPWR VGND sg13g2_decap_8
Xfanout36 net37 net36 VPWR VGND sg13g2_buf_1
Xfanout25 _098_ net25 VPWR VGND sg13g2_buf_1
XFILLER_8_6 VPWR VGND sg13g2_fill_1
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_2_604 VPWR VGND sg13g2_decap_8
XFILLER_46_836 VPWR VGND sg13g2_decap_8
XFILLER_45_368 VPWR VGND sg13g2_decap_8
XFILLER_49_641 VPWR VGND sg13g2_decap_8
XFILLER_1_681 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_37_814 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_28_814 VPWR VGND sg13g2_decap_8
Xclkbuf_4_5_0_clk_regs clknet_0_clk_regs clknet_4_5_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_43_839 VPWR VGND sg13g2_decap_4
XFILLER_40_55 VPWR VGND sg13g2_fill_1
XFILLER_2_478 VPWR VGND sg13g2_fill_2
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_27_891 VPWR VGND sg13g2_decap_8
XFILLER_34_839 VPWR VGND sg13g2_fill_2
XFILLER_34_828 VPWR VGND sg13g2_decap_8
XFILLER_46_633 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_814 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_42_861 VPWR VGND sg13g2_fill_1
X_288_ net31 VGND VPWR _048_ data\[41\] clknet_4_1_0_clk_regs sg13g2_dfrbpq_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
XFILLER_25_828 VPWR VGND sg13g2_decap_8
XFILLER_35_11 VPWR VGND sg13g2_fill_1
XFILLER_43_636 VPWR VGND sg13g2_decap_8
X_211_ data\[50\] data\[51\] net14 _058_ VPWR VGND sg13g2_mux2_1
X_142_ VGND VPWR u_shift_reg.bit_count\[0\] _097_ _000_ _104_ sg13g2_a21oi_1
XFILLER_42_146 VPWR VGND sg13g2_decap_8
XFILLER_3_732 VPWR VGND sg13g2_decap_8
XFILLER_2_253 VPWR VGND sg13g2_fill_1
XFILLER_46_430 VPWR VGND sg13g2_decap_8
XFILLER_30_842 VPWR VGND sg13g2_decap_8
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_decap_8
XFILLER_0_713 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_43_422 VPWR VGND sg13g2_decap_4
X_125_ _092_ _090_ osc_out _089_ adc_data\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_8_846 VPWR VGND sg13g2_fill_2
XFILLER_8_835 VPWR VGND sg13g2_decap_8
XFILLER_26_989 VPWR VGND sg13g2_decap_8
XFILLER_26_912 VPWR VGND sg13g2_decap_8
XFILLER_38_772 VPWR VGND sg13g2_decap_8
XFILLER_44_208 VPWR VGND sg13g2_fill_2
XFILLER_32_23 VPWR VGND sg13g2_decap_4
XFILLER_29_772 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_0_587 VPWR VGND sg13g2_decap_8
XFILLER_44_742 VPWR VGND sg13g2_decap_8
XFILLER_26_1010 VPWR VGND sg13g2_decap_8
XFILLER_3_370 VPWR VGND sg13g2_decap_4
XFILLER_35_786 VPWR VGND sg13g2_decap_8
XFILLER_27_45 VPWR VGND sg13g2_decap_8
XFILLER_26_786 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_49_823 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_0_395 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_17_786 VPWR VGND sg13g2_fill_1
Xfanout15 net16 net15 VPWR VGND sg13g2_buf_1
Xfanout26 net27 net26 VPWR VGND sg13g2_buf_1
Xfanout37 net42 net37 VPWR VGND sg13g2_buf_1
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_46_815 VPWR VGND sg13g2_decap_8
XFILLER_49_620 VPWR VGND sg13g2_decap_8
XFILLER_1_660 VPWR VGND sg13g2_decap_8
XFILLER_49_697 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_9_793 VPWR VGND sg13g2_decap_8
XFILLER_43_818 VPWR VGND sg13g2_decap_8
XFILLER_24_24 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_34_807 VPWR VGND sg13g2_decap_8
XFILLER_27_870 VPWR VGND sg13g2_decap_8
XFILLER_46_689 VPWR VGND sg13g2_decap_8
XFILLER_46_612 VPWR VGND sg13g2_decap_8
XFILLER_45_133 VPWR VGND sg13g2_decap_8
X_287_ net31 VGND VPWR _047_ data\[40\] clknet_4_0_0_clk_regs sg13g2_dfrbpq_1
XFILLER_39_4 VPWR VGND sg13g2_fill_2
XFILLER_49_494 VPWR VGND sg13g2_decap_8
XFILLER_25_807 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
XFILLER_43_615 VPWR VGND sg13g2_decap_8
X_210_ data\[49\] data\[50\] net14 _057_ VPWR VGND sg13g2_mux2_1
X_141_ VGND VPWR _097_ _102_ _104_ u_shift_reg.bit_count\[0\] sg13g2_a21oi_1
XFILLER_3_711 VPWR VGND sg13g2_decap_8
XFILLER_3_788 VPWR VGND sg13g2_decap_8
XFILLER_30_821 VPWR VGND sg13g2_decap_8
XFILLER_46_486 VPWR VGND sg13g2_decap_8
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
XFILLER_21_832 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_0_769 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
X_124_ VPWR net9 _091_ VGND sg13g2_inv_1
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_8_814 VPWR VGND sg13g2_decap_8
XFILLER_3_530 VPWR VGND sg13g2_fill_2
XFILLER_3_585 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_46_283 VPWR VGND sg13g2_decap_8
XFILLER_26_968 VPWR VGND sg13g2_decap_8
XFILLER_0_533 VPWR VGND sg13g2_fill_2
XFILLER_44_721 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_0_566 VPWR VGND sg13g2_decap_8
XFILLER_44_798 VPWR VGND sg13g2_decap_8
XFILLER_43_231 VPWR VGND sg13g2_fill_1
XFILLER_3_393 VPWR VGND sg13g2_decap_4
XFILLER_35_765 VPWR VGND sg13g2_decap_8
XFILLER_47_581 VPWR VGND sg13g2_decap_8
XFILLER_41_779 VPWR VGND sg13g2_decap_8
XFILLER_26_765 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_49_802 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_17_765 VPWR VGND sg13g2_decap_8
XFILLER_17_798 VPWR VGND sg13g2_decap_8
XFILLER_32_779 VPWR VGND sg13g2_decap_8
XFILLER_44_595 VPWR VGND sg13g2_decap_8
XFILLER_12_0 VPWR VGND sg13g2_fill_2
Xfanout16 net23 net16 VPWR VGND sg13g2_buf_1
Xfanout38 net39 net38 VPWR VGND sg13g2_buf_1
XFILLER_23_779 VPWR VGND sg13g2_decap_8
Xfanout27 _098_ net27 VPWR VGND sg13g2_buf_1
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_2_639 VPWR VGND sg13g2_decap_8
XFILLER_38_23 VPWR VGND sg13g2_decap_4
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_14_779 VPWR VGND sg13g2_decap_8
XFILLER_37_849 VPWR VGND sg13g2_decap_8
XFILLER_49_676 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_9_772 VPWR VGND sg13g2_decap_8
XFILLER_36_860 VPWR VGND sg13g2_fill_2
XFILLER_28_849 VPWR VGND sg13g2_decap_8
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_42_852 VPWR VGND sg13g2_decap_8
XFILLER_46_668 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
X_286_ net28 VGND VPWR _046_ data\[39\] clknet_4_0_0_clk_regs sg13g2_dfrbpq_1
XFILLER_10_793 VPWR VGND sg13g2_decap_8
XFILLER_6_786 VPWR VGND sg13g2_decap_8
XFILLER_49_473 VPWR VGND sg13g2_decap_8
XFILLER_19_47 VPWR VGND sg13g2_decap_8
XFILLER_19_36 VPWR VGND sg13g2_fill_1
XFILLER_19_25 VPWR VGND sg13g2_decap_8
X_140_ VPWR _103_ _102_ VGND sg13g2_inv_1
XFILLER_2_200 VPWR VGND sg13g2_fill_2
XFILLER_3_767 VPWR VGND sg13g2_decap_8
XFILLER_46_465 VPWR VGND sg13g2_decap_8
XFILLER_30_800 VPWR VGND sg13g2_decap_8
XFILLER_42_693 VPWR VGND sg13g2_decap_8
X_269_ net38 VGND VPWR _029_ data\[22\] clknet_4_13_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_21_811 VPWR VGND sg13g2_decap_8
XFILLER_21_48 VPWR VGND sg13g2_decap_8
XFILLER_0_748 VPWR VGND sg13g2_decap_8
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_12_800 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
X_123_ _091_ _090_ stable _089_ adc_data\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_542 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_46_262 VPWR VGND sg13g2_decap_8
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_26_947 VPWR VGND sg13g2_decap_8
XFILLER_5_807 VPWR VGND sg13g2_decap_8
XFILLER_0_545 VPWR VGND sg13g2_decap_8
XFILLER_44_700 VPWR VGND sg13g2_decap_8
XFILLER_44_777 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_fill_2
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_1_309 VPWR VGND sg13g2_decap_8
XFILLER_45_519 VPWR VGND sg13g2_decap_8
XFILLER_45_508 VPWR VGND sg13g2_decap_8
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_49_858 VPWR VGND sg13g2_decap_4
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_44_574 VPWR VGND sg13g2_decap_8
Xfanout28 net29 net28 VPWR VGND sg13g2_buf_1
XFILLER_13_27 VPWR VGND sg13g2_decap_4
Xfanout17 net23 net17 VPWR VGND sg13g2_buf_1
Xfanout39 net42 net39 VPWR VGND sg13g2_buf_1
XFILLER_13_49 VPWR VGND sg13g2_decap_8
XFILLER_2_618 VPWR VGND sg13g2_decap_8
XFILLER_37_828 VPWR VGND sg13g2_decap_8
XFILLER_49_655 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_1_695 VPWR VGND sg13g2_decap_8
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_45_861 VPWR VGND sg13g2_fill_1
XFILLER_44_371 VPWR VGND sg13g2_decap_8
XFILLER_28_828 VPWR VGND sg13g2_decap_8
XFILLER_24_48 VPWR VGND sg13g2_decap_8
XFILLER_2_426 VPWR VGND sg13g2_decap_8
XFILLER_46_647 VPWR VGND sg13g2_decap_8
XFILLER_49_67 VPWR VGND sg13g2_decap_8
XFILLER_42_831 VPWR VGND sg13g2_decap_8
XFILLER_45_168 VPWR VGND sg13g2_decap_8
X_285_ net38 VGND VPWR _045_ data\[38\] clknet_4_10_0_clk_regs sg13g2_dfrbpq_1
XFILLER_6_765 VPWR VGND sg13g2_decap_8
XFILLER_10_772 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_45_680 VPWR VGND sg13g2_decap_8
XFILLER_49_452 VPWR VGND sg13g2_decap_8
XFILLER_33_842 VPWR VGND sg13g2_decap_8
XFILLER_2_234 VPWR VGND sg13g2_fill_1
XFILLER_3_746 VPWR VGND sg13g2_decap_8
XFILLER_46_444 VPWR VGND sg13g2_decap_8
XFILLER_30_856 VPWR VGND sg13g2_decap_4
Xclkbuf_4_4_0_clk_regs clknet_0_clk_regs clknet_4_4_0_clk_regs VPWR VGND sg13g2_buf_8
X_199_ data\[38\] data\[39\] net14 _046_ VPWR VGND sg13g2_mux2_1
X_268_ net38 VGND VPWR _028_ data\[21\] clknet_4_13_0_clk_regs sg13g2_dfrbpq_1
XFILLER_2_95 VPWR VGND sg13g2_decap_8
XFILLER_0_727 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
X_122_ net5 net4 _090_ VPWR VGND sg13g2_nor2_1
XFILLER_16_8 VPWR VGND sg13g2_fill_1
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_46_241 VPWR VGND sg13g2_decap_8
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_26_926 VPWR VGND sg13g2_decap_8
XFILLER_38_786 VPWR VGND sg13g2_decap_8
XFILLER_16_16 VPWR VGND sg13g2_decap_8
XFILLER_16_27 VPWR VGND sg13g2_fill_2
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_44_756 VPWR VGND sg13g2_decap_8
XFILLER_29_786 VPWR VGND sg13g2_decap_8
XFILLER_43_200 VPWR VGND sg13g2_decap_8
XFILLER_25_992 VPWR VGND sg13g2_decap_8
XFILLER_26_1024 VPWR VGND sg13g2_decap_4
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_49_837 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_44_553 VPWR VGND sg13g2_decap_8
Xfanout29 net30 net29 VPWR VGND sg13g2_buf_1
Xfanout18 net23 net18 VPWR VGND sg13g2_buf_1
XFILLER_46_829 VPWR VGND sg13g2_decap_8
XFILLER_49_634 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_1_674 VPWR VGND sg13g2_decap_8
XFILLER_37_807 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_28_807 VPWR VGND sg13g2_decap_8
XFILLER_40_15 VPWR VGND sg13g2_fill_2
Xu_adc VPWR VGND data\[67\] data\[68\] data\[69\] data\[70\] data\[71\] data\[72\]
+ data\[73\] data\[74\] clknet_1_0__leaf_clk adc_data\[0\] adc_data\[1\] adc_data\[2\]
+ adc_data\[3\] adc_data\[4\] adc_data\[5\] adc_data\[6\] adc_data\[7\] u_adc/ready
+ data\[66\] adc
XFILLER_49_46 VPWR VGND sg13g2_decap_8
XFILLER_46_626 VPWR VGND sg13g2_decap_8
XFILLER_19_807 VPWR VGND sg13g2_decap_8
XFILLER_45_147 VPWR VGND sg13g2_fill_2
XFILLER_27_884 VPWR VGND sg13g2_decap_8
XFILLER_42_810 VPWR VGND sg13g2_decap_8
X_284_ net38 VGND VPWR _044_ data\[37\] clknet_4_10_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_431 VPWR VGND sg13g2_decap_8
XFILLER_33_821 VPWR VGND sg13g2_decap_8
XFILLER_43_629 VPWR VGND sg13g2_decap_8
XFILLER_24_821 VPWR VGND sg13g2_decap_8
XFILLER_2_202 VPWR VGND sg13g2_fill_1
XFILLER_3_725 VPWR VGND sg13g2_decap_8
XFILLER_2_246 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_15_843 VPWR VGND sg13g2_decap_4
XFILLER_46_423 VPWR VGND sg13g2_decap_8
XFILLER_30_835 VPWR VGND sg13g2_decap_8
X_267_ net38 VGND VPWR _027_ data\[20\] clknet_4_13_0_clk_regs sg13g2_dfrbpq_1
X_198_ data\[37\] data\[38\] net24 _045_ VPWR VGND sg13g2_mux2_1
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_21_846 VPWR VGND sg13g2_fill_2
XFILLER_0_706 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_43_415 VPWR VGND sg13g2_decap_8
XFILLER_43_426 VPWR VGND sg13g2_fill_1
X_121_ adc_data\[2\] _089_ net8 VPWR VGND sg13g2_and2_1
XFILLER_8_828 VPWR VGND sg13g2_decap_8
XFILLER_47_721 VPWR VGND sg13g2_decap_8
XFILLER_3_599 VPWR VGND sg13g2_decap_8
XFILLER_46_220 VPWR VGND sg13g2_decap_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_46_297 VPWR VGND sg13g2_decap_8
X_319_ net40 VGND VPWR _079_ data\[72\] clknet_4_12_0_clk_regs sg13g2_dfrbpq_1
Xclkbuf_1_0__f_clk clknet_1_0__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_26_905 VPWR VGND sg13g2_decap_8
XFILLER_38_765 VPWR VGND sg13g2_decap_8
XFILLER_32_16 VPWR VGND sg13g2_decap_8
XFILLER_32_27 VPWR VGND sg13g2_fill_2
XFILLER_29_765 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_44_735 VPWR VGND sg13g2_decap_8
XFILLER_25_971 VPWR VGND sg13g2_decap_8
XFILLER_26_1003 VPWR VGND sg13g2_decap_8
XFILLER_3_363 VPWR VGND sg13g2_decap_8
XFILLER_3_374 VPWR VGND sg13g2_fill_1
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_14_6 VPWR VGND sg13g2_fill_1
XFILLER_43_790 VPWR VGND sg13g2_decap_8
XFILLER_35_779 VPWR VGND sg13g2_decap_8
XFILLER_8_40 VPWR VGND sg13g2_decap_8
XFILLER_26_779 VPWR VGND sg13g2_decap_8
XFILLER_49_816 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_17_779 VPWR VGND sg13g2_decap_8
XFILLER_40_793 VPWR VGND sg13g2_decap_8
Xfanout19 net22 net19 VPWR VGND sg13g2_buf_1
XFILLER_47_392 VPWR VGND sg13g2_decap_8
XFILLER_31_793 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_46_808 VPWR VGND sg13g2_decap_8
XFILLER_45_329 VPWR VGND sg13g2_fill_1
XFILLER_22_793 VPWR VGND sg13g2_decap_8
XFILLER_49_613 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_fill_1
XFILLER_1_653 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_45_841 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_9_786 VPWR VGND sg13g2_decap_8
XFILLER_13_793 VPWR VGND sg13g2_decap_8
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_24_17 VPWR VGND sg13g2_decap_8
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_27_863 VPWR VGND sg13g2_decap_8
XFILLER_46_605 VPWR VGND sg13g2_decap_8
XFILLER_45_126 VPWR VGND sg13g2_decap_8
X_283_ net35 VGND VPWR _043_ data\[36\] clknet_4_10_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_fill_1
XFILLER_33_800 VPWR VGND sg13g2_decap_8
XFILLER_18_841 VPWR VGND sg13g2_decap_8
XFILLER_43_608 VPWR VGND sg13g2_decap_8
XFILLER_24_800 VPWR VGND sg13g2_decap_8
XFILLER_35_27 VPWR VGND sg13g2_fill_2
XFILLER_24_844 VPWR VGND sg13g2_decap_4
XFILLER_3_704 VPWR VGND sg13g2_decap_8
XFILLER_46_402 VPWR VGND sg13g2_decap_8
XFILLER_30_814 VPWR VGND sg13g2_decap_8
XFILLER_42_652 VPWR VGND sg13g2_decap_8
XFILLER_46_479 VPWR VGND sg13g2_decap_8
X_197_ data\[36\] data\[37\] net20 _044_ VPWR VGND sg13g2_mux2_1
X_266_ net39 VGND VPWR _026_ data\[19\] clknet_4_12_0_clk_regs sg13g2_dfrbpq_1
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_21_825 VPWR VGND sg13g2_decap_8
X_120_ adc_data\[1\] _089_ net7 VPWR VGND sg13g2_and2_1
XFILLER_8_807 VPWR VGND sg13g2_decap_8
XFILLER_12_814 VPWR VGND sg13g2_decap_8
XFILLER_3_523 VPWR VGND sg13g2_decap_8
XFILLER_3_556 VPWR VGND sg13g2_decap_4
XFILLER_3_578 VPWR VGND sg13g2_decap_8
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_47_700 VPWR VGND sg13g2_decap_8
XFILLER_46_276 VPWR VGND sg13g2_decap_8
XFILLER_42_482 VPWR VGND sg13g2_fill_2
X_318_ net40 VGND VPWR _078_ data\[71\] clknet_4_12_0_clk_regs sg13g2_dfrbpq_1
X_249_ net36 VGND VPWR _009_ data\[2\] clknet_4_7_0_clk_regs sg13g2_dfrbpq_1
XFILLER_0_526 VPWR VGND sg13g2_decap_8
XFILLER_44_714 VPWR VGND sg13g2_decap_8
XFILLER_0_559 VPWR VGND sg13g2_decap_8
XFILLER_25_950 VPWR VGND sg13g2_decap_8
XFILLER_3_320 VPWR VGND sg13g2_decap_8
XFILLER_3_331 VPWR VGND sg13g2_fill_2
XFILLER_21_8 VPWR VGND sg13g2_decap_4
XFILLER_3_397 VPWR VGND sg13g2_fill_2
XFILLER_47_574 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
XFILLER_40_772 VPWR VGND sg13g2_decap_8
XFILLER_44_588 VPWR VGND sg13g2_decap_8
XFILLER_48_861 VPWR VGND sg13g2_fill_1
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_31_772 VPWR VGND sg13g2_decap_8
XFILLER_38_27 VPWR VGND sg13g2_fill_2
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_22_772 VPWR VGND sg13g2_decap_8
XFILLER_49_669 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_1_632 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_45_820 VPWR VGND sg13g2_decap_8
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_9_765 VPWR VGND sg13g2_decap_8
XFILLER_13_772 VPWR VGND sg13g2_decap_8
XFILLER_36_842 VPWR VGND sg13g2_decap_8
XFILLER_40_17 VPWR VGND sg13g2_fill_1
XFILLER_42_845 VPWR VGND sg13g2_decap_8
XFILLER_27_842 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_45_149 VPWR VGND sg13g2_fill_1
X_282_ net34 VGND VPWR _042_ data\[35\] clknet_4_8_0_clk_regs sg13g2_dfrbpq_1
XFILLER_10_786 VPWR VGND sg13g2_decap_8
XFILLER_6_779 VPWR VGND sg13g2_decap_8
XFILLER_30_50 VPWR VGND sg13g2_decap_4
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_33_856 VPWR VGND sg13g2_decap_4
XFILLER_45_694 VPWR VGND sg13g2_decap_8
XFILLER_19_18 VPWR VGND sg13g2_decap_8
XFILLER_46_458 VPWR VGND sg13g2_decap_8
XFILLER_42_686 VPWR VGND sg13g2_decap_8
XFILLER_42_631 VPWR VGND sg13g2_decap_8
X_196_ data\[35\] data\[36\] net20 _043_ VPWR VGND sg13g2_mux2_1
X_265_ net39 VGND VPWR _025_ data\[18\] clknet_4_12_0_clk_regs sg13g2_dfrbpq_1
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_2_793 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_45_480 VPWR VGND sg13g2_decap_8
XFILLER_21_804 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_11_52 VPWR VGND sg13g2_decap_4
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_46_255 VPWR VGND sg13g2_decap_8
X_317_ net40 VGND VPWR _077_ data\[70\] clknet_4_12_0_clk_regs sg13g2_dfrbpq_1
X_179_ data\[18\] data\[19\] net25 _026_ VPWR VGND sg13g2_mux2_1
X_248_ net36 VGND VPWR _008_ data\[1\] clknet_4_6_0_clk_regs sg13g2_dfrbpq_1
XFILLER_0_505 VPWR VGND sg13g2_decap_4
Xclkbuf_4_3_0_clk_regs clknet_0_clk_regs clknet_4_3_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_22_51 VPWR VGND sg13g2_decap_4
XFILLER_4_800 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_0_379 VPWR VGND sg13g2_decap_4
XFILLER_0_357 VPWR VGND sg13g2_decap_4
XFILLER_44_567 VPWR VGND sg13g2_decap_8
XFILLER_48_840 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
XFILLER_1_611 VPWR VGND sg13g2_decap_8
XFILLER_49_648 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_1_688 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_45_854 VPWR VGND sg13g2_decap_8
XFILLER_44_364 VPWR VGND sg13g2_decap_8
XFILLER_5_54 VPWR VGND sg13g2_fill_2
XFILLER_5_32 VPWR VGND sg13g2_decap_4
XFILLER_36_821 VPWR VGND sg13g2_decap_8
XFILLER_27_821 VPWR VGND sg13g2_decap_8
XFILLER_27_898 VPWR VGND sg13g2_decap_8
XFILLER_42_824 VPWR VGND sg13g2_decap_8
X_281_ net34 VGND VPWR _041_ data\[34\] clknet_4_9_0_clk_regs sg13g2_dfrbpq_1
XFILLER_10_765 VPWR VGND sg13g2_decap_8
XFILLER_45_673 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_18_821 VPWR VGND sg13g2_decap_8
XFILLER_33_835 VPWR VGND sg13g2_decap_8
XFILLER_24_835 VPWR VGND sg13g2_decap_4
XFILLER_3_739 VPWR VGND sg13g2_decap_8
XFILLER_15_802 VPWR VGND sg13g2_decap_8
XFILLER_46_437 VPWR VGND sg13g2_decap_8
XFILLER_30_849 VPWR VGND sg13g2_decap_8
XFILLER_42_610 VPWR VGND sg13g2_decap_8
X_264_ net38 VGND VPWR _024_ data\[17\] clknet_4_12_0_clk_regs sg13g2_dfrbpq_1
X_195_ data\[34\] data\[35\] net19 _042_ VPWR VGND sg13g2_mux2_1
XFILLER_1_271 VPWR VGND sg13g2_fill_1
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_2_772 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_fill_2
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
XFILLER_46_234 VPWR VGND sg13g2_decap_8
X_316_ net40 VGND VPWR _076_ data\[69\] clknet_4_14_0_clk_regs sg13g2_dfrbpq_1
X_247_ net32 VGND VPWR _007_ data\[0\] clknet_4_5_0_clk_regs sg13g2_dfrbpq_1
XFILLER_42_462 VPWR VGND sg13g2_fill_2
XFILLER_42_484 VPWR VGND sg13g2_fill_1
X_178_ data\[17\] data\[18\] net24 _025_ VPWR VGND sg13g2_mux2_1
XFILLER_26_919 VPWR VGND sg13g2_decap_8
XFILLER_38_779 VPWR VGND sg13g2_decap_8
XFILLER_29_779 VPWR VGND sg13g2_decap_8
XFILLER_44_749 VPWR VGND sg13g2_decap_8
XFILLER_25_985 VPWR VGND sg13g2_decap_8
XFILLER_26_1017 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_8_54 VPWR VGND sg13g2_fill_2
XFILLER_34_793 VPWR VGND sg13g2_decap_8
XFILLER_1_804 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_44_546 VPWR VGND sg13g2_decap_8
XFILLER_17_41 VPWR VGND sg13g2_decap_8
XFILLER_25_793 VPWR VGND sg13g2_decap_8
XFILLER_3_196 VPWR VGND sg13g2_decap_4
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_1_667 VPWR VGND sg13g2_decap_8
XFILLER_49_627 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_36_800 VPWR VGND sg13g2_decap_8
XFILLER_48_693 VPWR VGND sg13g2_decap_8
XFILLER_49_39 VPWR VGND sg13g2_decap_8
XFILLER_27_800 VPWR VGND sg13g2_decap_8
XFILLER_46_619 VPWR VGND sg13g2_decap_8
XFILLER_27_877 VPWR VGND sg13g2_decap_8
XFILLER_42_803 VPWR VGND sg13g2_decap_8
X_280_ net34 VGND VPWR _040_ data\[33\] clknet_4_9_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_424 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_fill_2
XFILLER_33_814 VPWR VGND sg13g2_decap_8
XFILLER_45_652 VPWR VGND sg13g2_decap_8
XFILLER_18_800 VPWR VGND sg13g2_decap_8
XFILLER_44_140 VPWR VGND sg13g2_fill_1
XFILLER_48_490 VPWR VGND sg13g2_decap_8
XFILLER_24_814 VPWR VGND sg13g2_decap_8
XFILLER_35_19 VPWR VGND sg13g2_fill_2
XFILLER_3_718 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk_regs clknet_0_clk_regs clk_regs VPWR VGND sg13g2_buf_16
XFILLER_2_239 VPWR VGND sg13g2_decap_8
XFILLER_15_836 VPWR VGND sg13g2_decap_8
XFILLER_46_416 VPWR VGND sg13g2_decap_8
XFILLER_30_828 VPWR VGND sg13g2_decap_8
XFILLER_42_666 VPWR VGND sg13g2_decap_4
X_263_ net38 VGND VPWR _023_ data\[16\] clknet_4_13_0_clk_regs sg13g2_dfrbpq_1
XFILLER_15_847 VPWR VGND sg13g2_fill_1
X_194_ data\[33\] data\[34\] net19 _041_ VPWR VGND sg13g2_mux2_1
XFILLER_2_751 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
XFILLER_21_839 VPWR VGND sg13g2_decap_8
XFILLER_47_714 VPWR VGND sg13g2_decap_8
XFILLER_46_213 VPWR VGND sg13g2_decap_8
X_177_ data\[16\] data\[17\] net24 _024_ VPWR VGND sg13g2_mux2_1
X_315_ net40 VGND VPWR _075_ data\[68\] clknet_4_14_0_clk_regs sg13g2_dfrbpq_1
X_246_ net31 VGND VPWR _006_ u_shift_reg.bit_count\[6\] clknet_4_4_0_clk_regs sg13g2_dfrbpq_1
XFILLER_46_780 VPWR VGND sg13g2_decap_8
XFILLER_44_728 VPWR VGND sg13g2_decap_8
XFILLER_25_964 VPWR VGND sg13g2_decap_8
XFILLER_22_20 VPWR VGND sg13g2_fill_1
XFILLER_3_312 VPWR VGND sg13g2_fill_2
XFILLER_47_588 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_43_783 VPWR VGND sg13g2_decap_8
XFILLER_42_293 VPWR VGND sg13g2_decap_4
X_229_ data\[68\] data\[69\] net26 _076_ VPWR VGND sg13g2_mux2_1
XFILLER_34_772 VPWR VGND sg13g2_decap_8
XFILLER_49_809 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_25_772 VPWR VGND sg13g2_decap_8
XFILLER_40_786 VPWR VGND sg13g2_decap_8
XFILLER_3_164 VPWR VGND sg13g2_decap_4
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_31_786 VPWR VGND sg13g2_decap_8
XFILLER_43_580 VPWR VGND sg13g2_decap_8
XFILLER_16_772 VPWR VGND sg13g2_decap_8
XFILLER_39_831 VPWR VGND sg13g2_decap_8
XFILLER_22_786 VPWR VGND sg13g2_decap_8
XFILLER_49_606 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_1_646 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_45_834 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_13_786 VPWR VGND sg13g2_decap_8
XFILLER_44_84 VPWR VGND sg13g2_decap_8
XFILLER_9_779 VPWR VGND sg13g2_decap_8
XFILLER_48_672 VPWR VGND sg13g2_decap_8
XFILLER_36_856 VPWR VGND sg13g2_decap_4
XFILLER_47_182 VPWR VGND sg13g2_decap_8
XFILLER_49_18 VPWR VGND sg13g2_decap_8
XFILLER_27_856 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_42_859 VPWR VGND sg13g2_fill_2
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_39_40 VPWR VGND sg13g2_decap_8
XFILLER_45_631 VPWR VGND sg13g2_decap_8
Xu_multimode_dll VPWR VGND data\[38\] clk0_out data\[20\] data\[21\] data\[22\] data\[23\]
+ data\[24\] clk1_out data\[25\] data\[26\] data\[27\] data\[28\] data\[29\] clk2_out
+ data\[30\] data\[31\] data\[32\] data\[33\] data\[34\] data\[39\] ena data\[40\]
+ data\[50\] data\[51\] data\[52\] data\[53\] data\[54\] data\[55\] data\[56\] data\[57\]
+ data\[58\] data\[59\] data\[41\] data\[60\] data\[61\] data\[62\] data\[63\] data\[64\]
+ data\[65\] data\[42\] data\[43\] data\[44\] data\[45\] data\[46\] data\[47\] data\[48\]
+ data\[49\] data\[5\] data\[6\] data\[7\] data\[8\] data\[9\] data\[10\] data\[11\]
+ data\[12\] data\[13\] data\[14\] data\[15\] data\[16\] data\[17\] data\[18\] data\[19\]
+ data\[0\] data\[1\] data\[2\] data\[3\] data\[4\] data\[35\] data\[36\] data\[37\]
+ clknet_1_0__leaf_clk osc_out net34 stable multimode_dll
XFILLER_5_793 VPWR VGND sg13g2_decap_8
XFILLER_42_645 VPWR VGND sg13g2_decap_8
XFILLER_30_807 VPWR VGND sg13g2_decap_8
X_193_ data\[32\] data\[33\] net19 _040_ VPWR VGND sg13g2_mux2_1
X_262_ net38 VGND VPWR _022_ data\[15\] clknet_4_13_0_clk_regs sg13g2_dfrbpq_1
XFILLER_41_52 VPWR VGND sg13g2_decap_4
XFILLER_2_730 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_21_818 VPWR VGND sg13g2_decap_8
XFILLER_45_494 VPWR VGND sg13g2_decap_8
XFILLER_12_807 VPWR VGND sg13g2_decap_8
XFILLER_11_33 VPWR VGND sg13g2_fill_2
XFILLER_3_516 VPWR VGND sg13g2_decap_8
XFILLER_3_549 VPWR VGND sg13g2_decap_8
X_314_ net40 VGND VPWR _074_ data\[67\] clknet_4_14_0_clk_regs sg13g2_dfrbpq_1
XFILLER_46_269 VPWR VGND sg13g2_decap_8
XFILLER_42_464 VPWR VGND sg13g2_fill_1
XFILLER_42_475 VPWR VGND sg13g2_decap_8
X_176_ data\[15\] data\[16\] net24 _023_ VPWR VGND sg13g2_mux2_1
XFILLER_7_800 VPWR VGND sg13g2_decap_8
X_245_ net31 VGND VPWR _005_ u_shift_reg.bit_count\[5\] clknet_4_4_0_clk_regs sg13g2_dfrbpq_1
XFILLER_42_7 VPWR VGND sg13g2_decap_8
XFILLER_45_280 VPWR VGND sg13g2_decap_8
XFILLER_0_519 VPWR VGND sg13g2_decap_8
XFILLER_44_707 VPWR VGND sg13g2_decap_8
XFILLER_25_943 VPWR VGND sg13g2_decap_8
XFILLER_4_814 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
XFILLER_43_762 VPWR VGND sg13g2_decap_8
XFILLER_8_23 VPWR VGND sg13g2_decap_8
XFILLER_42_261 VPWR VGND sg13g2_decap_8
X_228_ data\[67\] data\[68\] net26 _075_ VPWR VGND sg13g2_mux2_1
X_159_ _114_ u_shift_reg.bit_count\[6\] _006_ VPWR VGND sg13g2_xor2_1
XFILLER_40_765 VPWR VGND sg13g2_decap_8
XFILLER_33_53 VPWR VGND sg13g2_fill_2
XFILLER_48_854 VPWR VGND sg13g2_decap_8
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_31_765 VPWR VGND sg13g2_decap_8
Xclkbuf_4_2_0_clk_regs clknet_0_clk_regs clknet_4_2_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_22_765 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_1_625 VPWR VGND sg13g2_decap_8
XFILLER_45_813 VPWR VGND sg13g2_decap_8
XFILLER_44_312 VPWR VGND sg13g2_decap_8
XFILLER_13_765 VPWR VGND sg13g2_decap_8
XFILLER_44_63 VPWR VGND sg13g2_decap_8
XFILLER_36_835 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_42_838 VPWR VGND sg13g2_decap_8
XFILLER_27_835 VPWR VGND sg13g2_decap_8
XFILLER_10_779 VPWR VGND sg13g2_decap_8
XFILLER_30_54 VPWR VGND sg13g2_fill_2
XFILLER_45_610 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_33_849 VPWR VGND sg13g2_decap_8
XFILLER_45_687 VPWR VGND sg13g2_decap_8
XFILLER_5_772 VPWR VGND sg13g2_decap_8
XFILLER_32_860 VPWR VGND sg13g2_fill_2
XFILLER_42_624 VPWR VGND sg13g2_decap_8
X_261_ net35 VGND VPWR _021_ data\[14\] clknet_4_9_0_clk_regs sg13g2_dfrbpq_1
X_192_ data\[31\] data\[32\] net19 _039_ VPWR VGND sg13g2_mux2_1
XFILLER_41_31 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_2_786 VPWR VGND sg13g2_decap_8
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_45_473 VPWR VGND sg13g2_decap_8
Xclkbuf_4_15_0_clk_regs clknet_0_clk_regs clknet_4_15_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_11_45 VPWR VGND sg13g2_decap_8
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_46_248 VPWR VGND sg13g2_decap_8
X_313_ net40 VGND VPWR _073_ data\[66\] clknet_4_14_0_clk_regs sg13g2_dfrbpq_1
X_244_ net32 VGND VPWR _004_ u_shift_reg.bit_count\[4\] clknet_4_4_0_clk_regs sg13g2_dfrbpq_1
X_175_ data\[14\] data\[15\] net24 _022_ VPWR VGND sg13g2_mux2_1
XFILLER_35_7 VPWR VGND sg13g2_decap_4
XFILLER_43_207 VPWR VGND sg13g2_fill_1
XFILLER_37_793 VPWR VGND sg13g2_decap_8
XFILLER_25_922 VPWR VGND sg13g2_decap_8
XFILLER_25_999 VPWR VGND sg13g2_decap_8
XFILLER_22_55 VPWR VGND sg13g2_fill_1
XFILLER_22_44 VPWR VGND sg13g2_decap_8
XFILLER_22_33 VPWR VGND sg13g2_fill_1
XFILLER_28_793 VPWR VGND sg13g2_decap_8
XFILLER_43_741 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
X_227_ data\[66\] data\[67\] net26 _074_ VPWR VGND sg13g2_mux2_1
X_158_ _114_ _115_ _005_ VPWR VGND sg13g2_nor2_1
XFILLER_19_793 VPWR VGND sg13g2_decap_8
XFILLER_25_1020 VPWR VGND sg13g2_decap_8
XFILLER_44_505 VPWR VGND sg13g2_fill_1
XFILLER_17_55 VPWR VGND sg13g2_fill_1
XFILLER_48_833 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_39_800 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_1_604 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_clk clknet_1_1__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_5_47 VPWR VGND sg13g2_decap_8
XFILLER_5_36 VPWR VGND sg13g2_fill_1
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_36_814 VPWR VGND sg13g2_decap_8
XFILLER_48_630 VPWR VGND sg13g2_decap_8
XFILLER_0_692 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_42_817 VPWR VGND sg13g2_decap_8
XFILLER_27_814 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_18_814 VPWR VGND sg13g2_decap_8
XFILLER_26_891 VPWR VGND sg13g2_decap_8
XFILLER_33_828 VPWR VGND sg13g2_decap_8
XFILLER_45_666 VPWR VGND sg13g2_decap_8
XFILLER_24_828 VPWR VGND sg13g2_decap_8
XFILLER_24_839 VPWR VGND sg13g2_fill_1
XFILLER_42_603 VPWR VGND sg13g2_decap_8
X_260_ net35 VGND VPWR _020_ data\[13\] clknet_4_8_0_clk_regs sg13g2_dfrbpq_1
XFILLER_25_11 VPWR VGND sg13g2_decap_8
X_191_ data\[30\] data\[31\] net16 _038_ VPWR VGND sg13g2_mux2_1
XFILLER_2_765 VPWR VGND sg13g2_decap_8
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_45_452 VPWR VGND sg13g2_decap_8
XFILLER_20_842 VPWR VGND sg13g2_decap_4
XFILLER_47_728 VPWR VGND sg13g2_decap_8
XFILLER_46_227 VPWR VGND sg13g2_decap_8
X_312_ net29 VGND VPWR _072_ data\[65\] clknet_4_0_0_clk_regs sg13g2_dfrbpq_1
XFILLER_11_842 VPWR VGND sg13g2_decap_4
X_243_ net32 VGND VPWR _003_ u_shift_reg.bit_count\[3\] clknet_4_5_0_clk_regs sg13g2_dfrbpq_1
X_174_ data\[13\] data\[14\] net20 _021_ VPWR VGND sg13g2_mux2_1
XFILLER_46_794 VPWR VGND sg13g2_decap_8
XFILLER_37_772 VPWR VGND sg13g2_decap_8
XFILLER_25_901 VPWR VGND sg13g2_decap_8
XFILLER_25_978 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_28_772 VPWR VGND sg13g2_decap_8
XFILLER_43_720 VPWR VGND sg13g2_decap_8
XFILLER_43_797 VPWR VGND sg13g2_decap_8
XFILLER_8_47 VPWR VGND sg13g2_decap_8
X_226_ data\[65\] data\[66\] net26 _073_ VPWR VGND sg13g2_mux2_1
X_157_ u_shift_reg.bit_count\[5\] _112_ _115_ VPWR VGND sg13g2_nor2_1
XFILLER_19_772 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
XFILLER_34_786 VPWR VGND sg13g2_decap_8
XFILLER_46_591 VPWR VGND sg13g2_decap_8
XFILLER_44_539 VPWR VGND sg13g2_decap_8
XFILLER_25_786 VPWR VGND sg13g2_decap_8
XFILLER_33_55 VPWR VGND sg13g2_fill_1
XFILLER_3_123 VPWR VGND sg13g2_decap_4
XFILLER_48_812 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_43_594 VPWR VGND sg13g2_decap_8
XFILLER_47_399 VPWR VGND sg13g2_decap_8
X_209_ data\[48\] data\[49\] net14 _056_ VPWR VGND sg13g2_mux2_1
XFILLER_39_845 VPWR VGND sg13g2_fill_1
XFILLER_3_690 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_28_22 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_45_848 VPWR VGND sg13g2_fill_2
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_44_98 VPWR VGND sg13g2_decap_8
XFILLER_0_671 VPWR VGND sg13g2_decap_8
XFILLER_48_686 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_8_793 VPWR VGND sg13g2_decap_8
XFILLER_14_24 VPWR VGND sg13g2_decap_4
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_39_54 VPWR VGND sg13g2_fill_2
XFILLER_33_807 VPWR VGND sg13g2_decap_8
XFILLER_45_645 VPWR VGND sg13g2_decap_8
XFILLER_44_133 VPWR VGND sg13g2_decap_8
XFILLER_26_870 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
XFILLER_24_807 VPWR VGND sg13g2_decap_8
XFILLER_46_409 VPWR VGND sg13g2_decap_8
XFILLER_42_659 VPWR VGND sg13g2_decap_8
X_190_ data\[29\] data\[30\] net16 _037_ VPWR VGND sg13g2_mux2_1
XFILLER_41_11 VPWR VGND sg13g2_fill_2
XFILLER_1_221 VPWR VGND sg13g2_fill_2
XFILLER_1_243 VPWR VGND sg13g2_fill_1
XFILLER_2_744 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_45_431 VPWR VGND sg13g2_decap_8
XFILLER_49_781 VPWR VGND sg13g2_decap_8
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_20_821 VPWR VGND sg13g2_decap_8
XFILLER_47_707 VPWR VGND sg13g2_decap_8
XFILLER_46_206 VPWR VGND sg13g2_decap_8
X_311_ net28 VGND VPWR _071_ data\[64\] clknet_4_3_0_clk_regs sg13g2_dfrbpq_1
X_173_ data\[12\] data\[13\] net19 _020_ VPWR VGND sg13g2_mux2_1
XFILLER_7_814 VPWR VGND sg13g2_decap_8
XFILLER_11_821 VPWR VGND sg13g2_decap_8
X_242_ net32 VGND VPWR _002_ u_shift_reg.bit_count\[2\] clknet_4_5_0_clk_regs sg13g2_dfrbpq_1
XFILLER_2_541 VPWR VGND sg13g2_fill_2
XFILLER_28_8 VPWR VGND sg13g2_decap_8
XFILLER_46_773 VPWR VGND sg13g2_decap_8
XFILLER_45_294 VPWR VGND sg13g2_decap_8
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_25_957 VPWR VGND sg13g2_decap_8
XFILLER_3_327 VPWR VGND sg13g2_decap_4
XFILLER_3_305 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
XFILLER_43_776 VPWR VGND sg13g2_decap_8
XFILLER_42_242 VPWR VGND sg13g2_decap_8
XFILLER_42_275 VPWR VGND sg13g2_fill_1
XFILLER_42_286 VPWR VGND sg13g2_decap_8
XFILLER_42_297 VPWR VGND sg13g2_fill_2
X_225_ data\[64\] data\[65\] net15 _072_ VPWR VGND sg13g2_mux2_1
X_156_ _088_ net17 _111_ _114_ VPWR VGND sg13g2_nor3_1
XFILLER_2_393 VPWR VGND sg13g2_decap_4
XFILLER_46_570 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_fill_2
XFILLER_34_765 VPWR VGND sg13g2_decap_8
XFILLER_17_24 VPWR VGND sg13g2_decap_8
XFILLER_25_765 VPWR VGND sg13g2_decap_8
XFILLER_40_779 VPWR VGND sg13g2_decap_8
XFILLER_3_102 VPWR VGND sg13g2_decap_8
XFILLER_3_168 VPWR VGND sg13g2_fill_1
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_31_779 VPWR VGND sg13g2_decap_8
XFILLER_43_573 VPWR VGND sg13g2_decap_8
XFILLER_16_765 VPWR VGND sg13g2_decap_8
X_208_ data\[47\] data\[48\] net15 _055_ VPWR VGND sg13g2_mux2_1
X_139_ _099_ _100_ u_shift_reg.bit_count\[6\] _102_ VPWR VGND _101_ sg13g2_nand4_1
XFILLER_39_824 VPWR VGND sg13g2_decap_8
XFILLER_22_779 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_1_639 VPWR VGND sg13g2_decap_8
XFILLER_45_827 VPWR VGND sg13g2_decap_8
XFILLER_44_326 VPWR VGND sg13g2_decap_4
XFILLER_13_779 VPWR VGND sg13g2_decap_8
XFILLER_44_77 VPWR VGND sg13g2_decap_8
XFILLER_21_790 VPWR VGND sg13g2_decap_8
XFILLER_0_650 VPWR VGND sg13g2_decap_8
XFILLER_36_849 VPWR VGND sg13g2_decap_8
XFILLER_48_665 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
XFILLER_8_772 VPWR VGND sg13g2_decap_8
XFILLER_27_849 VPWR VGND sg13g2_decap_8
Xclkbuf_4_1_0_clk_regs clknet_0_clk_regs clknet_4_1_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_39_33 VPWR VGND sg13g2_decap_8
XFILLER_45_624 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_5_786 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
XFILLER_0_491 VPWR VGND sg13g2_decap_8
XFILLER_42_638 VPWR VGND sg13g2_decap_8
XFILLER_41_45 VPWR VGND sg13g2_decap_8
XFILLER_2_723 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_45_410 VPWR VGND sg13g2_decap_8
XFILLER_45_487 VPWR VGND sg13g2_decap_8
XFILLER_49_4 VPWR VGND sg13g2_decap_8
XFILLER_49_760 VPWR VGND sg13g2_decap_8
XFILLER_20_800 VPWR VGND sg13g2_decap_8
XFILLER_11_26 VPWR VGND sg13g2_decap_8
XFILLER_3_509 VPWR VGND sg13g2_decap_8
X_310_ net28 VGND VPWR _070_ data\[63\] clknet_4_3_0_clk_regs sg13g2_dfrbpq_1
XFILLER_11_800 VPWR VGND sg13g2_decap_8
XFILLER_42_413 VPWR VGND sg13g2_fill_2
X_241_ net32 VGND VPWR _001_ u_shift_reg.bit_count\[1\] clknet_4_4_0_clk_regs sg13g2_dfrbpq_1
X_172_ data\[11\] data\[12\] net22 _019_ VPWR VGND sg13g2_mux2_1
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_597 VPWR VGND sg13g2_decap_8
XFILLER_46_752 VPWR VGND sg13g2_decap_8
XFILLER_45_273 VPWR VGND sg13g2_decap_8
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_25_936 VPWR VGND sg13g2_decap_8
XFILLER_4_807 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_43_755 VPWR VGND sg13g2_decap_8
X_224_ data\[63\] data\[64\] net14 _071_ VPWR VGND sg13g2_mux2_1
XFILLER_8_16 VPWR VGND sg13g2_decap_8
X_155_ _112_ _113_ _004_ VPWR VGND sg13g2_nor2_1
Xclkbuf_4_14_0_clk_regs clknet_0_clk_regs clknet_4_14_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_33_46 VPWR VGND sg13g2_decap_8
XFILLER_0_832 VPWR VGND sg13g2_decap_8
XFILLER_48_847 VPWR VGND sg13g2_decap_8
XFILLER_43_552 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_decap_8
X_207_ data\[46\] data\[47\] net15 _054_ VPWR VGND sg13g2_mux2_1
X_138_ u_shift_reg.bit_count\[2\] u_shift_reg.bit_count\[3\] _101_ VPWR VGND sg13g2_and2_1
XFILLER_1_618 VPWR VGND sg13g2_decap_8
XFILLER_45_806 VPWR VGND sg13g2_decap_8
XFILLER_44_305 VPWR VGND sg13g2_decap_8
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_36_828 VPWR VGND sg13g2_decap_8
XFILLER_48_644 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_27_828 VPWR VGND sg13g2_decap_8
XFILLER_45_603 VPWR VGND sg13g2_decap_8
XFILLER_1_459 VPWR VGND sg13g2_fill_2
XFILLER_18_828 VPWR VGND sg13g2_fill_2
XFILLER_5_765 VPWR VGND sg13g2_decap_8
XFILLER_48_441 VPWR VGND sg13g2_decap_8
XFILLER_32_842 VPWR VGND sg13g2_decap_8
XFILLER_42_617 VPWR VGND sg13g2_decap_8
XFILLER_15_809 VPWR VGND sg13g2_decap_8
XFILLER_23_842 VPWR VGND sg13g2_decap_4
XFILLER_41_24 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_702 VPWR VGND sg13g2_decap_8
XFILLER_2_779 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_45_466 VPWR VGND sg13g2_decap_8
XFILLER_1_790 VPWR VGND sg13g2_decap_8
X_240_ net31 VGND VPWR _000_ u_shift_reg.bit_count\[0\] clknet_4_4_0_clk_regs sg13g2_dfrbpq_1
XFILLER_42_425 VPWR VGND sg13g2_decap_8
XFILLER_42_436 VPWR VGND sg13g2_fill_1
X_171_ data\[10\] data\[11\] net21 _018_ VPWR VGND sg13g2_mux2_1
XFILLER_46_731 VPWR VGND sg13g2_decap_8
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_37_786 VPWR VGND sg13g2_decap_8
XFILLER_25_915 VPWR VGND sg13g2_decap_8
XFILLER_28_786 VPWR VGND sg13g2_decap_8
XFILLER_43_734 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
X_223_ data\[62\] data\[63\] net14 _070_ VPWR VGND sg13g2_mux2_1
XFILLER_3_830 VPWR VGND sg13g2_decap_8
X_154_ u_shift_reg.bit_count\[4\] _110_ _113_ VPWR VGND sg13g2_nor2_1
XFILLER_2_362 VPWR VGND sg13g2_decap_4
XFILLER_19_6 VPWR VGND sg13g2_fill_1
XFILLER_19_786 VPWR VGND sg13g2_decap_8
XFILLER_25_1013 VPWR VGND sg13g2_decap_8
XFILLER_17_48 VPWR VGND sg13g2_decap_8
XFILLER_48_826 VPWR VGND sg13g2_decap_8
XFILLER_0_811 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_decap_8
X_206_ data\[45\] data\[46\] net17 _053_ VPWR VGND sg13g2_mux2_1
X_137_ u_shift_reg.bit_count\[0\] u_shift_reg.bit_count\[1\] _100_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_36_807 VPWR VGND sg13g2_decap_8
XFILLER_48_623 VPWR VGND sg13g2_decap_8
XFILLER_0_685 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_27_807 VPWR VGND sg13g2_decap_8
XFILLER_15_0 VPWR VGND sg13g2_fill_2
XFILLER_18_807 VPWR VGND sg13g2_decap_8
XFILLER_26_884 VPWR VGND sg13g2_decap_8
XFILLER_41_821 VPWR VGND sg13g2_decap_8
XFILLER_45_659 VPWR VGND sg13g2_decap_8
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_17_840 VPWR VGND sg13g2_decap_8
XFILLER_32_821 VPWR VGND sg13g2_decap_8
XFILLER_23_821 VPWR VGND sg13g2_decap_8
XFILLER_2_758 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_45_445 VPWR VGND sg13g2_decap_8
XFILLER_49_795 VPWR VGND sg13g2_decap_8
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_20_846 VPWR VGND sg13g2_fill_2
XFILLER_20_835 VPWR VGND sg13g2_decap_8
XFILLER_11_846 VPWR VGND sg13g2_fill_2
XFILLER_11_835 VPWR VGND sg13g2_decap_8
X_170_ data\[9\] data\[10\] net21 _017_ VPWR VGND sg13g2_mux2_1
XFILLER_46_710 VPWR VGND sg13g2_decap_8
XFILLER_46_787 VPWR VGND sg13g2_decap_8
XFILLER_45_231 VPWR VGND sg13g2_decap_8
X_299_ net28 VGND VPWR _059_ data\[52\] clknet_4_0_0_clk_regs sg13g2_dfrbpq_1
XFILLER_37_765 VPWR VGND sg13g2_decap_8
XFILLER_49_592 VPWR VGND sg13g2_decap_8
XFILLER_3_95 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_28_765 VPWR VGND sg13g2_decap_8
XFILLER_43_713 VPWR VGND sg13g2_decap_8
X_222_ data\[61\] data\[62\] net14 _069_ VPWR VGND sg13g2_mux2_1
X_153_ u_shift_reg.bit_count\[4\] _097_ _101_ _105_ _112_ VPWR VGND sg13g2_and4_1
XFILLER_42_256 VPWR VGND sg13g2_fill_2
XFILLER_19_765 VPWR VGND sg13g2_decap_8
XFILLER_34_779 VPWR VGND sg13g2_decap_8
XFILLER_46_584 VPWR VGND sg13g2_decap_8
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_25_779 VPWR VGND sg13g2_decap_8
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_48_805 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_43_587 VPWR VGND sg13g2_decap_8
XFILLER_16_779 VPWR VGND sg13g2_fill_1
X_136_ u_shift_reg.bit_count\[4\] u_shift_reg.bit_count\[5\] _099_ VPWR VGND sg13g2_nor2_1
X_205_ data\[44\] data\[45\] net18 _052_ VPWR VGND sg13g2_mux2_1
XFILLER_2_193 VPWR VGND sg13g2_decap_8
XFILLER_3_683 VPWR VGND sg13g2_decap_8
XFILLER_39_838 VPWR VGND sg13g2_decap_8
XFILLER_17_4 VPWR VGND sg13g2_fill_2
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_46_381 VPWR VGND sg13g2_decap_8
XFILLER_30_793 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_28_15 VPWR VGND sg13g2_decap_8
XFILLER_38_860 VPWR VGND sg13g2_fill_2
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_48_602 VPWR VGND sg13g2_decap_8
XFILLER_0_664 VPWR VGND sg13g2_decap_8
XFILLER_29_860 VPWR VGND sg13g2_fill_2
XFILLER_48_679 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
X_119_ adc_data\[0\] _089_ net6 VPWR VGND sg13g2_and2_1
XFILLER_8_786 VPWR VGND sg13g2_decap_8
XFILLER_12_793 VPWR VGND sg13g2_decap_8
XFILLER_14_17 VPWR VGND sg13g2_decap_8
XFILLER_14_28 VPWR VGND sg13g2_fill_1
XFILLER_39_47 VPWR VGND sg13g2_decap_8
XFILLER_45_638 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_41_800 VPWR VGND sg13g2_decap_8
XFILLER_26_863 VPWR VGND sg13g2_decap_8
XFILLER_0_472 VPWR VGND sg13g2_decap_8
XFILLER_32_800 VPWR VGND sg13g2_decap_8
XFILLER_44_693 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_23_800 VPWR VGND sg13g2_decap_8
XFILLER_1_214 VPWR VGND sg13g2_decap_8
XFILLER_2_737 VPWR VGND sg13g2_decap_8
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_14_800 VPWR VGND sg13g2_decap_8
XFILLER_45_424 VPWR VGND sg13g2_decap_8
XFILLER_49_774 VPWR VGND sg13g2_decap_8
XFILLER_0_291 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_20_814 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_clk_regs clknet_0_clk_regs clknet_4_0_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_7_807 VPWR VGND sg13g2_decap_8
XFILLER_11_814 VPWR VGND sg13g2_decap_8
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_46_766 VPWR VGND sg13g2_decap_8
XFILLER_45_287 VPWR VGND sg13g2_decap_8
X_298_ net28 VGND VPWR _058_ data\[51\] clknet_4_0_0_clk_regs sg13g2_dfrbpq_1
XFILLER_3_74 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_43_769 VPWR VGND sg13g2_decap_8
XFILLER_42_213 VPWR VGND sg13g2_fill_2
XFILLER_42_268 VPWR VGND sg13g2_decap_8
X_221_ data\[60\] data\[61\] net15 _068_ VPWR VGND sg13g2_mux2_1
X_152_ _101_ _105_ u_shift_reg.bit_count\[4\] _111_ VPWR VGND sg13g2_nand3_1
XFILLER_2_397 VPWR VGND sg13g2_fill_2
XFILLER_2_331 VPWR VGND sg13g2_decap_4
XFILLER_2_320 VPWR VGND sg13g2_decap_8
XFILLER_46_563 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_4
XFILLER_17_17 VPWR VGND sg13g2_decap_8
XFILLER_0_846 VPWR VGND sg13g2_fill_2
XFILLER_43_566 VPWR VGND sg13g2_decap_8
X_204_ data\[43\] data\[44\] net18 _051_ VPWR VGND sg13g2_mux2_1
X_135_ _098_ net2 u_shift_reg.locked VPWR VGND sg13g2_nand2b_1
XFILLER_3_662 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_fill_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_46_360 VPWR VGND sg13g2_decap_8
XFILLER_30_772 VPWR VGND sg13g2_decap_8
XFILLER_44_319 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_clk_regs clknet_0_clk_regs clknet_4_13_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_0_643 VPWR VGND sg13g2_decap_8
XFILLER_48_658 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_8_765 VPWR VGND sg13g2_decap_8
XFILLER_12_772 VPWR VGND sg13g2_decap_8
X_118_ net5 net4 _089_ VPWR VGND sg13g2_nor2b_1
XFILLER_3_470 VPWR VGND sg13g2_fill_2
XFILLER_26_842 VPWR VGND sg13g2_decap_8
XFILLER_45_617 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_5_779 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_32_856 VPWR VGND sg13g2_decap_4
XFILLER_44_672 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XFILLER_43_193 VPWR VGND sg13g2_decap_8
XANTENNA_1 VPWR VGND data\[65\] sg13g2_antennanp
XFILLER_41_38 VPWR VGND sg13g2_decap_8
XFILLER_2_716 VPWR VGND sg13g2_decap_8
XFILLER_45_403 VPWR VGND sg13g2_decap_8
Xheichips25_template_50 VPWR VGND uo_out[0] sg13g2_tielo
XFILLER_49_753 VPWR VGND sg13g2_decap_8
XFILLER_0_270 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_44_491 VPWR VGND sg13g2_decap_8
XFILLER_11_19 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_decap_8
XFILLER_46_745 VPWR VGND sg13g2_decap_8
XFILLER_45_266 VPWR VGND sg13g2_decap_8
X_297_ net28 VGND VPWR _057_ data\[50\] clknet_4_3_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_550 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_1_590 VPWR VGND sg13g2_decap_8
XFILLER_25_929 VPWR VGND sg13g2_decap_8
XFILLER_22_29 VPWR VGND sg13g2_decap_4
XFILLER_43_748 VPWR VGND sg13g2_decap_8
X_220_ data\[59\] data\[60\] net16 _067_ VPWR VGND sg13g2_mux2_1
X_151_ VGND VPWR _087_ _108_ _003_ _110_ sg13g2_a21oi_1
XFILLER_3_844 VPWR VGND sg13g2_decap_4
XFILLER_46_542 VPWR VGND sg13g2_decap_8
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
XFILLER_43_545 VPWR VGND sg13g2_decap_8
X_203_ data\[42\] data\[43\] net17 _050_ VPWR VGND sg13g2_mux2_1
XFILLER_3_641 VPWR VGND sg13g2_decap_8
X_134_ u_shift_reg.locked net2 _097_ VPWR VGND sg13g2_nor2b_1
XFILLER_47_840 VPWR VGND sg13g2_decap_8
XFILLER_39_807 VPWR VGND sg13g2_fill_1
XFILLER_17_6 VPWR VGND sg13g2_fill_1
XFILLER_2_151 VPWR VGND sg13g2_decap_8
XFILLER_31_8 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_48_637 VPWR VGND sg13g2_decap_8
XFILLER_0_622 VPWR VGND sg13g2_decap_8
XFILLER_0_699 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
X_117_ VPWR _088_ u_shift_reg.bit_count\[5\] VGND sg13g2_inv_1
XFILLER_3_482 VPWR VGND sg13g2_decap_8
XFILLER_35_821 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_fill_2
XFILLER_26_898 VPWR VGND sg13g2_decap_8
XFILLER_26_821 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_32_835 VPWR VGND sg13g2_decap_8
XFILLER_44_651 VPWR VGND sg13g2_decap_8
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_fill_1
XFILLER_23_835 VPWR VGND sg13g2_decap_8
XFILLER_23_846 VPWR VGND sg13g2_fill_2
XFILLER_41_17 VPWR VGND sg13g2_decap_8
Xheichips25_template_51 VPWR VGND uo_out[1] sg13g2_tielo
XFILLER_15_51 VPWR VGND sg13g2_decap_4
XFILLER_45_459 VPWR VGND sg13g2_decap_8
XFILLER_49_732 VPWR VGND sg13g2_decap_8
XFILLER_1_783 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_44_470 VPWR VGND sg13g2_decap_8
XFILLER_27_982 VPWR VGND sg13g2_decap_8
XFILLER_46_724 VPWR VGND sg13g2_decap_8
XFILLER_45_245 VPWR VGND sg13g2_decap_8
X_296_ net28 VGND VPWR _056_ data\[49\] clknet_4_0_0_clk_regs sg13g2_dfrbpq_1
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_37_779 VPWR VGND sg13g2_decap_8
XFILLER_25_908 VPWR VGND sg13g2_decap_8
XFILLER_28_779 VPWR VGND sg13g2_decap_8
XFILLER_43_727 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
X_150_ u_shift_reg.bit_count\[0\] u_shift_reg.bit_count\[1\] _097_ _101_ _110_ VPWR
+ VGND sg13g2_and4_1
XFILLER_3_823 VPWR VGND sg13g2_decap_8
XFILLER_46_598 VPWR VGND sg13g2_decap_8
XFILLER_46_521 VPWR VGND sg13g2_decap_8
XFILLER_19_779 VPWR VGND sg13g2_decap_8
XFILLER_42_782 VPWR VGND sg13g2_decap_8
X_279_ net34 VGND VPWR _039_ data\[32\] clknet_4_8_0_clk_regs sg13g2_dfrbpq_1
XFILLER_25_1006 VPWR VGND sg13g2_decap_8
XFILLER_33_793 VPWR VGND sg13g2_decap_8
XFILLER_48_819 VPWR VGND sg13g2_decap_8
XFILLER_0_804 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
X_133_ net13 _095_ _096_ VPWR VGND sg13g2_nand2_1
XFILLER_24_793 VPWR VGND sg13g2_decap_8
X_202_ data\[41\] data\[42\] net17 _049_ VPWR VGND sg13g2_mux2_1
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_3_620 VPWR VGND sg13g2_decap_8
XFILLER_3_697 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_15_793 VPWR VGND sg13g2_decap_4
XFILLER_46_395 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_44_28 VPWR VGND sg13g2_decap_8
XFILLER_0_601 VPWR VGND sg13g2_decap_8
XFILLER_48_616 VPWR VGND sg13g2_decap_8
XFILLER_0_678 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_44_833 VPWR VGND sg13g2_fill_2
XFILLER_43_354 VPWR VGND sg13g2_decap_8
X_116_ VPWR _087_ u_shift_reg.bit_count\[3\] VGND sg13g2_inv_1
XFILLER_35_800 VPWR VGND sg13g2_decap_8
XFILLER_47_693 VPWR VGND sg13g2_decap_8
XFILLER_46_192 VPWR VGND sg13g2_decap_8
XFILLER_30_19 VPWR VGND sg13g2_decap_4
XFILLER_26_877 VPWR VGND sg13g2_decap_8
XFILLER_41_814 VPWR VGND sg13g2_decap_8
XFILLER_26_800 VPWR VGND sg13g2_decap_8
XFILLER_0_442 VPWR VGND sg13g2_decap_8
XFILLER_0_453 VPWR VGND sg13g2_fill_2
XFILLER_44_630 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_17_833 VPWR VGND sg13g2_decap_8
XFILLER_32_814 VPWR VGND sg13g2_decap_8
XFILLER_23_814 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
Xheichips25_template_52 VPWR VGND uo_out[2] sg13g2_tielo
XFILLER_45_438 VPWR VGND sg13g2_decap_8
XFILLER_14_814 VPWR VGND sg13g2_decap_8
XFILLER_49_711 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_49_788 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_20_828 VPWR VGND sg13g2_decap_8
XFILLER_11_828 VPWR VGND sg13g2_decap_8
XFILLER_2_537 VPWR VGND sg13g2_decap_4
Xdelaybuf_0_clk delaynet_0_clk clk VPWR VGND sg13g2_buf_16
XFILLER_27_961 VPWR VGND sg13g2_decap_8
XFILLER_46_703 VPWR VGND sg13g2_decap_8
XFILLER_45_224 VPWR VGND sg13g2_decap_8
X_295_ net29 VGND VPWR _055_ data\[48\] clknet_4_2_0_clk_regs sg13g2_dfrbpq_1
XFILLER_6_821 VPWR VGND sg13g2_decap_8
XFILLER_42_83 VPWR VGND sg13g2_fill_2
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_49_585 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_43_706 VPWR VGND sg13g2_decap_8
XFILLER_42_249 VPWR VGND sg13g2_decap_8
XFILLER_3_802 VPWR VGND sg13g2_decap_8
XFILLER_46_500 VPWR VGND sg13g2_decap_8
XFILLER_42_761 VPWR VGND sg13g2_decap_8
XFILLER_46_577 VPWR VGND sg13g2_decap_8
X_278_ net30 VGND VPWR _038_ data\[31\] clknet_4_2_0_clk_regs sg13g2_dfrbpq_1
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_33_772 VPWR VGND sg13g2_decap_8
XFILLER_3_109 VPWR VGND sg13g2_decap_8
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_24_772 VPWR VGND sg13g2_decap_8
X_201_ data\[40\] data\[41\] net17 _048_ VPWR VGND sg13g2_mux2_1
X_132_ _096_ _090_ clk0_out _089_ adc_data\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_3_676 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_46_374 VPWR VGND sg13g2_decap_8
XFILLER_15_772 VPWR VGND sg13g2_decap_8
XFILLER_30_786 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_fill_1
XFILLER_38_842 VPWR VGND sg13g2_decap_8
XFILLER_21_797 VPWR VGND sg13g2_decap_8
XFILLER_44_812 VPWR VGND sg13g2_decap_8
XFILLER_29_842 VPWR VGND sg13g2_decap_8
XFILLER_0_657 VPWR VGND sg13g2_decap_8
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_34_51 VPWR VGND sg13g2_decap_4
XFILLER_8_779 VPWR VGND sg13g2_decap_8
XFILLER_12_786 VPWR VGND sg13g2_decap_8
XFILLER_47_672 VPWR VGND sg13g2_decap_8
XFILLER_46_171 VPWR VGND sg13g2_decap_8
XFILLER_44_119 VPWR VGND sg13g2_decap_8
XFILLER_26_856 VPWR VGND sg13g2_decap_8
XFILLER_0_465 VPWR VGND sg13g2_decap_8
XFILLER_0_498 VPWR VGND sg13g2_decap_8
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_17_812 VPWR VGND sg13g2_decap_8
XFILLER_44_686 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_4_793 VPWR VGND sg13g2_decap_8
Xclkbuf_4_12_0_clk_regs clknet_0_clk_regs clknet_4_12_0_clk_regs VPWR VGND sg13g2_buf_8
Xheichips25_template_53 VPWR VGND uo_out[3] sg13g2_tielo
XFILLER_45_417 VPWR VGND sg13g2_decap_8
Xoutput6 net6 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_31_41 VPWR VGND sg13g2_decap_8
XFILLER_49_767 VPWR VGND sg13g2_decap_8
XFILLER_0_284 VPWR VGND sg13g2_decap_8
XFILLER_1_730 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_20_807 VPWR VGND sg13g2_decap_8
XFILLER_44_450 VPWR VGND sg13g2_decap_8
.ends

