module heichips25_template (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire \adc_data[0] ;
 wire \adc_data[1] ;
 wire \adc_data[2] ;
 wire \adc_data[3] ;
 wire \adc_data[4] ;
 wire \adc_data[5] ;
 wire \adc_data[6] ;
 wire \adc_data[7] ;
 wire adc_ready;
 wire clk0_out;
 wire clk1_out;
 wire clk2_out;
 wire clk_delayed;
 wire \data[0] ;
 wire \data[10] ;
 wire \data[11] ;
 wire \data[12] ;
 wire \data[13] ;
 wire \data[14] ;
 wire \data[15] ;
 wire \data[16] ;
 wire \data[17] ;
 wire \data[18] ;
 wire \data[19] ;
 wire \data[1] ;
 wire \data[20] ;
 wire \data[21] ;
 wire \data[22] ;
 wire \data[23] ;
 wire \data[24] ;
 wire \data[25] ;
 wire \data[26] ;
 wire \data[27] ;
 wire \data[28] ;
 wire \data[29] ;
 wire \data[2] ;
 wire \data[30] ;
 wire \data[31] ;
 wire \data[32] ;
 wire \data[33] ;
 wire \data[34] ;
 wire \data[35] ;
 wire \data[36] ;
 wire \data[37] ;
 wire \data[38] ;
 wire \data[39] ;
 wire \data[3] ;
 wire \data[40] ;
 wire \data[41] ;
 wire \data[42] ;
 wire \data[43] ;
 wire \data[44] ;
 wire \data[45] ;
 wire \data[46] ;
 wire \data[47] ;
 wire \data[48] ;
 wire \data[49] ;
 wire \data[4] ;
 wire \data[50] ;
 wire \data[51] ;
 wire \data[52] ;
 wire \data[53] ;
 wire \data[54] ;
 wire \data[55] ;
 wire \data[56] ;
 wire \data[57] ;
 wire \data[58] ;
 wire \data[59] ;
 wire \data[5] ;
 wire \data[60] ;
 wire \data[61] ;
 wire \data[62] ;
 wire \data[63] ;
 wire \data[64] ;
 wire \data[65] ;
 wire \data[66] ;
 wire \data[67] ;
 wire \data[68] ;
 wire \data[69] ;
 wire \data[6] ;
 wire \data[70] ;
 wire \data[71] ;
 wire \data[72] ;
 wire \data[73] ;
 wire \data[74] ;
 wire \data[75] ;
 wire \data[76] ;
 wire \data[77] ;
 wire \data[78] ;
 wire \data[7] ;
 wire \data[8] ;
 wire \data[9] ;
 wire osc_out;
 wire net1;
 wire stable;
 wire \u_shift_reg.bit_count[0] ;
 wire \u_shift_reg.bit_count[1] ;
 wire \u_shift_reg.bit_count[2] ;
 wire \u_shift_reg.bit_count[3] ;
 wire \u_shift_reg.bit_count[4] ;
 wire \u_shift_reg.bit_count[5] ;
 wire \u_shift_reg.bit_count[6] ;
 wire \u_shift_reg.locked ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire clk_regs;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;

 sg13g2_inv_1 _116_ (.Y(_087_),
    .A(\u_shift_reg.bit_count[3] ));
 sg13g2_inv_1 _117_ (.Y(_088_),
    .A(\u_shift_reg.bit_count[5] ));
 sg13g2_nor2b_1 _118_ (.A(net5),
    .B_N(net4),
    .Y(_089_));
 sg13g2_and2_1 _119_ (.A(\adc_data[0] ),
    .B(_089_),
    .X(net6));
 sg13g2_and2_1 _120_ (.A(\adc_data[1] ),
    .B(_089_),
    .X(net7));
 sg13g2_and2_1 _121_ (.A(\adc_data[2] ),
    .B(_089_),
    .X(net8));
 sg13g2_nor2_1 _122_ (.A(net5),
    .B(net4),
    .Y(_090_));
 sg13g2_a22oi_1 _123_ (.Y(_091_),
    .B1(_090_),
    .B2(stable),
    .A2(_089_),
    .A1(\adc_data[3] ));
 sg13g2_inv_1 _124_ (.Y(net9),
    .A(_091_));
 sg13g2_a22oi_1 _125_ (.Y(_092_),
    .B1(_090_),
    .B2(osc_out),
    .A2(_089_),
    .A1(\adc_data[4] ));
 sg13g2_inv_1 _126_ (.Y(net10),
    .A(_092_));
 sg13g2_a22oi_1 _127_ (.Y(_093_),
    .B1(_090_),
    .B2(clk2_out),
    .A2(_089_),
    .A1(\adc_data[5] ));
 sg13g2_inv_1 _128_ (.Y(net11),
    .A(_093_));
 sg13g2_a22oi_1 _129_ (.Y(_094_),
    .B1(_090_),
    .B2(clk1_out),
    .A2(_089_),
    .A1(\adc_data[6] ));
 sg13g2_inv_1 _130_ (.Y(net12),
    .A(_094_));
 sg13g2_nand3b_1 _131_ (.B(clk_delayed),
    .C(net5),
    .Y(_095_),
    .A_N(net4));
 sg13g2_a22oi_1 _132_ (.Y(_096_),
    .B1(_090_),
    .B2(clk0_out),
    .A2(_089_),
    .A1(\adc_data[7] ));
 sg13g2_nand2_1 _133_ (.Y(net13),
    .A(_095_),
    .B(_096_));
 sg13g2_nor2b_1 _134_ (.A(\u_shift_reg.locked ),
    .B_N(net2),
    .Y(_097_));
 sg13g2_nand2b_1 _135_ (.Y(_098_),
    .B(net2),
    .A_N(\u_shift_reg.locked ));
 sg13g2_nor2_1 _136_ (.A(\u_shift_reg.bit_count[4] ),
    .B(\u_shift_reg.bit_count[5] ),
    .Y(_099_));
 sg13g2_nor2b_1 _137_ (.A(\u_shift_reg.bit_count[0] ),
    .B_N(\u_shift_reg.bit_count[1] ),
    .Y(_100_));
 sg13g2_and2_1 _138_ (.A(\u_shift_reg.bit_count[2] ),
    .B(\u_shift_reg.bit_count[3] ),
    .X(_101_));
 sg13g2_nand4_1 _139_ (.B(_099_),
    .C(_100_),
    .A(\u_shift_reg.bit_count[6] ),
    .Y(_102_),
    .D(_101_));
 sg13g2_inv_1 _140_ (.Y(_103_),
    .A(_102_));
 sg13g2_a21oi_1 _141_ (.A1(_097_),
    .A2(_102_),
    .Y(_104_),
    .B1(\u_shift_reg.bit_count[0] ));
 sg13g2_a21oi_1 _142_ (.A1(\u_shift_reg.bit_count[0] ),
    .A2(_097_),
    .Y(_000_),
    .B1(_104_));
 sg13g2_and2_1 _143_ (.A(\u_shift_reg.bit_count[0] ),
    .B(\u_shift_reg.bit_count[1] ),
    .X(_105_));
 sg13g2_and3_1 _144_ (.X(_106_),
    .A(\u_shift_reg.bit_count[0] ),
    .B(\u_shift_reg.bit_count[1] ),
    .C(_097_));
 sg13g2_a21oi_1 _145_ (.A1(\u_shift_reg.bit_count[0] ),
    .A2(_097_),
    .Y(_107_),
    .B1(\u_shift_reg.bit_count[1] ));
 sg13g2_nor2_1 _146_ (.A(_106_),
    .B(_107_),
    .Y(_001_));
 sg13g2_nand4_1 _147_ (.B(\u_shift_reg.bit_count[1] ),
    .C(\u_shift_reg.bit_count[2] ),
    .A(\u_shift_reg.bit_count[0] ),
    .Y(_108_),
    .D(_097_));
 sg13g2_o21ai_1 _148_ (.B1(_108_),
    .Y(_109_),
    .A1(\u_shift_reg.bit_count[2] ),
    .A2(_106_));
 sg13g2_inv_1 _149_ (.Y(_002_),
    .A(_109_));
 sg13g2_and4_1 _150_ (.A(\u_shift_reg.bit_count[0] ),
    .B(\u_shift_reg.bit_count[1] ),
    .C(_097_),
    .D(_101_),
    .X(_110_));
 sg13g2_a21oi_1 _151_ (.A1(_087_),
    .A2(_108_),
    .Y(_003_),
    .B1(_110_));
 sg13g2_nand3_1 _152_ (.B(_101_),
    .C(_105_),
    .A(\u_shift_reg.bit_count[4] ),
    .Y(_111_));
 sg13g2_and4_1 _153_ (.A(\u_shift_reg.bit_count[4] ),
    .B(_097_),
    .C(_101_),
    .D(_105_),
    .X(_112_));
 sg13g2_nor2_1 _154_ (.A(\u_shift_reg.bit_count[4] ),
    .B(_110_),
    .Y(_113_));
 sg13g2_nor2_1 _155_ (.A(_112_),
    .B(_113_),
    .Y(_004_));
 sg13g2_nor3_1 _156_ (.A(_088_),
    .B(net17),
    .C(_111_),
    .Y(_114_));
 sg13g2_nor2_1 _157_ (.A(\u_shift_reg.bit_count[5] ),
    .B(_112_),
    .Y(_115_));
 sg13g2_nor2_1 _158_ (.A(_114_),
    .B(_115_),
    .Y(_005_));
 sg13g2_xor2_1 _159_ (.B(_114_),
    .A(\u_shift_reg.bit_count[6] ),
    .X(_006_));
 sg13g2_mux2_1 _160_ (.A0(\data[0] ),
    .A1(net3),
    .S(_097_),
    .X(_007_));
 sg13g2_mux2_1 _161_ (.A0(\data[0] ),
    .A1(\data[1] ),
    .S(net21),
    .X(_008_));
 sg13g2_mux2_1 _162_ (.A0(\data[1] ),
    .A1(\data[2] ),
    .S(net21),
    .X(_009_));
 sg13g2_mux2_1 _163_ (.A0(\data[2] ),
    .A1(\data[3] ),
    .S(net21),
    .X(_010_));
 sg13g2_mux2_1 _164_ (.A0(\data[3] ),
    .A1(\data[4] ),
    .S(net21),
    .X(_011_));
 sg13g2_mux2_1 _165_ (.A0(\data[4] ),
    .A1(\data[5] ),
    .S(net21),
    .X(_012_));
 sg13g2_mux2_1 _166_ (.A0(\data[5] ),
    .A1(\data[6] ),
    .S(net25),
    .X(_013_));
 sg13g2_mux2_1 _167_ (.A0(\data[6] ),
    .A1(\data[7] ),
    .S(net25),
    .X(_014_));
 sg13g2_mux2_1 _168_ (.A0(\data[7] ),
    .A1(\data[8] ),
    .S(net25),
    .X(_015_));
 sg13g2_mux2_1 _169_ (.A0(\data[8] ),
    .A1(\data[9] ),
    .S(net25),
    .X(_016_));
 sg13g2_mux2_1 _170_ (.A0(\data[9] ),
    .A1(\data[10] ),
    .S(net21),
    .X(_017_));
 sg13g2_mux2_1 _171_ (.A0(\data[10] ),
    .A1(\data[11] ),
    .S(net21),
    .X(_018_));
 sg13g2_mux2_1 _172_ (.A0(\data[11] ),
    .A1(\data[12] ),
    .S(net22),
    .X(_019_));
 sg13g2_mux2_1 _173_ (.A0(\data[12] ),
    .A1(\data[13] ),
    .S(net19),
    .X(_020_));
 sg13g2_mux2_1 _174_ (.A0(\data[13] ),
    .A1(\data[14] ),
    .S(net20),
    .X(_021_));
 sg13g2_mux2_1 _175_ (.A0(\data[14] ),
    .A1(\data[15] ),
    .S(net24),
    .X(_022_));
 sg13g2_mux2_1 _176_ (.A0(\data[15] ),
    .A1(\data[16] ),
    .S(net24),
    .X(_023_));
 sg13g2_mux2_1 _177_ (.A0(\data[16] ),
    .A1(\data[17] ),
    .S(net24),
    .X(_024_));
 sg13g2_mux2_1 _178_ (.A0(\data[17] ),
    .A1(\data[18] ),
    .S(net24),
    .X(_025_));
 sg13g2_mux2_1 _179_ (.A0(\data[18] ),
    .A1(\data[19] ),
    .S(net25),
    .X(_026_));
 sg13g2_mux2_1 _180_ (.A0(\data[19] ),
    .A1(\data[20] ),
    .S(net24),
    .X(_027_));
 sg13g2_mux2_1 _181_ (.A0(\data[20] ),
    .A1(\data[21] ),
    .S(net24),
    .X(_028_));
 sg13g2_mux2_1 _182_ (.A0(\data[21] ),
    .A1(\data[22] ),
    .S(net24),
    .X(_029_));
 sg13g2_mux2_1 _183_ (.A0(\data[22] ),
    .A1(\data[23] ),
    .S(net20),
    .X(_030_));
 sg13g2_mux2_1 _184_ (.A0(\data[23] ),
    .A1(\data[24] ),
    .S(net20),
    .X(_031_));
 sg13g2_mux2_1 _185_ (.A0(\data[24] ),
    .A1(\data[25] ),
    .S(net20),
    .X(_032_));
 sg13g2_mux2_1 _186_ (.A0(\data[25] ),
    .A1(\data[26] ),
    .S(net20),
    .X(_033_));
 sg13g2_mux2_1 _187_ (.A0(\data[26] ),
    .A1(\data[27] ),
    .S(net19),
    .X(_034_));
 sg13g2_mux2_1 _188_ (.A0(\data[27] ),
    .A1(\data[28] ),
    .S(net19),
    .X(_035_));
 sg13g2_mux2_1 _189_ (.A0(\data[28] ),
    .A1(\data[29] ),
    .S(net19),
    .X(_036_));
 sg13g2_mux2_1 _190_ (.A0(\data[29] ),
    .A1(\data[30] ),
    .S(net16),
    .X(_037_));
 sg13g2_mux2_1 _191_ (.A0(\data[30] ),
    .A1(\data[31] ),
    .S(net16),
    .X(_038_));
 sg13g2_mux2_1 _192_ (.A0(\data[31] ),
    .A1(\data[32] ),
    .S(net19),
    .X(_039_));
 sg13g2_mux2_1 _193_ (.A0(\data[32] ),
    .A1(\data[33] ),
    .S(net19),
    .X(_040_));
 sg13g2_mux2_1 _194_ (.A0(\data[33] ),
    .A1(\data[34] ),
    .S(net19),
    .X(_041_));
 sg13g2_mux2_1 _195_ (.A0(\data[34] ),
    .A1(\data[35] ),
    .S(net19),
    .X(_042_));
 sg13g2_mux2_1 _196_ (.A0(\data[35] ),
    .A1(\data[36] ),
    .S(net20),
    .X(_043_));
 sg13g2_mux2_1 _197_ (.A0(\data[36] ),
    .A1(\data[37] ),
    .S(net20),
    .X(_044_));
 sg13g2_mux2_1 _198_ (.A0(\data[37] ),
    .A1(\data[38] ),
    .S(net24),
    .X(_045_));
 sg13g2_mux2_1 _199_ (.A0(\data[38] ),
    .A1(\data[39] ),
    .S(net14),
    .X(_046_));
 sg13g2_mux2_1 _200_ (.A0(\data[39] ),
    .A1(\data[40] ),
    .S(net17),
    .X(_047_));
 sg13g2_mux2_1 _201_ (.A0(\data[40] ),
    .A1(\data[41] ),
    .S(net17),
    .X(_048_));
 sg13g2_mux2_1 _202_ (.A0(\data[41] ),
    .A1(\data[42] ),
    .S(net17),
    .X(_049_));
 sg13g2_mux2_1 _203_ (.A0(\data[42] ),
    .A1(\data[43] ),
    .S(net17),
    .X(_050_));
 sg13g2_mux2_1 _204_ (.A0(\data[43] ),
    .A1(\data[44] ),
    .S(net18),
    .X(_051_));
 sg13g2_mux2_1 _205_ (.A0(\data[44] ),
    .A1(\data[45] ),
    .S(net18),
    .X(_052_));
 sg13g2_mux2_1 _206_ (.A0(\data[45] ),
    .A1(\data[46] ),
    .S(net17),
    .X(_053_));
 sg13g2_mux2_1 _207_ (.A0(\data[46] ),
    .A1(\data[47] ),
    .S(net15),
    .X(_054_));
 sg13g2_mux2_1 _208_ (.A0(\data[47] ),
    .A1(\data[48] ),
    .S(net15),
    .X(_055_));
 sg13g2_mux2_1 _209_ (.A0(\data[48] ),
    .A1(\data[49] ),
    .S(net14),
    .X(_056_));
 sg13g2_mux2_1 _210_ (.A0(\data[49] ),
    .A1(\data[50] ),
    .S(net14),
    .X(_057_));
 sg13g2_mux2_1 _211_ (.A0(\data[50] ),
    .A1(\data[51] ),
    .S(net14),
    .X(_058_));
 sg13g2_mux2_1 _212_ (.A0(\data[51] ),
    .A1(\data[52] ),
    .S(net14),
    .X(_059_));
 sg13g2_mux2_1 _213_ (.A0(\data[52] ),
    .A1(\data[53] ),
    .S(net15),
    .X(_060_));
 sg13g2_mux2_1 _214_ (.A0(\data[53] ),
    .A1(\data[54] ),
    .S(net17),
    .X(_061_));
 sg13g2_mux2_1 _215_ (.A0(\data[54] ),
    .A1(\data[55] ),
    .S(net17),
    .X(_062_));
 sg13g2_mux2_1 _216_ (.A0(\data[55] ),
    .A1(\data[56] ),
    .S(net18),
    .X(_063_));
 sg13g2_mux2_1 _217_ (.A0(\data[56] ),
    .A1(\data[57] ),
    .S(net18),
    .X(_064_));
 sg13g2_mux2_1 _218_ (.A0(\data[57] ),
    .A1(\data[58] ),
    .S(net21),
    .X(_065_));
 sg13g2_mux2_1 _219_ (.A0(\data[58] ),
    .A1(\data[59] ),
    .S(net16),
    .X(_066_));
 sg13g2_mux2_1 _220_ (.A0(\data[59] ),
    .A1(\data[60] ),
    .S(net16),
    .X(_067_));
 sg13g2_mux2_1 _221_ (.A0(\data[60] ),
    .A1(\data[61] ),
    .S(net15),
    .X(_068_));
 sg13g2_mux2_1 _222_ (.A0(\data[61] ),
    .A1(\data[62] ),
    .S(net14),
    .X(_069_));
 sg13g2_mux2_1 _223_ (.A0(\data[62] ),
    .A1(\data[63] ),
    .S(net14),
    .X(_070_));
 sg13g2_mux2_1 _224_ (.A0(\data[63] ),
    .A1(\data[64] ),
    .S(net14),
    .X(_071_));
 sg13g2_mux2_1 _225_ (.A0(\data[64] ),
    .A1(\data[65] ),
    .S(net15),
    .X(_072_));
 sg13g2_mux2_1 _226_ (.A0(\data[65] ),
    .A1(\data[66] ),
    .S(net26),
    .X(_073_));
 sg13g2_mux2_1 _227_ (.A0(\data[66] ),
    .A1(\data[67] ),
    .S(net26),
    .X(_074_));
 sg13g2_mux2_1 _228_ (.A0(\data[67] ),
    .A1(\data[68] ),
    .S(net26),
    .X(_075_));
 sg13g2_mux2_1 _229_ (.A0(\data[68] ),
    .A1(\data[69] ),
    .S(net26),
    .X(_076_));
 sg13g2_mux2_1 _230_ (.A0(\data[69] ),
    .A1(\data[70] ),
    .S(net26),
    .X(_077_));
 sg13g2_mux2_1 _231_ (.A0(\data[70] ),
    .A1(\data[71] ),
    .S(net26),
    .X(_078_));
 sg13g2_mux2_1 _232_ (.A0(\data[71] ),
    .A1(\data[72] ),
    .S(net26),
    .X(_079_));
 sg13g2_mux2_1 _233_ (.A0(\data[72] ),
    .A1(\data[73] ),
    .S(net26),
    .X(_080_));
 sg13g2_mux2_1 _234_ (.A0(\data[73] ),
    .A1(\data[74] ),
    .S(net27),
    .X(_081_));
 sg13g2_mux2_1 _235_ (.A0(\data[74] ),
    .A1(\data[75] ),
    .S(net27),
    .X(_082_));
 sg13g2_mux2_1 _236_ (.A0(\data[75] ),
    .A1(\data[76] ),
    .S(net27),
    .X(_083_));
 sg13g2_mux2_1 _237_ (.A0(\data[76] ),
    .A1(\data[77] ),
    .S(net27),
    .X(_084_));
 sg13g2_mux2_1 _238_ (.A0(\data[77] ),
    .A1(\data[78] ),
    .S(net27),
    .X(_085_));
 sg13g2_a21o_1 _239_ (.A2(_103_),
    .A1(net2),
    .B1(\u_shift_reg.locked ),
    .X(_086_));
 sg13g2_dfrbpq_1 _240_ (.RESET_B(net31),
    .D(_000_),
    .Q(\u_shift_reg.bit_count[0] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _241_ (.RESET_B(net32),
    .D(_001_),
    .Q(\u_shift_reg.bit_count[1] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _242_ (.RESET_B(net32),
    .D(_002_),
    .Q(\u_shift_reg.bit_count[2] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _243_ (.RESET_B(net32),
    .D(_003_),
    .Q(\u_shift_reg.bit_count[3] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _244_ (.RESET_B(net32),
    .D(_004_),
    .Q(\u_shift_reg.bit_count[4] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _245_ (.RESET_B(net31),
    .D(_005_),
    .Q(\u_shift_reg.bit_count[5] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _246_ (.RESET_B(net31),
    .D(_006_),
    .Q(\u_shift_reg.bit_count[6] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _247_ (.RESET_B(net32),
    .D(_007_),
    .Q(\data[0] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _248_ (.RESET_B(net36),
    .D(_008_),
    .Q(\data[1] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _249_ (.RESET_B(net36),
    .D(_009_),
    .Q(\data[2] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _250_ (.RESET_B(net36),
    .D(_010_),
    .Q(\data[3] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _251_ (.RESET_B(net36),
    .D(_011_),
    .Q(\data[4] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _252_ (.RESET_B(net39),
    .D(_012_),
    .Q(\data[5] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _253_ (.RESET_B(net39),
    .D(_013_),
    .Q(\data[6] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _254_ (.RESET_B(net39),
    .D(_014_),
    .Q(\data[7] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _255_ (.RESET_B(net39),
    .D(_015_),
    .Q(\data[8] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _256_ (.RESET_B(net39),
    .D(_016_),
    .Q(\data[9] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _257_ (.RESET_B(net36),
    .D(_017_),
    .Q(\data[10] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _258_ (.RESET_B(net36),
    .D(_018_),
    .Q(\data[11] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _259_ (.RESET_B(net37),
    .D(_019_),
    .Q(\data[12] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _260_ (.RESET_B(net35),
    .D(_020_),
    .Q(\data[13] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _261_ (.RESET_B(net35),
    .D(_021_),
    .Q(\data[14] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _262_ (.RESET_B(net38),
    .D(_022_),
    .Q(\data[15] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _263_ (.RESET_B(net38),
    .D(_023_),
    .Q(\data[16] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _264_ (.RESET_B(net38),
    .D(_024_),
    .Q(\data[17] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _265_ (.RESET_B(net39),
    .D(_025_),
    .Q(\data[18] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _266_ (.RESET_B(net39),
    .D(_026_),
    .Q(\data[19] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _267_ (.RESET_B(net38),
    .D(_027_),
    .Q(\data[20] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _268_ (.RESET_B(net38),
    .D(_028_),
    .Q(\data[21] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _269_ (.RESET_B(net38),
    .D(_029_),
    .Q(\data[22] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _270_ (.RESET_B(net35),
    .D(_030_),
    .Q(\data[23] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _271_ (.RESET_B(net35),
    .D(_031_),
    .Q(\data[24] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _272_ (.RESET_B(net35),
    .D(_032_),
    .Q(\data[25] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _273_ (.RESET_B(net35),
    .D(_033_),
    .Q(\data[26] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _274_ (.RESET_B(net34),
    .D(_034_),
    .Q(\data[27] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _275_ (.RESET_B(net34),
    .D(_035_),
    .Q(\data[28] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _276_ (.RESET_B(net34),
    .D(_036_),
    .Q(\data[29] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _277_ (.RESET_B(net30),
    .D(_037_),
    .Q(\data[30] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _278_ (.RESET_B(net30),
    .D(_038_),
    .Q(\data[31] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _279_ (.RESET_B(net34),
    .D(_039_),
    .Q(\data[32] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _280_ (.RESET_B(net34),
    .D(_040_),
    .Q(\data[33] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _281_ (.RESET_B(net34),
    .D(_041_),
    .Q(\data[34] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _282_ (.RESET_B(net34),
    .D(_042_),
    .Q(\data[35] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _283_ (.RESET_B(net35),
    .D(_043_),
    .Q(\data[36] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _284_ (.RESET_B(net38),
    .D(_044_),
    .Q(\data[37] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _285_ (.RESET_B(net38),
    .D(_045_),
    .Q(\data[38] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _286_ (.RESET_B(net28),
    .D(_046_),
    .Q(\data[39] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _287_ (.RESET_B(net31),
    .D(_047_),
    .Q(\data[40] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _288_ (.RESET_B(net31),
    .D(_048_),
    .Q(\data[41] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _289_ (.RESET_B(net32),
    .D(_049_),
    .Q(\data[42] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _290_ (.RESET_B(net33),
    .D(_050_),
    .Q(\data[43] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _291_ (.RESET_B(net33),
    .D(_051_),
    .Q(\data[44] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _292_ (.RESET_B(net33),
    .D(_052_),
    .Q(\data[45] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _293_ (.RESET_B(net31),
    .D(_053_),
    .Q(\data[46] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _294_ (.RESET_B(net29),
    .D(_054_),
    .Q(\data[47] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _295_ (.RESET_B(net29),
    .D(_055_),
    .Q(\data[48] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _296_ (.RESET_B(net28),
    .D(_056_),
    .Q(\data[49] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _297_ (.RESET_B(net28),
    .D(_057_),
    .Q(\data[50] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _298_ (.RESET_B(net28),
    .D(_058_),
    .Q(\data[51] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _299_ (.RESET_B(net28),
    .D(_059_),
    .Q(\data[52] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _300_ (.RESET_B(net31),
    .D(_060_),
    .Q(\data[53] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _301_ (.RESET_B(net31),
    .D(_061_),
    .Q(\data[54] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _302_ (.RESET_B(net33),
    .D(_062_),
    .Q(\data[55] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _303_ (.RESET_B(net33),
    .D(_063_),
    .Q(\data[56] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _304_ (.RESET_B(net36),
    .D(_064_),
    .Q(\data[57] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _305_ (.RESET_B(net36),
    .D(_065_),
    .Q(\data[58] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _306_ (.RESET_B(net30),
    .D(_066_),
    .Q(\data[59] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _307_ (.RESET_B(net30),
    .D(_067_),
    .Q(\data[60] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _308_ (.RESET_B(net29),
    .D(_068_),
    .Q(\data[61] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _309_ (.RESET_B(net28),
    .D(_069_),
    .Q(\data[62] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _310_ (.RESET_B(net28),
    .D(_070_),
    .Q(\data[63] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _311_ (.RESET_B(net28),
    .D(_071_),
    .Q(\data[64] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _312_ (.RESET_B(net29),
    .D(_072_),
    .Q(\data[65] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _313_ (.RESET_B(net40),
    .D(_073_),
    .Q(\data[66] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _314_ (.RESET_B(net40),
    .D(_074_),
    .Q(\data[67] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _315_ (.RESET_B(net40),
    .D(_075_),
    .Q(\data[68] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _316_ (.RESET_B(net40),
    .D(_076_),
    .Q(\data[69] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _317_ (.RESET_B(net40),
    .D(_077_),
    .Q(\data[70] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _318_ (.RESET_B(net40),
    .D(_078_),
    .Q(\data[71] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _319_ (.RESET_B(net40),
    .D(_079_),
    .Q(\data[72] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _320_ (.RESET_B(net40),
    .D(_080_),
    .Q(\data[73] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _321_ (.RESET_B(net41),
    .D(_081_),
    .Q(\data[74] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _322_ (.RESET_B(net41),
    .D(_082_),
    .Q(\data[75] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _323_ (.RESET_B(net41),
    .D(_083_),
    .Q(\data[76] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _324_ (.RESET_B(net41),
    .D(_084_),
    .Q(\data[77] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _325_ (.RESET_B(net41),
    .D(_085_),
    .Q(\data[78] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _326_ (.RESET_B(net32),
    .D(_086_),
    .Q(\u_shift_reg.locked ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_tielo heichips25_template_43 (.L_LO(net43));
 sg13g2_tielo heichips25_template_44 (.L_LO(net44));
 sg13g2_tielo heichips25_template_45 (.L_LO(net45));
 sg13g2_tielo heichips25_template_46 (.L_LO(net46));
 sg13g2_tielo heichips25_template_47 (.L_LO(net47));
 sg13g2_tielo heichips25_template_48 (.L_LO(net48));
 sg13g2_tielo heichips25_template_49 (.L_LO(net49));
 sg13g2_tielo heichips25_template_50 (.L_LO(net50));
 sg13g2_tielo heichips25_template_51 (.L_LO(net51));
 sg13g2_tielo heichips25_template_52 (.L_LO(net52));
 sg13g2_tielo heichips25_template_53 (.L_LO(net53));
 sg13g2_tielo heichips25_template_54 (.L_LO(net54));
 sg13g2_tielo heichips25_template_55 (.L_LO(net55));
 sg13g2_tielo heichips25_template_56 (.L_LO(net56));
 sg13g2_tielo heichips25_template_57 (.L_LO(net57));
 sg13g2_buf_16 clkbuf_regs_0_clk (.X(clk_regs),
    .A(clk));
 adc u_adc (.clk(clknet_1_0__leaf_clk),
    .ready(adc_ready),
    .start(\data[66] ),
    .analog_in({\data[74] ,
    \data[73] ,
    \data[72] ,
    \data[71] ,
    \data[70] ,
    \data[69] ,
    \data[68] ,
    \data[67] }),
    .data_out({\adc_data[7] ,
    \adc_data[6] ,
    \adc_data[5] ,
    \adc_data[4] ,
    \adc_data[3] ,
    \adc_data[2] ,
    \adc_data[1] ,
    \adc_data[0] }));
 delay_line u_delay_line (.clk(clknet_1_1__leaf_clk),
    .clk_delayed(clk_delayed),
    .delay({\data[78] ,
    \data[77] ,
    \data[76] ,
    \data[75] }));
 multimode_dll u_multimode_dll (.bias(\data[38] ),
    .clk0_out(clk0_out),
    .clk1_out(clk1_out),
    .clk2_out(clk2_out),
    .dco(\data[39] ),
    .enable(ena),
    .osc(clknet_1_0__leaf_clk),
    .osc_out(osc_out),
    .resetb(net34),
    .stable(stable),
    .clk0_phase_sel({\data[24] ,
    \data[23] ,
    \data[22] ,
    \data[21] ,
    \data[20] }),
    .clk1_phase_sel({\data[29] ,
    \data[28] ,
    \data[27] ,
    \data[26] ,
    \data[25] }),
    .clk2_phase_sel({\data[34] ,
    \data[33] ,
    \data[32] ,
    \data[31] ,
    \data[30] }),
    .ext_trim({\data[65] ,
    \data[64] ,
    \data[63] ,
    \data[62] ,
    \data[61] ,
    \data[60] ,
    \data[59] ,
    \data[58] ,
    \data[57] ,
    \data[56] ,
    \data[55] ,
    \data[54] ,
    \data[53] ,
    \data[52] ,
    \data[51] ,
    \data[50] ,
    \data[49] ,
    \data[48] ,
    \data[47] ,
    \data[46] ,
    \data[45] ,
    \data[44] ,
    \data[43] ,
    \data[42] ,
    \data[41] ,
    \data[40] }),
    .f_clk0_divider({\data[9] ,
    \data[8] ,
    \data[7] ,
    \data[6] ,
    \data[5] }),
    .f_clk1_divider({\data[14] ,
    \data[13] ,
    \data[12] ,
    \data[11] ,
    \data[10] }),
    .f_clk2_divider({\data[19] ,
    \data[18] ,
    \data[17] ,
    \data[16] ,
    \data[15] }),
    .f_osc_multiply_factor({\data[4] ,
    \data[3] ,
    \data[2] ,
    \data[1] ,
    \data[0] }),
    .mode_xor({\data[37] ,
    \data[36] ,
    \data[35] }));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[7]));
 sg13g2_buf_1 fanout14 (.A(net15),
    .X(net14));
 sg13g2_buf_1 fanout15 (.A(net16),
    .X(net15));
 sg13g2_buf_1 fanout16 (.A(net23),
    .X(net16));
 sg13g2_buf_1 fanout17 (.A(net23),
    .X(net17));
 sg13g2_buf_1 fanout18 (.A(net23),
    .X(net18));
 sg13g2_buf_1 fanout19 (.A(net22),
    .X(net19));
 sg13g2_buf_1 fanout20 (.A(net22),
    .X(net20));
 sg13g2_buf_1 fanout21 (.A(net22),
    .X(net21));
 sg13g2_buf_1 fanout22 (.A(net23),
    .X(net22));
 sg13g2_buf_1 fanout23 (.A(_098_),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(net25),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(_098_),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(net27),
    .X(net26));
 sg13g2_buf_1 fanout27 (.A(_098_),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(net29),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(net30),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(net42),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net33),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(net42),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(net37),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net37),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(net37),
    .X(net36));
 sg13g2_buf_1 fanout37 (.A(net42),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(net39),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(net42),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net42),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(net1),
    .X(net42));
 sg13g2_tielo heichips25_template (.L_LO(net));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(delaynet_0_clk));
 sg13g2_buf_16 clkbuf_1_0__f_clk (.X(clknet_1_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_1_1__f_clk (.X(clknet_1_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_0_clk_regs (.X(clknet_0_clk_regs),
    .A(clk_regs));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_4_14_0_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_4_15_0_clk_regs));
 sg13g2_buf_16 delaybuf_0_clk (.X(delaynet_0_clk),
    .A(clk));
 sg13g2_antennanp ANTENNA_1 (.A(\data[65] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_fill_1 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_fill_1 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_fill_1 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_4 FILLER_0_357 ();
 sg13g2_fill_1 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_4 FILLER_0_379 ();
 sg13g2_fill_2 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_fill_2 FILLER_0_402 ();
 sg13g2_fill_1 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_4 FILLER_0_449 ();
 sg13g2_fill_2 FILLER_0_453 ();
 sg13g2_decap_8 FILLER_0_465 ();
 sg13g2_decap_8 FILLER_0_472 ();
 sg13g2_fill_2 FILLER_0_479 ();
 sg13g2_decap_8 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_498 ();
 sg13g2_decap_4 FILLER_0_505 ();
 sg13g2_decap_8 FILLER_0_519 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_fill_2 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_545 ();
 sg13g2_decap_8 FILLER_0_552 ();
 sg13g2_decap_8 FILLER_0_559 ();
 sg13g2_decap_8 FILLER_0_566 ();
 sg13g2_decap_8 FILLER_0_573 ();
 sg13g2_decap_8 FILLER_0_580 ();
 sg13g2_decap_8 FILLER_0_587 ();
 sg13g2_decap_8 FILLER_0_594 ();
 sg13g2_decap_8 FILLER_0_601 ();
 sg13g2_decap_8 FILLER_0_608 ();
 sg13g2_decap_8 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_636 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_decap_8 FILLER_0_678 ();
 sg13g2_decap_8 FILLER_0_685 ();
 sg13g2_decap_8 FILLER_0_692 ();
 sg13g2_decap_8 FILLER_0_699 ();
 sg13g2_decap_8 FILLER_0_706 ();
 sg13g2_decap_8 FILLER_0_713 ();
 sg13g2_decap_8 FILLER_0_720 ();
 sg13g2_decap_8 FILLER_0_727 ();
 sg13g2_decap_8 FILLER_0_734 ();
 sg13g2_decap_8 FILLER_0_741 ();
 sg13g2_decap_8 FILLER_0_748 ();
 sg13g2_decap_8 FILLER_0_755 ();
 sg13g2_decap_8 FILLER_0_762 ();
 sg13g2_decap_8 FILLER_0_769 ();
 sg13g2_decap_8 FILLER_0_776 ();
 sg13g2_decap_8 FILLER_0_783 ();
 sg13g2_decap_8 FILLER_0_790 ();
 sg13g2_decap_8 FILLER_0_797 ();
 sg13g2_decap_8 FILLER_0_804 ();
 sg13g2_decap_8 FILLER_0_811 ();
 sg13g2_decap_4 FILLER_0_818 ();
 sg13g2_decap_8 FILLER_0_832 ();
 sg13g2_decap_8 FILLER_0_839 ();
 sg13g2_fill_2 FILLER_0_846 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_4 FILLER_1_182 ();
 sg13g2_fill_1 FILLER_1_186 ();
 sg13g2_decap_8 FILLER_1_214 ();
 sg13g2_fill_2 FILLER_1_221 ();
 sg13g2_fill_1 FILLER_1_243 ();
 sg13g2_fill_1 FILLER_1_271 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_fill_2 FILLER_1_316 ();
 sg13g2_fill_1 FILLER_1_355 ();
 sg13g2_fill_2 FILLER_1_383 ();
 sg13g2_fill_1 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_fill_2 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_459 ();
 sg13g2_decap_8 FILLER_1_569 ();
 sg13g2_decap_8 FILLER_1_576 ();
 sg13g2_decap_8 FILLER_1_583 ();
 sg13g2_decap_8 FILLER_1_590 ();
 sg13g2_decap_8 FILLER_1_597 ();
 sg13g2_decap_8 FILLER_1_604 ();
 sg13g2_decap_8 FILLER_1_611 ();
 sg13g2_decap_8 FILLER_1_618 ();
 sg13g2_decap_8 FILLER_1_625 ();
 sg13g2_decap_8 FILLER_1_632 ();
 sg13g2_decap_8 FILLER_1_639 ();
 sg13g2_decap_8 FILLER_1_646 ();
 sg13g2_decap_8 FILLER_1_653 ();
 sg13g2_decap_8 FILLER_1_660 ();
 sg13g2_decap_8 FILLER_1_667 ();
 sg13g2_decap_8 FILLER_1_674 ();
 sg13g2_decap_8 FILLER_1_681 ();
 sg13g2_decap_8 FILLER_1_688 ();
 sg13g2_decap_8 FILLER_1_695 ();
 sg13g2_decap_8 FILLER_1_702 ();
 sg13g2_decap_8 FILLER_1_709 ();
 sg13g2_decap_8 FILLER_1_716 ();
 sg13g2_decap_8 FILLER_1_723 ();
 sg13g2_decap_8 FILLER_1_730 ();
 sg13g2_decap_8 FILLER_1_737 ();
 sg13g2_decap_8 FILLER_1_769 ();
 sg13g2_decap_8 FILLER_1_776 ();
 sg13g2_decap_8 FILLER_1_783 ();
 sg13g2_decap_8 FILLER_1_790 ();
 sg13g2_decap_8 FILLER_1_797 ();
 sg13g2_decap_8 FILLER_1_804 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_4 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_fill_2 FILLER_2_200 ();
 sg13g2_fill_1 FILLER_2_202 ();
 sg13g2_decap_4 FILLER_2_230 ();
 sg13g2_fill_1 FILLER_2_234 ();
 sg13g2_decap_8 FILLER_2_239 ();
 sg13g2_decap_8 FILLER_2_246 ();
 sg13g2_fill_1 FILLER_2_253 ();
 sg13g2_fill_2 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_320 ();
 sg13g2_decap_4 FILLER_2_331 ();
 sg13g2_decap_4 FILLER_2_362 ();
 sg13g2_decap_4 FILLER_2_393 ();
 sg13g2_fill_2 FILLER_2_397 ();
 sg13g2_decap_8 FILLER_2_426 ();
 sg13g2_fill_1 FILLER_2_433 ();
 sg13g2_decap_8 FILLER_2_471 ();
 sg13g2_fill_2 FILLER_2_478 ();
 sg13g2_fill_2 FILLER_2_507 ();
 sg13g2_fill_1 FILLER_2_509 ();
 sg13g2_decap_4 FILLER_2_537 ();
 sg13g2_fill_2 FILLER_2_541 ();
 sg13g2_decap_8 FILLER_2_597 ();
 sg13g2_decap_8 FILLER_2_604 ();
 sg13g2_decap_8 FILLER_2_611 ();
 sg13g2_decap_8 FILLER_2_618 ();
 sg13g2_decap_8 FILLER_2_625 ();
 sg13g2_decap_8 FILLER_2_632 ();
 sg13g2_decap_8 FILLER_2_639 ();
 sg13g2_decap_8 FILLER_2_646 ();
 sg13g2_decap_8 FILLER_2_653 ();
 sg13g2_decap_8 FILLER_2_660 ();
 sg13g2_decap_8 FILLER_2_667 ();
 sg13g2_decap_8 FILLER_2_674 ();
 sg13g2_decap_8 FILLER_2_681 ();
 sg13g2_decap_8 FILLER_2_688 ();
 sg13g2_decap_8 FILLER_2_695 ();
 sg13g2_decap_8 FILLER_2_702 ();
 sg13g2_decap_8 FILLER_2_709 ();
 sg13g2_decap_8 FILLER_2_716 ();
 sg13g2_decap_8 FILLER_2_723 ();
 sg13g2_decap_8 FILLER_2_730 ();
 sg13g2_decap_8 FILLER_2_737 ();
 sg13g2_decap_8 FILLER_2_744 ();
 sg13g2_decap_8 FILLER_2_751 ();
 sg13g2_decap_8 FILLER_2_758 ();
 sg13g2_decap_8 FILLER_2_765 ();
 sg13g2_decap_8 FILLER_2_772 ();
 sg13g2_decap_8 FILLER_2_779 ();
 sg13g2_decap_8 FILLER_2_786 ();
 sg13g2_decap_8 FILLER_2_793 ();
 sg13g2_decap_8 FILLER_2_800 ();
 sg13g2_decap_8 FILLER_2_807 ();
 sg13g2_decap_8 FILLER_2_814 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_4 FILLER_3_123 ();
 sg13g2_decap_4 FILLER_3_164 ();
 sg13g2_fill_1 FILLER_3_168 ();
 sg13g2_decap_4 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_200 ();
 sg13g2_fill_2 FILLER_3_212 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_4 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_320 ();
 sg13g2_decap_4 FILLER_3_327 ();
 sg13g2_fill_2 FILLER_3_331 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_4 FILLER_3_370 ();
 sg13g2_fill_1 FILLER_3_374 ();
 sg13g2_decap_4 FILLER_3_393 ();
 sg13g2_fill_2 FILLER_3_397 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_fill_2 FILLER_3_430 ();
 sg13g2_fill_1 FILLER_3_432 ();
 sg13g2_decap_4 FILLER_3_466 ();
 sg13g2_fill_2 FILLER_3_470 ();
 sg13g2_decap_8 FILLER_3_482 ();
 sg13g2_decap_8 FILLER_3_489 ();
 sg13g2_fill_2 FILLER_3_496 ();
 sg13g2_fill_1 FILLER_3_498 ();
 sg13g2_decap_8 FILLER_3_509 ();
 sg13g2_decap_8 FILLER_3_516 ();
 sg13g2_decap_8 FILLER_3_523 ();
 sg13g2_fill_2 FILLER_3_530 ();
 sg13g2_decap_8 FILLER_3_542 ();
 sg13g2_decap_8 FILLER_3_549 ();
 sg13g2_decap_4 FILLER_3_556 ();
 sg13g2_fill_1 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_571 ();
 sg13g2_decap_8 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_585 ();
 sg13g2_decap_8 FILLER_3_592 ();
 sg13g2_decap_8 FILLER_3_599 ();
 sg13g2_decap_8 FILLER_3_606 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_decap_8 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_648 ();
 sg13g2_decap_8 FILLER_3_655 ();
 sg13g2_decap_8 FILLER_3_662 ();
 sg13g2_decap_8 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_676 ();
 sg13g2_decap_8 FILLER_3_683 ();
 sg13g2_decap_8 FILLER_3_690 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_8 FILLER_3_704 ();
 sg13g2_decap_8 FILLER_3_711 ();
 sg13g2_decap_8 FILLER_3_718 ();
 sg13g2_decap_8 FILLER_3_725 ();
 sg13g2_decap_8 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_8 FILLER_3_746 ();
 sg13g2_decap_8 FILLER_3_753 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_decap_8 FILLER_3_767 ();
 sg13g2_decap_8 FILLER_3_774 ();
 sg13g2_decap_8 FILLER_3_781 ();
 sg13g2_decap_8 FILLER_3_788 ();
 sg13g2_decap_8 FILLER_3_795 ();
 sg13g2_decap_8 FILLER_3_802 ();
 sg13g2_decap_8 FILLER_3_809 ();
 sg13g2_decap_8 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_3_823 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_837 ();
 sg13g2_decap_4 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_fill_2 FILLER_4_53 ();
 sg13g2_fill_1 FILLER_4_55 ();
 sg13g2_decap_8 FILLER_4_765 ();
 sg13g2_decap_8 FILLER_4_772 ();
 sg13g2_decap_8 FILLER_4_779 ();
 sg13g2_decap_8 FILLER_4_786 ();
 sg13g2_decap_8 FILLER_4_793 ();
 sg13g2_decap_8 FILLER_4_800 ();
 sg13g2_decap_8 FILLER_4_807 ();
 sg13g2_decap_8 FILLER_4_814 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_4 FILLER_5_32 ();
 sg13g2_fill_1 FILLER_5_36 ();
 sg13g2_decap_8 FILLER_5_47 ();
 sg13g2_fill_2 FILLER_5_54 ();
 sg13g2_decap_8 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_8 FILLER_5_786 ();
 sg13g2_decap_8 FILLER_5_793 ();
 sg13g2_decap_8 FILLER_5_800 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_decap_4 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_4 FILLER_5_842 ();
 sg13g2_fill_2 FILLER_5_846 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_4 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_765 ();
 sg13g2_decap_8 FILLER_6_772 ();
 sg13g2_decap_8 FILLER_6_779 ();
 sg13g2_decap_8 FILLER_6_786 ();
 sg13g2_decap_8 FILLER_6_793 ();
 sg13g2_decap_8 FILLER_6_800 ();
 sg13g2_decap_8 FILLER_6_807 ();
 sg13g2_decap_8 FILLER_6_814 ();
 sg13g2_decap_8 FILLER_6_821 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_fill_2 FILLER_6_845 ();
 sg13g2_fill_1 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_765 ();
 sg13g2_decap_8 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_779 ();
 sg13g2_decap_8 FILLER_7_786 ();
 sg13g2_decap_8 FILLER_7_793 ();
 sg13g2_decap_8 FILLER_7_800 ();
 sg13g2_decap_8 FILLER_7_807 ();
 sg13g2_decap_8 FILLER_7_814 ();
 sg13g2_fill_2 FILLER_8_4 ();
 sg13g2_fill_1 FILLER_8_6 ();
 sg13g2_decap_8 FILLER_8_16 ();
 sg13g2_decap_8 FILLER_8_23 ();
 sg13g2_decap_8 FILLER_8_40 ();
 sg13g2_decap_8 FILLER_8_47 ();
 sg13g2_fill_2 FILLER_8_54 ();
 sg13g2_decap_8 FILLER_8_765 ();
 sg13g2_decap_8 FILLER_8_772 ();
 sg13g2_decap_8 FILLER_8_779 ();
 sg13g2_decap_8 FILLER_8_786 ();
 sg13g2_decap_8 FILLER_8_793 ();
 sg13g2_decap_8 FILLER_8_800 ();
 sg13g2_decap_8 FILLER_8_807 ();
 sg13g2_decap_8 FILLER_8_814 ();
 sg13g2_decap_8 FILLER_8_821 ();
 sg13g2_decap_8 FILLER_8_828 ();
 sg13g2_decap_8 FILLER_8_835 ();
 sg13g2_decap_4 FILLER_8_842 ();
 sg13g2_fill_2 FILLER_8_846 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_4 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_765 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_8 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_786 ();
 sg13g2_decap_8 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_835 ();
 sg13g2_decap_4 FILLER_9_842 ();
 sg13g2_fill_2 FILLER_9_846 ();
 sg13g2_decap_4 FILLER_10_50 ();
 sg13g2_fill_2 FILLER_10_54 ();
 sg13g2_decap_8 FILLER_10_765 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_4 FILLER_10_842 ();
 sg13g2_fill_2 FILLER_10_846 ();
 sg13g2_decap_8 FILLER_11_19 ();
 sg13g2_decap_8 FILLER_11_26 ();
 sg13g2_fill_2 FILLER_11_33 ();
 sg13g2_decap_8 FILLER_11_45 ();
 sg13g2_decap_4 FILLER_11_52 ();
 sg13g2_decap_8 FILLER_11_765 ();
 sg13g2_decap_8 FILLER_11_772 ();
 sg13g2_decap_8 FILLER_11_779 ();
 sg13g2_decap_8 FILLER_11_786 ();
 sg13g2_decap_8 FILLER_11_793 ();
 sg13g2_decap_8 FILLER_11_800 ();
 sg13g2_decap_8 FILLER_11_807 ();
 sg13g2_decap_8 FILLER_11_814 ();
 sg13g2_decap_8 FILLER_11_821 ();
 sg13g2_decap_8 FILLER_11_828 ();
 sg13g2_decap_8 FILLER_11_835 ();
 sg13g2_decap_4 FILLER_11_842 ();
 sg13g2_fill_2 FILLER_11_846 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_772 ();
 sg13g2_decap_8 FILLER_12_779 ();
 sg13g2_decap_8 FILLER_12_786 ();
 sg13g2_decap_8 FILLER_12_793 ();
 sg13g2_decap_8 FILLER_12_800 ();
 sg13g2_decap_8 FILLER_12_807 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_8 FILLER_13_13 ();
 sg13g2_decap_8 FILLER_13_20 ();
 sg13g2_decap_4 FILLER_13_27 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_772 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_decap_8 FILLER_13_793 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_4 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_835 ();
 sg13g2_decap_4 FILLER_13_842 ();
 sg13g2_fill_2 FILLER_13_846 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_6 ();
 sg13g2_decap_8 FILLER_14_17 ();
 sg13g2_decap_4 FILLER_14_24 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_44 ();
 sg13g2_decap_4 FILLER_15_51 ();
 sg13g2_fill_1 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_8 FILLER_15_772 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_8 FILLER_15_786 ();
 sg13g2_decap_4 FILLER_15_793 ();
 sg13g2_fill_1 FILLER_15_797 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_8 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_4 FILLER_15_843 ();
 sg13g2_fill_1 FILLER_15_847 ();
 sg13g2_decap_4 FILLER_16_4 ();
 sg13g2_fill_1 FILLER_16_8 ();
 sg13g2_decap_8 FILLER_16_16 ();
 sg13g2_decap_4 FILLER_16_23 ();
 sg13g2_fill_2 FILLER_16_27 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_779 ();
 sg13g2_fill_1 FILLER_16_820 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_6 ();
 sg13g2_decap_8 FILLER_17_17 ();
 sg13g2_decap_8 FILLER_17_24 ();
 sg13g2_decap_8 FILLER_17_41 ();
 sg13g2_decap_8 FILLER_17_48 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_decap_8 FILLER_17_765 ();
 sg13g2_decap_8 FILLER_17_772 ();
 sg13g2_decap_8 FILLER_17_779 ();
 sg13g2_fill_1 FILLER_17_786 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_fill_1 FILLER_17_847 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_fill_2 FILLER_18_828 ();
 sg13g2_fill_1 FILLER_18_830 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_6 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_4 FILLER_19_32 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_decap_8 FILLER_19_47 ();
 sg13g2_fill_2 FILLER_19_54 ();
 sg13g2_decap_8 FILLER_19_765 ();
 sg13g2_decap_8 FILLER_19_772 ();
 sg13g2_decap_8 FILLER_19_779 ();
 sg13g2_decap_8 FILLER_19_786 ();
 sg13g2_decap_8 FILLER_19_793 ();
 sg13g2_decap_8 FILLER_19_800 ();
 sg13g2_decap_8 FILLER_19_807 ();
 sg13g2_decap_8 FILLER_19_814 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_decap_4 FILLER_20_24 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_765 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_779 ();
 sg13g2_decap_8 FILLER_20_786 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_8 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_814 ();
 sg13g2_decap_8 FILLER_20_821 ();
 sg13g2_decap_8 FILLER_20_828 ();
 sg13g2_decap_8 FILLER_20_835 ();
 sg13g2_decap_4 FILLER_20_842 ();
 sg13g2_fill_2 FILLER_20_846 ();
 sg13g2_decap_4 FILLER_21_8 ();
 sg13g2_fill_2 FILLER_21_12 ();
 sg13g2_decap_8 FILLER_21_41 ();
 sg13g2_decap_8 FILLER_21_48 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_decap_8 FILLER_21_790 ();
 sg13g2_decap_8 FILLER_21_797 ();
 sg13g2_decap_8 FILLER_21_804 ();
 sg13g2_decap_8 FILLER_21_811 ();
 sg13g2_decap_8 FILLER_21_818 ();
 sg13g2_decap_8 FILLER_21_825 ();
 sg13g2_decap_8 FILLER_21_832 ();
 sg13g2_decap_8 FILLER_21_839 ();
 sg13g2_fill_2 FILLER_21_846 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_20 ();
 sg13g2_decap_4 FILLER_22_29 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_decap_8 FILLER_22_44 ();
 sg13g2_decap_4 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_decap_8 FILLER_22_779 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_793 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_decap_8 FILLER_22_835 ();
 sg13g2_decap_4 FILLER_22_842 ();
 sg13g2_fill_2 FILLER_22_846 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_765 ();
 sg13g2_decap_8 FILLER_23_772 ();
 sg13g2_decap_8 FILLER_23_779 ();
 sg13g2_decap_8 FILLER_23_786 ();
 sg13g2_decap_8 FILLER_23_793 ();
 sg13g2_decap_8 FILLER_23_800 ();
 sg13g2_decap_8 FILLER_23_807 ();
 sg13g2_decap_8 FILLER_23_814 ();
 sg13g2_decap_8 FILLER_23_821 ();
 sg13g2_decap_8 FILLER_23_828 ();
 sg13g2_decap_8 FILLER_23_835 ();
 sg13g2_decap_4 FILLER_23_842 ();
 sg13g2_fill_2 FILLER_23_846 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_17 ();
 sg13g2_decap_8 FILLER_24_24 ();
 sg13g2_decap_8 FILLER_24_31 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_786 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_4 FILLER_24_835 ();
 sg13g2_fill_1 FILLER_24_839 ();
 sg13g2_decap_4 FILLER_24_844 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_fill_1 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_fill_1 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_873 ();
 sg13g2_decap_8 FILLER_25_880 ();
 sg13g2_decap_8 FILLER_25_887 ();
 sg13g2_decap_8 FILLER_25_894 ();
 sg13g2_decap_8 FILLER_25_901 ();
 sg13g2_decap_8 FILLER_25_908 ();
 sg13g2_decap_8 FILLER_25_915 ();
 sg13g2_decap_8 FILLER_25_922 ();
 sg13g2_decap_8 FILLER_25_929 ();
 sg13g2_decap_8 FILLER_25_936 ();
 sg13g2_decap_8 FILLER_25_943 ();
 sg13g2_decap_8 FILLER_25_950 ();
 sg13g2_decap_8 FILLER_25_957 ();
 sg13g2_decap_8 FILLER_25_964 ();
 sg13g2_decap_8 FILLER_25_971 ();
 sg13g2_decap_8 FILLER_25_978 ();
 sg13g2_decap_8 FILLER_25_985 ();
 sg13g2_decap_8 FILLER_25_992 ();
 sg13g2_decap_8 FILLER_25_999 ();
 sg13g2_decap_8 FILLER_25_1006 ();
 sg13g2_decap_8 FILLER_25_1013 ();
 sg13g2_decap_8 FILLER_25_1020 ();
 sg13g2_fill_2 FILLER_25_1027 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_4 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_765 ();
 sg13g2_decap_8 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_779 ();
 sg13g2_decap_8 FILLER_26_786 ();
 sg13g2_decap_8 FILLER_26_793 ();
 sg13g2_decap_8 FILLER_26_800 ();
 sg13g2_decap_8 FILLER_26_807 ();
 sg13g2_decap_8 FILLER_26_814 ();
 sg13g2_decap_8 FILLER_26_821 ();
 sg13g2_decap_8 FILLER_26_828 ();
 sg13g2_decap_8 FILLER_26_835 ();
 sg13g2_decap_8 FILLER_26_842 ();
 sg13g2_decap_8 FILLER_26_849 ();
 sg13g2_decap_8 FILLER_26_856 ();
 sg13g2_decap_8 FILLER_26_863 ();
 sg13g2_decap_8 FILLER_26_870 ();
 sg13g2_decap_8 FILLER_26_877 ();
 sg13g2_decap_8 FILLER_26_884 ();
 sg13g2_decap_8 FILLER_26_891 ();
 sg13g2_decap_8 FILLER_26_898 ();
 sg13g2_decap_8 FILLER_26_905 ();
 sg13g2_decap_8 FILLER_26_912 ();
 sg13g2_decap_8 FILLER_26_919 ();
 sg13g2_decap_8 FILLER_26_926 ();
 sg13g2_decap_8 FILLER_26_933 ();
 sg13g2_decap_8 FILLER_26_940 ();
 sg13g2_decap_8 FILLER_26_947 ();
 sg13g2_decap_8 FILLER_26_954 ();
 sg13g2_decap_8 FILLER_26_961 ();
 sg13g2_decap_8 FILLER_26_968 ();
 sg13g2_decap_8 FILLER_26_975 ();
 sg13g2_decap_8 FILLER_26_982 ();
 sg13g2_decap_8 FILLER_26_989 ();
 sg13g2_decap_8 FILLER_26_996 ();
 sg13g2_decap_8 FILLER_26_1003 ();
 sg13g2_decap_8 FILLER_26_1010 ();
 sg13g2_decap_8 FILLER_26_1017 ();
 sg13g2_decap_4 FILLER_26_1024 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_45 ();
 sg13g2_decap_4 FILLER_27_52 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_decap_8 FILLER_27_772 ();
 sg13g2_decap_8 FILLER_27_779 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_decap_8 FILLER_27_954 ();
 sg13g2_decap_8 FILLER_27_961 ();
 sg13g2_decap_8 FILLER_27_968 ();
 sg13g2_decap_8 FILLER_27_975 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_4 FILLER_27_1024 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_28_8 ();
 sg13g2_decap_8 FILLER_28_15 ();
 sg13g2_decap_8 FILLER_28_22 ();
 sg13g2_decap_8 FILLER_28_765 ();
 sg13g2_decap_8 FILLER_28_772 ();
 sg13g2_decap_8 FILLER_28_779 ();
 sg13g2_decap_8 FILLER_28_786 ();
 sg13g2_decap_8 FILLER_28_793 ();
 sg13g2_decap_8 FILLER_28_800 ();
 sg13g2_decap_8 FILLER_28_807 ();
 sg13g2_decap_8 FILLER_28_814 ();
 sg13g2_decap_8 FILLER_28_821 ();
 sg13g2_decap_8 FILLER_28_828 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_decap_8 FILLER_28_842 ();
 sg13g2_decap_8 FILLER_28_849 ();
 sg13g2_decap_4 FILLER_28_856 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_27 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_decap_8 FILLER_29_45 ();
 sg13g2_decap_4 FILLER_29_52 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_19 ();
 sg13g2_decap_4 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_772 ();
 sg13g2_decap_8 FILLER_30_779 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_4 FILLER_30_856 ();
 sg13g2_fill_2 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_31_8 ();
 sg13g2_decap_8 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_41 ();
 sg13g2_decap_8 FILLER_31_48 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_765 ();
 sg13g2_decap_8 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_786 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_fill_2 FILLER_31_821 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_16 ();
 sg13g2_decap_4 FILLER_32_23 ();
 sg13g2_fill_2 FILLER_32_27 ();
 sg13g2_decap_8 FILLER_32_765 ();
 sg13g2_decap_8 FILLER_32_772 ();
 sg13g2_decap_8 FILLER_32_779 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_decap_8 FILLER_32_793 ();
 sg13g2_decap_8 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_814 ();
 sg13g2_decap_8 FILLER_32_821 ();
 sg13g2_decap_8 FILLER_32_828 ();
 sg13g2_decap_8 FILLER_32_835 ();
 sg13g2_decap_8 FILLER_32_842 ();
 sg13g2_decap_8 FILLER_32_849 ();
 sg13g2_decap_4 FILLER_32_856 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_53 ();
 sg13g2_fill_1 FILLER_33_55 ();
 sg13g2_decap_8 FILLER_33_765 ();
 sg13g2_decap_8 FILLER_33_772 ();
 sg13g2_decap_8 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_decap_8 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_33_828 ();
 sg13g2_decap_8 FILLER_33_835 ();
 sg13g2_decap_8 FILLER_33_842 ();
 sg13g2_decap_8 FILLER_33_849 ();
 sg13g2_decap_4 FILLER_33_856 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_13 ();
 sg13g2_fill_1 FILLER_34_17 ();
 sg13g2_decap_4 FILLER_34_23 ();
 sg13g2_decap_8 FILLER_34_44 ();
 sg13g2_decap_4 FILLER_34_51 ();
 sg13g2_fill_1 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_765 ();
 sg13g2_decap_8 FILLER_34_772 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_8 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_793 ();
 sg13g2_decap_8 FILLER_34_800 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_decap_8 FILLER_34_814 ();
 sg13g2_decap_8 FILLER_34_821 ();
 sg13g2_decap_8 FILLER_34_828 ();
 sg13g2_decap_4 FILLER_34_835 ();
 sg13g2_fill_2 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_851 ();
 sg13g2_decap_4 FILLER_34_858 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_fill_2 FILLER_35_19 ();
 sg13g2_fill_1 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_27 ();
 sg13g2_decap_8 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_772 ();
 sg13g2_decap_8 FILLER_35_779 ();
 sg13g2_decap_8 FILLER_35_786 ();
 sg13g2_decap_8 FILLER_35_793 ();
 sg13g2_decap_8 FILLER_35_800 ();
 sg13g2_decap_8 FILLER_35_807 ();
 sg13g2_decap_8 FILLER_35_814 ();
 sg13g2_decap_8 FILLER_35_821 ();
 sg13g2_decap_8 FILLER_35_828 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_765 ();
 sg13g2_decap_8 FILLER_36_772 ();
 sg13g2_decap_8 FILLER_36_779 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_8 FILLER_36_793 ();
 sg13g2_decap_8 FILLER_36_800 ();
 sg13g2_decap_8 FILLER_36_807 ();
 sg13g2_decap_8 FILLER_36_814 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_decap_8 FILLER_36_828 ();
 sg13g2_decap_8 FILLER_36_835 ();
 sg13g2_decap_8 FILLER_36_842 ();
 sg13g2_decap_8 FILLER_36_849 ();
 sg13g2_decap_4 FILLER_36_856 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_18 ();
 sg13g2_fill_1 FILLER_37_20 ();
 sg13g2_fill_1 FILLER_37_27 ();
 sg13g2_fill_2 FILLER_37_38 ();
 sg13g2_decap_8 FILLER_37_765 ();
 sg13g2_decap_8 FILLER_37_772 ();
 sg13g2_decap_8 FILLER_37_779 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_807 ();
 sg13g2_decap_8 FILLER_37_814 ();
 sg13g2_decap_8 FILLER_37_821 ();
 sg13g2_decap_8 FILLER_37_828 ();
 sg13g2_decap_8 FILLER_37_835 ();
 sg13g2_decap_8 FILLER_37_842 ();
 sg13g2_decap_8 FILLER_37_849 ();
 sg13g2_decap_4 FILLER_37_856 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_decap_4 FILLER_38_23 ();
 sg13g2_fill_2 FILLER_38_27 ();
 sg13g2_decap_8 FILLER_38_765 ();
 sg13g2_decap_8 FILLER_38_772 ();
 sg13g2_decap_8 FILLER_38_779 ();
 sg13g2_decap_8 FILLER_38_786 ();
 sg13g2_decap_8 FILLER_38_793 ();
 sg13g2_decap_8 FILLER_38_800 ();
 sg13g2_decap_8 FILLER_38_807 ();
 sg13g2_decap_8 FILLER_38_814 ();
 sg13g2_decap_8 FILLER_38_821 ();
 sg13g2_decap_8 FILLER_38_828 ();
 sg13g2_decap_8 FILLER_38_835 ();
 sg13g2_decap_8 FILLER_38_842 ();
 sg13g2_decap_8 FILLER_38_849 ();
 sg13g2_decap_4 FILLER_38_856 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_33 ();
 sg13g2_decap_8 FILLER_39_40 ();
 sg13g2_decap_8 FILLER_39_47 ();
 sg13g2_fill_2 FILLER_39_54 ();
 sg13g2_decap_8 FILLER_39_765 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_fill_1 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_824 ();
 sg13g2_decap_8 FILLER_39_831 ();
 sg13g2_decap_8 FILLER_39_838 ();
 sg13g2_fill_1 FILLER_39_845 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_15 ();
 sg13g2_fill_1 FILLER_40_17 ();
 sg13g2_fill_1 FILLER_40_55 ();
 sg13g2_decap_8 FILLER_40_765 ();
 sg13g2_decap_8 FILLER_40_772 ();
 sg13g2_decap_8 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_828 ();
 sg13g2_decap_4 FILLER_40_835 ();
 sg13g2_fill_2 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_11 ();
 sg13g2_decap_8 FILLER_41_17 ();
 sg13g2_decap_8 FILLER_41_24 ();
 sg13g2_decap_8 FILLER_41_31 ();
 sg13g2_decap_8 FILLER_41_38 ();
 sg13g2_decap_8 FILLER_41_45 ();
 sg13g2_decap_4 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_765 ();
 sg13g2_decap_8 FILLER_41_772 ();
 sg13g2_decap_8 FILLER_41_779 ();
 sg13g2_decap_8 FILLER_41_786 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_828 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_76 ();
 sg13g2_fill_2 FILLER_42_83 ();
 sg13g2_fill_1 FILLER_42_95 ();
 sg13g2_decap_8 FILLER_42_123 ();
 sg13g2_decap_4 FILLER_42_130 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_decap_8 FILLER_42_146 ();
 sg13g2_decap_8 FILLER_42_163 ();
 sg13g2_fill_2 FILLER_42_170 ();
 sg13g2_decap_4 FILLER_42_209 ();
 sg13g2_fill_2 FILLER_42_213 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_decap_8 FILLER_42_249 ();
 sg13g2_fill_2 FILLER_42_256 ();
 sg13g2_decap_8 FILLER_42_261 ();
 sg13g2_decap_8 FILLER_42_268 ();
 sg13g2_fill_1 FILLER_42_275 ();
 sg13g2_decap_8 FILLER_42_286 ();
 sg13g2_decap_4 FILLER_42_293 ();
 sg13g2_fill_2 FILLER_42_297 ();
 sg13g2_decap_8 FILLER_42_326 ();
 sg13g2_decap_4 FILLER_42_333 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_fill_2 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_425 ();
 sg13g2_fill_1 FILLER_42_436 ();
 sg13g2_fill_2 FILLER_42_462 ();
 sg13g2_fill_1 FILLER_42_464 ();
 sg13g2_decap_8 FILLER_42_475 ();
 sg13g2_fill_2 FILLER_42_482 ();
 sg13g2_fill_1 FILLER_42_484 ();
 sg13g2_decap_8 FILLER_42_561 ();
 sg13g2_decap_8 FILLER_42_568 ();
 sg13g2_decap_8 FILLER_42_575 ();
 sg13g2_decap_8 FILLER_42_582 ();
 sg13g2_decap_8 FILLER_42_589 ();
 sg13g2_decap_8 FILLER_42_596 ();
 sg13g2_decap_8 FILLER_42_603 ();
 sg13g2_decap_8 FILLER_42_610 ();
 sg13g2_decap_8 FILLER_42_617 ();
 sg13g2_decap_8 FILLER_42_624 ();
 sg13g2_decap_8 FILLER_42_631 ();
 sg13g2_decap_8 FILLER_42_638 ();
 sg13g2_decap_8 FILLER_42_645 ();
 sg13g2_decap_8 FILLER_42_652 ();
 sg13g2_decap_8 FILLER_42_659 ();
 sg13g2_decap_4 FILLER_42_666 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_4 FILLER_42_707 ();
 sg13g2_fill_2 FILLER_42_711 ();
 sg13g2_decap_8 FILLER_42_726 ();
 sg13g2_decap_8 FILLER_42_733 ();
 sg13g2_decap_8 FILLER_42_740 ();
 sg13g2_decap_8 FILLER_42_747 ();
 sg13g2_decap_8 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_decap_8 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_789 ();
 sg13g2_decap_8 FILLER_42_796 ();
 sg13g2_decap_8 FILLER_42_803 ();
 sg13g2_decap_8 FILLER_42_810 ();
 sg13g2_decap_8 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_824 ();
 sg13g2_decap_8 FILLER_42_831 ();
 sg13g2_decap_8 FILLER_42_838 ();
 sg13g2_decap_8 FILLER_42_845 ();
 sg13g2_decap_8 FILLER_42_852 ();
 sg13g2_fill_2 FILLER_42_859 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_4 FILLER_43_133 ();
 sg13g2_fill_2 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_166 ();
 sg13g2_fill_1 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_179 ();
 sg13g2_decap_8 FILLER_43_186 ();
 sg13g2_decap_8 FILLER_43_193 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_fill_1 FILLER_43_207 ();
 sg13g2_fill_1 FILLER_43_231 ();
 sg13g2_decap_4 FILLER_43_272 ();
 sg13g2_decap_4 FILLER_43_303 ();
 sg13g2_decap_8 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_415 ();
 sg13g2_decap_4 FILLER_43_422 ();
 sg13g2_fill_1 FILLER_43_426 ();
 sg13g2_decap_8 FILLER_43_454 ();
 sg13g2_decap_8 FILLER_43_545 ();
 sg13g2_decap_8 FILLER_43_552 ();
 sg13g2_decap_8 FILLER_43_559 ();
 sg13g2_decap_8 FILLER_43_566 ();
 sg13g2_decap_8 FILLER_43_573 ();
 sg13g2_decap_8 FILLER_43_580 ();
 sg13g2_decap_8 FILLER_43_587 ();
 sg13g2_decap_8 FILLER_43_594 ();
 sg13g2_decap_8 FILLER_43_601 ();
 sg13g2_decap_8 FILLER_43_608 ();
 sg13g2_decap_8 FILLER_43_615 ();
 sg13g2_decap_8 FILLER_43_622 ();
 sg13g2_decap_8 FILLER_43_629 ();
 sg13g2_decap_8 FILLER_43_636 ();
 sg13g2_decap_8 FILLER_43_643 ();
 sg13g2_decap_8 FILLER_43_650 ();
 sg13g2_decap_8 FILLER_43_657 ();
 sg13g2_decap_8 FILLER_43_664 ();
 sg13g2_decap_8 FILLER_43_671 ();
 sg13g2_decap_8 FILLER_43_678 ();
 sg13g2_decap_8 FILLER_43_685 ();
 sg13g2_decap_8 FILLER_43_692 ();
 sg13g2_decap_8 FILLER_43_699 ();
 sg13g2_decap_8 FILLER_43_706 ();
 sg13g2_decap_8 FILLER_43_713 ();
 sg13g2_decap_8 FILLER_43_720 ();
 sg13g2_decap_8 FILLER_43_727 ();
 sg13g2_decap_8 FILLER_43_734 ();
 sg13g2_decap_8 FILLER_43_741 ();
 sg13g2_decap_8 FILLER_43_748 ();
 sg13g2_decap_8 FILLER_43_755 ();
 sg13g2_decap_8 FILLER_43_762 ();
 sg13g2_decap_8 FILLER_43_769 ();
 sg13g2_decap_8 FILLER_43_776 ();
 sg13g2_decap_8 FILLER_43_783 ();
 sg13g2_decap_8 FILLER_43_790 ();
 sg13g2_decap_8 FILLER_43_797 ();
 sg13g2_decap_8 FILLER_43_804 ();
 sg13g2_decap_8 FILLER_43_811 ();
 sg13g2_decap_8 FILLER_43_818 ();
 sg13g2_decap_8 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_4 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_853 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_236 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_decap_8 FILLER_44_250 ();
 sg13g2_decap_8 FILLER_44_257 ();
 sg13g2_decap_8 FILLER_44_264 ();
 sg13g2_decap_8 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_decap_8 FILLER_44_285 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_4 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_decap_8 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_44_415 ();
 sg13g2_decap_8 FILLER_44_422 ();
 sg13g2_decap_8 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_44_436 ();
 sg13g2_decap_8 FILLER_44_443 ();
 sg13g2_decap_8 FILLER_44_450 ();
 sg13g2_decap_8 FILLER_44_457 ();
 sg13g2_fill_2 FILLER_44_464 ();
 sg13g2_decap_8 FILLER_44_470 ();
 sg13g2_decap_8 FILLER_44_477 ();
 sg13g2_decap_8 FILLER_44_484 ();
 sg13g2_decap_8 FILLER_44_491 ();
 sg13g2_decap_8 FILLER_44_498 ();
 sg13g2_fill_1 FILLER_44_505 ();
 sg13g2_decap_8 FILLER_44_539 ();
 sg13g2_decap_8 FILLER_44_546 ();
 sg13g2_decap_8 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_8 FILLER_44_567 ();
 sg13g2_decap_8 FILLER_44_574 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_decap_8 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_609 ();
 sg13g2_decap_8 FILLER_44_616 ();
 sg13g2_decap_8 FILLER_44_623 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_decap_8 FILLER_44_637 ();
 sg13g2_decap_8 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_651 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_693 ();
 sg13g2_decap_8 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_714 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_fill_2 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_45_147 ();
 sg13g2_fill_1 FILLER_45_149 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_fill_1 FILLER_45_329 ();
 sg13g2_decap_4 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_354 ();
 sg13g2_decap_8 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_396 ();
 sg13g2_decap_8 FILLER_45_403 ();
 sg13g2_decap_8 FILLER_45_410 ();
 sg13g2_decap_8 FILLER_45_417 ();
 sg13g2_decap_8 FILLER_45_424 ();
 sg13g2_decap_8 FILLER_45_431 ();
 sg13g2_decap_8 FILLER_45_438 ();
 sg13g2_decap_8 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_decap_8 FILLER_45_459 ();
 sg13g2_decap_8 FILLER_45_466 ();
 sg13g2_decap_8 FILLER_45_473 ();
 sg13g2_decap_8 FILLER_45_480 ();
 sg13g2_decap_8 FILLER_45_487 ();
 sg13g2_decap_8 FILLER_45_494 ();
 sg13g2_decap_8 FILLER_45_501 ();
 sg13g2_decap_8 FILLER_45_508 ();
 sg13g2_fill_1 FILLER_45_515 ();
 sg13g2_decap_8 FILLER_45_519 ();
 sg13g2_decap_8 FILLER_45_526 ();
 sg13g2_decap_8 FILLER_45_533 ();
 sg13g2_decap_8 FILLER_45_540 ();
 sg13g2_decap_8 FILLER_45_547 ();
 sg13g2_decap_8 FILLER_45_554 ();
 sg13g2_decap_8 FILLER_45_561 ();
 sg13g2_decap_8 FILLER_45_568 ();
 sg13g2_decap_8 FILLER_45_575 ();
 sg13g2_decap_8 FILLER_45_582 ();
 sg13g2_decap_8 FILLER_45_589 ();
 sg13g2_decap_8 FILLER_45_596 ();
 sg13g2_decap_8 FILLER_45_603 ();
 sg13g2_decap_8 FILLER_45_610 ();
 sg13g2_decap_8 FILLER_45_617 ();
 sg13g2_decap_8 FILLER_45_624 ();
 sg13g2_decap_8 FILLER_45_631 ();
 sg13g2_decap_8 FILLER_45_638 ();
 sg13g2_decap_8 FILLER_45_645 ();
 sg13g2_decap_8 FILLER_45_652 ();
 sg13g2_decap_8 FILLER_45_659 ();
 sg13g2_decap_8 FILLER_45_666 ();
 sg13g2_decap_8 FILLER_45_673 ();
 sg13g2_decap_8 FILLER_45_680 ();
 sg13g2_decap_8 FILLER_45_687 ();
 sg13g2_decap_8 FILLER_45_694 ();
 sg13g2_decap_8 FILLER_45_701 ();
 sg13g2_decap_8 FILLER_45_708 ();
 sg13g2_decap_8 FILLER_45_715 ();
 sg13g2_decap_8 FILLER_45_722 ();
 sg13g2_decap_8 FILLER_45_729 ();
 sg13g2_decap_8 FILLER_45_736 ();
 sg13g2_decap_8 FILLER_45_743 ();
 sg13g2_decap_8 FILLER_45_750 ();
 sg13g2_decap_8 FILLER_45_757 ();
 sg13g2_decap_8 FILLER_45_764 ();
 sg13g2_decap_8 FILLER_45_771 ();
 sg13g2_decap_8 FILLER_45_778 ();
 sg13g2_decap_8 FILLER_45_785 ();
 sg13g2_decap_8 FILLER_45_792 ();
 sg13g2_decap_8 FILLER_45_799 ();
 sg13g2_decap_8 FILLER_45_806 ();
 sg13g2_decap_8 FILLER_45_813 ();
 sg13g2_decap_8 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_827 ();
 sg13g2_decap_8 FILLER_45_834 ();
 sg13g2_decap_8 FILLER_45_841 ();
 sg13g2_fill_2 FILLER_45_848 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_136 ();
 sg13g2_decap_8 FILLER_46_143 ();
 sg13g2_decap_8 FILLER_46_150 ();
 sg13g2_decap_8 FILLER_46_157 ();
 sg13g2_decap_8 FILLER_46_164 ();
 sg13g2_decap_8 FILLER_46_171 ();
 sg13g2_decap_8 FILLER_46_178 ();
 sg13g2_decap_8 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_192 ();
 sg13g2_decap_8 FILLER_46_199 ();
 sg13g2_decap_8 FILLER_46_206 ();
 sg13g2_decap_8 FILLER_46_213 ();
 sg13g2_decap_8 FILLER_46_220 ();
 sg13g2_decap_8 FILLER_46_227 ();
 sg13g2_decap_8 FILLER_46_234 ();
 sg13g2_decap_8 FILLER_46_241 ();
 sg13g2_decap_8 FILLER_46_248 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_decap_8 FILLER_46_262 ();
 sg13g2_decap_8 FILLER_46_269 ();
 sg13g2_decap_8 FILLER_46_276 ();
 sg13g2_decap_8 FILLER_46_283 ();
 sg13g2_decap_8 FILLER_46_290 ();
 sg13g2_decap_8 FILLER_46_297 ();
 sg13g2_decap_8 FILLER_46_304 ();
 sg13g2_decap_8 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_318 ();
 sg13g2_decap_8 FILLER_46_325 ();
 sg13g2_decap_8 FILLER_46_332 ();
 sg13g2_decap_8 FILLER_46_339 ();
 sg13g2_decap_8 FILLER_46_346 ();
 sg13g2_decap_8 FILLER_46_353 ();
 sg13g2_decap_8 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_46_409 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_46_430 ();
 sg13g2_decap_8 FILLER_46_437 ();
 sg13g2_decap_8 FILLER_46_444 ();
 sg13g2_decap_8 FILLER_46_451 ();
 sg13g2_decap_8 FILLER_46_458 ();
 sg13g2_decap_8 FILLER_46_465 ();
 sg13g2_decap_8 FILLER_46_472 ();
 sg13g2_decap_8 FILLER_46_479 ();
 sg13g2_decap_8 FILLER_46_486 ();
 sg13g2_decap_8 FILLER_46_493 ();
 sg13g2_decap_8 FILLER_46_500 ();
 sg13g2_decap_8 FILLER_46_507 ();
 sg13g2_decap_8 FILLER_46_514 ();
 sg13g2_decap_8 FILLER_46_521 ();
 sg13g2_decap_8 FILLER_46_528 ();
 sg13g2_decap_8 FILLER_46_535 ();
 sg13g2_decap_8 FILLER_46_542 ();
 sg13g2_decap_8 FILLER_46_549 ();
 sg13g2_decap_8 FILLER_46_556 ();
 sg13g2_decap_8 FILLER_46_563 ();
 sg13g2_decap_8 FILLER_46_570 ();
 sg13g2_decap_8 FILLER_46_577 ();
 sg13g2_decap_8 FILLER_46_584 ();
 sg13g2_decap_8 FILLER_46_591 ();
 sg13g2_decap_8 FILLER_46_598 ();
 sg13g2_decap_8 FILLER_46_605 ();
 sg13g2_decap_8 FILLER_46_612 ();
 sg13g2_decap_8 FILLER_46_619 ();
 sg13g2_decap_8 FILLER_46_626 ();
 sg13g2_decap_8 FILLER_46_633 ();
 sg13g2_decap_8 FILLER_46_640 ();
 sg13g2_decap_8 FILLER_46_647 ();
 sg13g2_decap_8 FILLER_46_654 ();
 sg13g2_decap_8 FILLER_46_661 ();
 sg13g2_decap_8 FILLER_46_668 ();
 sg13g2_decap_8 FILLER_46_675 ();
 sg13g2_decap_8 FILLER_46_682 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_decap_8 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_703 ();
 sg13g2_decap_8 FILLER_46_710 ();
 sg13g2_decap_8 FILLER_46_717 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_745 ();
 sg13g2_decap_8 FILLER_46_752 ();
 sg13g2_decap_8 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_766 ();
 sg13g2_decap_8 FILLER_46_773 ();
 sg13g2_decap_8 FILLER_46_780 ();
 sg13g2_decap_8 FILLER_46_787 ();
 sg13g2_decap_8 FILLER_46_794 ();
 sg13g2_decap_8 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_4 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_298 ();
 sg13g2_decap_8 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_312 ();
 sg13g2_decap_8 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_decap_8 FILLER_49_340 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_8 FILLER_49_424 ();
 sg13g2_decap_8 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_494 ();
 sg13g2_decap_8 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_508 ();
 sg13g2_decap_8 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_522 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_550 ();
 sg13g2_decap_8 FILLER_49_557 ();
 sg13g2_decap_8 FILLER_49_564 ();
 sg13g2_decap_8 FILLER_49_571 ();
 sg13g2_decap_8 FILLER_49_578 ();
 sg13g2_decap_8 FILLER_49_585 ();
 sg13g2_decap_8 FILLER_49_592 ();
 sg13g2_decap_8 FILLER_49_599 ();
 sg13g2_decap_8 FILLER_49_606 ();
 sg13g2_decap_8 FILLER_49_613 ();
 sg13g2_decap_8 FILLER_49_620 ();
 sg13g2_decap_8 FILLER_49_627 ();
 sg13g2_decap_8 FILLER_49_634 ();
 sg13g2_decap_8 FILLER_49_641 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_decap_8 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_662 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_decap_8 FILLER_49_683 ();
 sg13g2_decap_8 FILLER_49_690 ();
 sg13g2_decap_8 FILLER_49_697 ();
 sg13g2_decap_8 FILLER_49_704 ();
 sg13g2_decap_8 FILLER_49_711 ();
 sg13g2_decap_8 FILLER_49_718 ();
 sg13g2_decap_8 FILLER_49_725 ();
 sg13g2_decap_8 FILLER_49_732 ();
 sg13g2_decap_8 FILLER_49_739 ();
 sg13g2_decap_8 FILLER_49_746 ();
 sg13g2_decap_8 FILLER_49_753 ();
 sg13g2_decap_8 FILLER_49_760 ();
 sg13g2_decap_8 FILLER_49_767 ();
 sg13g2_decap_8 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_781 ();
 sg13g2_decap_8 FILLER_49_788 ();
 sg13g2_decap_8 FILLER_49_795 ();
 sg13g2_decap_8 FILLER_49_802 ();
 sg13g2_decap_8 FILLER_49_809 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_decap_8 FILLER_49_823 ();
 sg13g2_decap_8 FILLER_49_830 ();
 sg13g2_decap_8 FILLER_49_837 ();
 sg13g2_decap_8 FILLER_49_844 ();
 sg13g2_decap_8 FILLER_49_851 ();
 sg13g2_decap_4 FILLER_49_858 ();
 assign uio_oe[0] = net;
 assign uio_oe[1] = net43;
 assign uio_oe[2] = net44;
 assign uio_oe[3] = net45;
 assign uio_oe[4] = net46;
 assign uio_oe[5] = net47;
 assign uio_oe[6] = net48;
 assign uio_oe[7] = net49;
 assign uo_out[0] = net50;
 assign uo_out[1] = net51;
 assign uo_out[2] = net52;
 assign uo_out[3] = net53;
 assign uo_out[4] = net54;
 assign uo_out[5] = net55;
 assign uo_out[6] = net56;
 assign uo_out[7] = net57;
endmodule
