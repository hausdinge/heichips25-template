module heichips25_internal (analog_adc,
    analog_pin0,
    analog_pin1,
    clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 inout analog_adc;
 inout analog_pin0;
 inout analog_pin1;
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire \adc_data[0] ;
 wire \adc_data[1] ;
 wire \adc_data[2] ;
 wire \adc_data[3] ;
 wire \adc_data[4] ;
 wire \adc_data[5] ;
 wire \adc_data[6] ;
 wire \adc_data[7] ;
 wire adc_ready;
 wire clk0_out;
 wire clk1_out;
 wire clk2_out;
 wire clk_delayed;
 wire \data[0] ;
 wire \data[10] ;
 wire \data[11] ;
 wire \data[12] ;
 wire \data[13] ;
 wire \data[14] ;
 wire \data[15] ;
 wire \data[16] ;
 wire \data[17] ;
 wire \data[18] ;
 wire \data[19] ;
 wire \data[1] ;
 wire \data[20] ;
 wire \data[21] ;
 wire \data[22] ;
 wire \data[23] ;
 wire \data[24] ;
 wire \data[25] ;
 wire \data[26] ;
 wire \data[27] ;
 wire \data[28] ;
 wire \data[29] ;
 wire \data[2] ;
 wire \data[30] ;
 wire \data[31] ;
 wire \data[32] ;
 wire \data[33] ;
 wire \data[34] ;
 wire \data[35] ;
 wire \data[36] ;
 wire \data[37] ;
 wire \data[38] ;
 wire \data[39] ;
 wire \data[3] ;
 wire \data[40] ;
 wire \data[41] ;
 wire \data[42] ;
 wire \data[43] ;
 wire \data[44] ;
 wire \data[45] ;
 wire \data[46] ;
 wire \data[47] ;
 wire \data[48] ;
 wire \data[49] ;
 wire \data[4] ;
 wire \data[50] ;
 wire \data[51] ;
 wire \data[52] ;
 wire \data[53] ;
 wire \data[54] ;
 wire \data[55] ;
 wire \data[56] ;
 wire \data[57] ;
 wire \data[58] ;
 wire \data[59] ;
 wire \data[5] ;
 wire \data[60] ;
 wire \data[61] ;
 wire \data[62] ;
 wire \data[63] ;
 wire \data[64] ;
 wire \data[65] ;
 wire \data[66] ;
 wire \data[67] ;
 wire \data[68] ;
 wire \data[69] ;
 wire \data[6] ;
 wire \data[70] ;
 wire \data[71] ;
 wire \data[72] ;
 wire \data[73] ;
 wire \data[74] ;
 wire \data[75] ;
 wire \data[76] ;
 wire \data[77] ;
 wire \data[78] ;
 wire \data[79] ;
 wire \data[7] ;
 wire \data[80] ;
 wire \data[81] ;
 wire \data[82] ;
 wire \data[83] ;
 wire \data[84] ;
 wire \data[85] ;
 wire \data[8] ;
 wire \data[9] ;
 wire osc_out;
 wire net1;
 wire stable;
 wire \u_custom_cells.u_latch0.D ;
 wire \u_custom_cells.u_latch0.Q ;
 wire \u_shift_reg.bit_count[0] ;
 wire \u_shift_reg.bit_count[1] ;
 wire \u_shift_reg.bit_count[2] ;
 wire \u_shift_reg.bit_count[3] ;
 wire \u_shift_reg.bit_count[4] ;
 wire \u_shift_reg.bit_count[5] ;
 wire \u_shift_reg.bit_count[6] ;
 wire \u_shift_reg.locked ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire clk_regs;
 wire VDD;
 wire VSS;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;

 sg13g2_inv_1 _128_ (.VDD(VPWR),
    .Y(_095_),
    .A(\u_shift_reg.bit_count[2] ),
    .VSS(VGND));
 sg13g2_inv_1 _129_ (.VDD(VPWR),
    .Y(_096_),
    .A(\data[83] ),
    .VSS(VGND));
 sg13g2_mux2_1 _130_ (.A0(\data[80] ),
    .A1(\data[81] ),
    .S(\data[82] ),
    .X(_097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _131_ (.A0(\data[78] ),
    .A1(\data[79] ),
    .S(\data[82] ),
    .X(_098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _132_ (.A(\data[83] ),
    .B(_098_),
    .Y(_099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _133_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\data[83] ),
    .A2(_097_),
    .Y(_000_),
    .B1(_099_));
 sg13g2_nor2b_1 _134_ (.A(net5),
    .B_N(net4),
    .Y(_100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _135_ (.A(\adc_data[0] ),
    .B(_100_),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _136_ (.A(\adc_data[1] ),
    .B(_100_),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _137_ (.A(\adc_data[2] ),
    .B(_100_),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _138_ (.A(_096_),
    .B(_098_),
    .Y(_101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _139_ (.A(net5),
    .B(net4),
    .X(_102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _140_ (.B1(_102_),
    .VDD(VPWR),
    .Y(_103_),
    .VSS(VGND),
    .A1(\data[83] ),
    .A2(\u_custom_cells.u_latch0.Q ));
 sg13g2_nor2_1 _141_ (.A(net5),
    .B(net4),
    .Y(_104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _142_ (.Y(_105_),
    .B1(_104_),
    .B2(stable),
    .A2(_100_),
    .A1(\adc_data[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _143_ (.B1(_105_),
    .VDD(VPWR),
    .Y(net9),
    .VSS(VGND),
    .A1(_101_),
    .A2(_103_));
 sg13g2_nand2_1 _144_ (.Y(_106_),
    .A(\adc_data[4] ),
    .B(_100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _145_ (.Y(_107_),
    .B1(_104_),
    .B2(osc_out),
    .A2(_102_),
    .A1(\u_custom_cells.u_latch0.D ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _146_ (.Y(net10),
    .A(_106_),
    .B(_107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _147_ (.Y(_108_),
    .A(\adc_data[5] ),
    .B(_100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _148_ (.Y(_109_),
    .B1(_104_),
    .B2(clk2_out),
    .A2(_102_),
    .A1(\u_custom_cells.u_latch0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _149_ (.Y(net11),
    .A(_108_),
    .B(_109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _150_ (.Y(_110_),
    .B(_102_),
    .A_N(_097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _151_ (.Y(_111_),
    .B1(_104_),
    .B2(clk1_out),
    .A2(_100_),
    .A1(\adc_data[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _152_ (.Y(net12),
    .A(_110_),
    .B(_111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _153_ (.S0(net4),
    .A0(clk0_out),
    .A1(\adc_data[7] ),
    .A2(clk_delayed),
    .A3(_098_),
    .S1(net5),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _154_ (.A(\u_shift_reg.locked ),
    .B_N(net2),
    .Y(_112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _155_ (.Y(_113_),
    .B(net2),
    .A_N(\u_shift_reg.locked ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _156_ (.A(\u_shift_reg.bit_count[0] ),
    .B(\u_shift_reg.bit_count[2] ),
    .X(_114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _157_ (.A(\u_shift_reg.bit_count[1] ),
    .B(\u_shift_reg.bit_count[3] ),
    .C(\u_shift_reg.bit_count[5] ),
    .Y(_115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _158_ (.B(\u_shift_reg.bit_count[6] ),
    .C(_114_),
    .A(\u_shift_reg.bit_count[4] ),
    .Y(_116_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_115_));
 sg13g2_inv_1 _159_ (.VDD(VPWR),
    .Y(_117_),
    .A(_116_),
    .VSS(VGND));
 sg13g2_nand3_1 _160_ (.B(net29),
    .C(_116_),
    .A(\u_shift_reg.bit_count[0] ),
    .Y(_118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _161_ (.A2(_116_),
    .A1(net29),
    .B1(\u_shift_reg.bit_count[0] ),
    .X(_119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _162_ (.A(_118_),
    .B(_119_),
    .X(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _163_ (.B(\u_shift_reg.bit_count[1] ),
    .C(net29),
    .A(\u_shift_reg.bit_count[0] ),
    .Y(_120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _164_ (.Y(_002_),
    .A(\u_shift_reg.bit_count[1] ),
    .B(_118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _165_ (.X(_121_),
    .A(\u_shift_reg.bit_count[1] ),
    .B(net29),
    .C(_114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _166_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_095_),
    .A2(_120_),
    .Y(_003_),
    .B1(_121_));
 sg13g2_xor2_1 _167_ (.B(_121_),
    .A(\u_shift_reg.bit_count[3] ),
    .X(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _168_ (.A(\u_shift_reg.bit_count[3] ),
    .B(\u_shift_reg.bit_count[4] ),
    .X(_122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _169_ (.A(\u_shift_reg.bit_count[1] ),
    .B(net29),
    .C(_114_),
    .D(_122_),
    .X(_123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _170_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_shift_reg.bit_count[3] ),
    .A2(_121_),
    .Y(_124_),
    .B1(\u_shift_reg.bit_count[4] ));
 sg13g2_nor2_1 _171_ (.A(_123_),
    .B(_124_),
    .Y(_005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _172_ (.Y(_125_),
    .A(\u_shift_reg.bit_count[5] ),
    .B(_123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _173_ (.B(_123_),
    .A(\u_shift_reg.bit_count[5] ),
    .X(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _174_ (.Y(_007_),
    .A(\u_shift_reg.bit_count[6] ),
    .B(_125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _175_ (.A0(\data[0] ),
    .A1(net3),
    .S(net29),
    .X(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _176_ (.A0(\data[0] ),
    .A1(\data[1] ),
    .S(net22),
    .X(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _177_ (.A0(\data[1] ),
    .A1(\data[2] ),
    .S(net22),
    .X(_010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _178_ (.A0(\data[2] ),
    .A1(\data[3] ),
    .S(net21),
    .X(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _179_ (.A0(\data[3] ),
    .A1(\data[4] ),
    .S(net21),
    .X(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _180_ (.A0(\data[4] ),
    .A1(\data[5] ),
    .S(net25),
    .X(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _181_ (.A0(\data[5] ),
    .A1(\data[6] ),
    .S(net25),
    .X(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _182_ (.A0(\data[6] ),
    .A1(\data[7] ),
    .S(net25),
    .X(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _183_ (.A0(\data[7] ),
    .A1(\data[8] ),
    .S(net25),
    .X(_016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _184_ (.A0(\data[8] ),
    .A1(\data[9] ),
    .S(net25),
    .X(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _185_ (.A0(\data[9] ),
    .A1(\data[10] ),
    .S(net21),
    .X(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _186_ (.A0(\data[10] ),
    .A1(\data[11] ),
    .S(net21),
    .X(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _187_ (.A0(\data[11] ),
    .A1(\data[12] ),
    .S(net21),
    .X(_020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _188_ (.A0(\data[12] ),
    .A1(\data[13] ),
    .S(net19),
    .X(_021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _189_ (.A0(\data[13] ),
    .A1(\data[14] ),
    .S(net19),
    .X(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _190_ (.A0(\data[14] ),
    .A1(\data[15] ),
    .S(net24),
    .X(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _191_ (.A0(\data[15] ),
    .A1(\data[16] ),
    .S(net24),
    .X(_024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _192_ (.A0(\data[16] ),
    .A1(\data[17] ),
    .S(net24),
    .X(_025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _193_ (.A0(\data[17] ),
    .A1(\data[18] ),
    .S(net25),
    .X(_026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _194_ (.A0(\data[18] ),
    .A1(\data[19] ),
    .S(net25),
    .X(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _195_ (.A0(\data[19] ),
    .A1(\data[20] ),
    .S(net24),
    .X(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _196_ (.A0(\data[20] ),
    .A1(\data[21] ),
    .S(net24),
    .X(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _197_ (.A0(\data[21] ),
    .A1(\data[22] ),
    .S(net24),
    .X(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _198_ (.A0(\data[22] ),
    .A1(\data[23] ),
    .S(net24),
    .X(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _199_ (.A0(\data[23] ),
    .A1(\data[24] ),
    .S(net20),
    .X(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _200_ (.A0(\data[24] ),
    .A1(\data[25] ),
    .S(net20),
    .X(_033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _201_ (.A0(\data[25] ),
    .A1(\data[26] ),
    .S(net19),
    .X(_034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _202_ (.A0(\data[26] ),
    .A1(\data[27] ),
    .S(net20),
    .X(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _203_ (.A0(\data[27] ),
    .A1(\data[28] ),
    .S(net20),
    .X(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _204_ (.A0(\data[28] ),
    .A1(\data[29] ),
    .S(net19),
    .X(_037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _205_ (.A0(\data[29] ),
    .A1(\data[30] ),
    .S(net19),
    .X(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _206_ (.A0(\data[30] ),
    .A1(\data[31] ),
    .S(net16),
    .X(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _207_ (.A0(\data[31] ),
    .A1(\data[32] ),
    .S(net16),
    .X(_040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _208_ (.A0(\data[32] ),
    .A1(\data[33] ),
    .S(net19),
    .X(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _209_ (.A0(\data[33] ),
    .A1(\data[34] ),
    .S(net19),
    .X(_042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _210_ (.A0(\data[34] ),
    .A1(\data[35] ),
    .S(net19),
    .X(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _211_ (.A0(\data[35] ),
    .A1(\data[36] ),
    .S(net20),
    .X(_044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _212_ (.A0(\data[36] ),
    .A1(\data[37] ),
    .S(net20),
    .X(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _213_ (.A0(\data[37] ),
    .A1(\data[38] ),
    .S(net20),
    .X(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _214_ (.A0(\data[38] ),
    .A1(\data[39] ),
    .S(net14),
    .X(_047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _215_ (.A0(\data[39] ),
    .A1(\data[40] ),
    .S(net17),
    .X(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _216_ (.A0(\data[40] ),
    .A1(\data[41] ),
    .S(net17),
    .X(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _217_ (.A0(\data[41] ),
    .A1(\data[42] ),
    .S(net17),
    .X(_050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _218_ (.A0(\data[42] ),
    .A1(\data[43] ),
    .S(net17),
    .X(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _219_ (.A0(\data[43] ),
    .A1(\data[44] ),
    .S(net17),
    .X(_052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _220_ (.A0(\data[44] ),
    .A1(\data[45] ),
    .S(net18),
    .X(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _221_ (.A0(\data[45] ),
    .A1(\data[46] ),
    .S(net17),
    .X(_054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _222_ (.A0(\data[46] ),
    .A1(\data[47] ),
    .S(net16),
    .X(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _223_ (.A0(\data[47] ),
    .A1(\data[48] ),
    .S(net14),
    .X(_056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _224_ (.A0(\data[48] ),
    .A1(\data[49] ),
    .S(net14),
    .X(_057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _225_ (.A0(\data[49] ),
    .A1(\data[50] ),
    .S(net14),
    .X(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _226_ (.A0(\data[50] ),
    .A1(\data[51] ),
    .S(net14),
    .X(_059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _227_ (.A0(\data[51] ),
    .A1(\data[52] ),
    .S(net15),
    .X(_060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _228_ (.A0(\data[52] ),
    .A1(\data[53] ),
    .S(net15),
    .X(_061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _229_ (.A0(\data[53] ),
    .A1(\data[54] ),
    .S(net17),
    .X(_062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _230_ (.A0(\data[54] ),
    .A1(\data[55] ),
    .S(net17),
    .X(_063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _231_ (.A0(\data[55] ),
    .A1(\data[56] ),
    .S(net18),
    .X(_064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _232_ (.A0(\data[56] ),
    .A1(\data[57] ),
    .S(net18),
    .X(_065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _233_ (.A0(\data[57] ),
    .A1(\data[58] ),
    .S(net18),
    .X(_066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _234_ (.A0(\data[58] ),
    .A1(\data[59] ),
    .S(net16),
    .X(_067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _235_ (.A0(\data[59] ),
    .A1(\data[60] ),
    .S(net16),
    .X(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _236_ (.A0(\data[60] ),
    .A1(\data[61] ),
    .S(net16),
    .X(_069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _237_ (.A0(\data[61] ),
    .A1(\data[62] ),
    .S(net14),
    .X(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _238_ (.A0(\data[62] ),
    .A1(\data[63] ),
    .S(net14),
    .X(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _239_ (.A0(\data[63] ),
    .A1(\data[64] ),
    .S(net14),
    .X(_072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _240_ (.A0(\data[64] ),
    .A1(\data[65] ),
    .S(net15),
    .X(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _241_ (.A0(\data[65] ),
    .A1(\data[66] ),
    .S(net28),
    .X(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _242_ (.A0(\data[66] ),
    .A1(\data[67] ),
    .S(net26),
    .X(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _243_ (.A0(\data[67] ),
    .A1(\data[68] ),
    .S(net26),
    .X(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _244_ (.A0(\data[68] ),
    .A1(\data[69] ),
    .S(net26),
    .X(_077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _245_ (.A0(\data[69] ),
    .A1(\data[70] ),
    .S(net26),
    .X(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _246_ (.A0(\data[70] ),
    .A1(\data[71] ),
    .S(net26),
    .X(_079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _247_ (.A0(\data[71] ),
    .A1(\data[72] ),
    .S(net26),
    .X(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _248_ (.A0(\data[72] ),
    .A1(\data[73] ),
    .S(net26),
    .X(_081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _249_ (.A0(\data[73] ),
    .A1(\data[74] ),
    .S(net26),
    .X(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _250_ (.A0(\data[74] ),
    .A1(\data[75] ),
    .S(net27),
    .X(_083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _251_ (.A0(\data[75] ),
    .A1(\data[76] ),
    .S(net27),
    .X(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _252_ (.A0(\data[76] ),
    .A1(\data[77] ),
    .S(net27),
    .X(_085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _253_ (.A0(\data[78] ),
    .A1(\data[77] ),
    .S(net29),
    .X(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _254_ (.A0(\data[78] ),
    .A1(\data[79] ),
    .S(net28),
    .X(_087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _255_ (.A0(\data[79] ),
    .A1(\data[80] ),
    .S(net21),
    .X(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _256_ (.A0(\data[80] ),
    .A1(\data[81] ),
    .S(net21),
    .X(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _257_ (.A0(\data[82] ),
    .A1(\data[81] ),
    .S(net29),
    .X(_090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _258_ (.A(\data[82] ),
    .B(net21),
    .Y(_126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _259_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_096_),
    .A2(net22),
    .Y(_091_),
    .B1(_126_));
 sg13g2_nor2_1 _260_ (.A(\data[84] ),
    .B(_112_),
    .Y(_127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_096_),
    .A2(_112_),
    .Y(_092_),
    .B1(_127_));
 sg13g2_mux2_1 _262_ (.A0(\data[84] ),
    .A1(\data[85] ),
    .S(net24),
    .X(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _263_ (.A2(_117_),
    .A1(net2),
    .B1(\u_shift_reg.locked ),
    .X(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _264_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_001_),
    .Q(\u_shift_reg.bit_count[0] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _265_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_002_),
    .Q(\u_shift_reg.bit_count[1] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _266_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_003_),
    .Q(\u_shift_reg.bit_count[2] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _267_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_004_),
    .Q(\u_shift_reg.bit_count[3] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _268_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_005_),
    .Q(\u_shift_reg.bit_count[4] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _269_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_006_),
    .Q(\u_shift_reg.bit_count[5] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _270_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_007_),
    .Q(\u_shift_reg.bit_count[6] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _271_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_008_),
    .Q(\data[0] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _272_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_009_),
    .Q(\data[1] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _273_ (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_010_),
    .Q(\data[2] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _274_ (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_011_),
    .Q(\data[3] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _275_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_012_),
    .Q(\data[4] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _276_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_013_),
    .Q(\data[5] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _277_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_014_),
    .Q(\data[6] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _278_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_015_),
    .Q(\data[7] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _279_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_016_),
    .Q(\data[8] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _280_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_017_),
    .Q(\data[9] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _281_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_018_),
    .Q(\data[10] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _282_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_019_),
    .Q(\data[11] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _283_ (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_020_),
    .Q(\data[12] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _284_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_021_),
    .Q(\data[13] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _285_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_022_),
    .Q(\data[14] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _286_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_023_),
    .Q(\data[15] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _287_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_024_),
    .Q(\data[16] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _288_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_025_),
    .Q(\data[17] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _289_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_026_),
    .Q(\data[18] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _290_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_027_),
    .Q(\data[19] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _291_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_028_),
    .Q(\data[20] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _292_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_029_),
    .Q(\data[21] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _293_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_030_),
    .Q(\data[22] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _294_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_031_),
    .Q(\data[23] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _295_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_032_),
    .Q(\data[24] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _296_ (.RESET_B(net36),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_033_),
    .Q(\data[25] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _297_ (.RESET_B(net36),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_034_),
    .Q(\data[26] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _298_ (.RESET_B(net36),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_035_),
    .Q(\data[27] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _299_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_036_),
    .Q(\data[28] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _300_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_037_),
    .Q(\data[29] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _301_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_038_),
    .Q(\data[30] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _302_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_039_),
    .Q(\data[31] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _303_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_040_),
    .Q(\data[32] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _304_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_041_),
    .Q(\data[33] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _305_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_042_),
    .Q(\data[34] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _306_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_043_),
    .Q(\data[35] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _307_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_044_),
    .Q(\data[36] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _308_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_045_),
    .Q(\data[37] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _309_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_046_),
    .Q(\data[38] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _310_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_047_),
    .Q(\data[39] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _311_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_048_),
    .Q(\data[40] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _312_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_049_),
    .Q(\data[41] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _313_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_050_),
    .Q(\data[42] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _314_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_051_),
    .Q(\data[43] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _315_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_052_),
    .Q(\data[44] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _316_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_053_),
    .Q(\data[45] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _317_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_054_),
    .Q(\data[46] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _318_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_055_),
    .Q(\data[47] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _319_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_056_),
    .Q(\data[48] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _320_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_057_),
    .Q(\data[49] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _321_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_058_),
    .Q(\data[50] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _322_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_059_),
    .Q(\data[51] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _323_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_060_),
    .Q(\data[52] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _324_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_061_),
    .Q(\data[53] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _325_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_062_),
    .Q(\data[54] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _326_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_063_),
    .Q(\data[55] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _327_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_064_),
    .Q(\data[56] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _328_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_065_),
    .Q(\data[57] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _329_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_066_),
    .Q(\data[58] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _330_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_067_),
    .Q(\data[59] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _331_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_068_),
    .Q(\data[60] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _332_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_069_),
    .Q(\data[61] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _333_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_070_),
    .Q(\data[62] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _334_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_071_),
    .Q(\data[63] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _335_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_072_),
    .Q(\data[64] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _336_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_073_),
    .Q(\data[65] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _337_ (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_074_),
    .Q(\data[66] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _338_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_075_),
    .Q(\data[67] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _339_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_076_),
    .Q(\data[68] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _340_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_077_),
    .Q(\data[69] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _341_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_078_),
    .Q(\data[70] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _342_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_079_),
    .Q(\data[71] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _343_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_080_),
    .Q(\data[72] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _344_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_081_),
    .Q(\data[73] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _345_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_082_),
    .Q(\data[74] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _346_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_083_),
    .Q(\data[75] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _347_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_084_),
    .Q(\data[76] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _348_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_085_),
    .Q(\data[77] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _349_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_086_),
    .Q(\data[78] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _350_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_087_),
    .Q(\data[79] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _351_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_088_),
    .Q(\data[80] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _352_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_089_),
    .Q(\data[81] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _353_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_090_),
    .Q(\data[82] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _354_ (.RESET_B(net41),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_091_),
    .Q(\data[83] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _355_ (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_092_),
    .Q(\data[84] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _356_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_093_),
    .Q(\data[85] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _357_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_094_),
    .Q(\u_shift_reg.locked ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dlhq_1 _358_ (.D(_000_),
    .GATE(\data[84] ),
    .Q(\u_custom_cells.u_latch0.D ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _359_ (.D(\u_custom_cells.u_latch0.D ),
    .GATE(\data[85] ),
    .Q(\u_custom_cells.u_latch0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_internal_47 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net47));
 sg13g2_tielo heichips25_internal_48 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net48));
 sg13g2_tielo heichips25_internal_49 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net49));
 sg13g2_tielo heichips25_internal_50 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net50));
 sg13g2_tielo heichips25_internal_51 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net51));
 sg13g2_tielo heichips25_internal_52 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net52));
 sg13g2_tielo heichips25_internal_53 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net53));
 sg13g2_tielo heichips25_internal_54 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net54));
 sg13g2_tielo heichips25_internal_55 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net55));
 sg13g2_tielo heichips25_internal_56 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net56));
 sg13g2_tielo heichips25_internal_57 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net57));
 sg13g2_tielo heichips25_internal_58 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net58));
 sg13g2_tielo heichips25_internal_59 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net59));
 sg13g2_tielo heichips25_internal_60 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net60));
 sg13g2_tielo heichips25_internal_61 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net61));
 sg13g2_buf_16 clkbuf_regs_0_clk (.X(clk_regs),
    .A(clk),
    .VDD(VPWR),
    .VSS(VGND));
 adc u_adc (.VDD(VPWR),
    .VSS(VGND),
    .analog_in(analog_adc),
    .clk(clknet_1_1__leaf_clk),
    .ready(adc_ready),
    .start(\data[66] ),
    .data_out({\adc_data[7] ,
    \adc_data[6] ,
    \adc_data[5] ,
    \adc_data[4] ,
    \adc_data[3] ,
    \adc_data[2] ,
    \adc_data[1] ,
    \adc_data[0] }));
 sg13g2_buf_16 \u_clkbuf_analog_pin0.u_buf  (.X(analog_pin0),
    .A(clk0_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 \u_clkbuf_analog_pin1.u_buf  (.X(analog_pin1),
    .A(clk1_out),
    .VDD(VPWR),
    .VSS(VGND));
 delay_line u_delay_line (.VDD(VPWR),
    .VSS(VGND),
    .clk(clknet_1_0__leaf_clk),
    .clk_delayed(clk_delayed),
    .reset(net44),
    .sel({\data[77] ,
    \data[76] ,
    \data[75] }),
    .trim({\data[74] ,
    \data[73] ,
    \data[72] ,
    \data[71] ,
    \data[70] ,
    \data[69] ,
    \data[68] ,
    \data[67] }));
 multimode_dll u_multimode_dll (.VDD(VPWR),
    .VSS(VGND),
    .bias(\data[38] ),
    .clk0_out(clk0_out),
    .clk1_out(clk1_out),
    .clk2_out(clk2_out),
    .dco(\data[39] ),
    .enable(ena),
    .osc(clknet_1_0__leaf_clk),
    .osc_out(osc_out),
    .resetb(net35),
    .stable(stable),
    .clk0_phase_sel({\data[24] ,
    \data[23] ,
    \data[22] ,
    \data[21] ,
    \data[20] }),
    .clk1_phase_sel({\data[29] ,
    \data[28] ,
    \data[27] ,
    \data[26] ,
    \data[25] }),
    .clk2_phase_sel({\data[34] ,
    \data[33] ,
    \data[32] ,
    \data[31] ,
    \data[30] }),
    .ext_trim({\data[65] ,
    \data[64] ,
    \data[63] ,
    \data[62] ,
    \data[61] ,
    \data[60] ,
    \data[59] ,
    \data[58] ,
    \data[57] ,
    \data[56] ,
    \data[55] ,
    \data[54] ,
    \data[53] ,
    \data[52] ,
    \data[51] ,
    \data[50] ,
    \data[49] ,
    \data[48] ,
    \data[47] ,
    \data[46] ,
    \data[45] ,
    \data[44] ,
    \data[43] ,
    \data[42] ,
    \data[41] ,
    \data[40] }),
    .f_clk0_divider({\data[9] ,
    \data[8] ,
    \data[7] ,
    \data[6] ,
    \data[5] }),
    .f_clk1_divider({\data[14] ,
    \data[13] ,
    \data[12] ,
    \data[11] ,
    \data[10] }),
    .f_clk2_divider({\data[19] ,
    \data[18] ,
    \data[17] ,
    \data[16] ,
    \data[15] }),
    .f_osc_multiply_factor({\data[4] ,
    \data[3] ,
    \data[2] ,
    \data[1] ,
    \data[0] }),
    .mode_xor({\data[37] ,
    \data[36] ,
    \data[35] }));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout14 (.A(net15),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout15 (.A(net16),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout16 (.A(net23),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout17 (.A(net23),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout18 (.A(net23),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout19 (.A(net20),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout20 (.A(net23),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout21 (.A(net22),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout22 (.A(net23),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout23 (.A(_113_),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout24 (.A(net25),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout25 (.A(net28),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout26 (.A(net27),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout27 (.A(net28),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout28 (.A(_113_),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout29 (.A(_112_),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout30 (.A(net31),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout31 (.A(net32),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout32 (.A(net41),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout33 (.A(net41),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout34 (.A(net41),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout35 (.A(net36),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout36 (.A(net37),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout37 (.A(net41),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout38 (.A(net39),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout39 (.A(net40),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout40 (.A(net41),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout41 (.A(net1),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout42 (.A(net43),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout43 (.A(net46),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout44 (.A(net46),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout45 (.A(net46),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout46 (.A(net1),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_internal (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(delaynet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_1_0__f_clk (.X(clknet_1_0__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_1_1__f_clk (.X(clknet_1_1__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_0_clk_regs (.X(clknet_0_clk_regs),
    .A(clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload0 (.VDD(VPWR),
    .A(clknet_4_7_0_clk_regs),
    .VSS(VGND));
 sg13g2_inv_1 clkload1 (.VDD(VPWR),
    .A(clknet_4_15_0_clk_regs),
    .VSS(VGND));
 sg13g2_buf_16 delaybuf_0_clk (.X(delaynet_0_clk),
    .A(clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(\adc_data[6] ));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(_101_));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(\adc_data[0] ));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(\adc_data[0] ));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(\adc_data[2] ));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_860 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net;
 assign uio_oe[1] = net47;
 assign uio_oe[2] = net48;
 assign uio_oe[3] = net49;
 assign uio_oe[4] = net50;
 assign uio_oe[5] = net51;
 assign uio_oe[6] = net52;
 assign uio_oe[7] = net53;
 assign uo_out[0] = net54;
 assign uo_out[1] = net55;
 assign uo_out[2] = net56;
 assign uo_out[3] = net57;
 assign uo_out[4] = net58;
 assign uo_out[5] = net59;
 assign uo_out[6] = net60;
 assign uo_out[7] = net61;
endmodule
