magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771728784
<< metal1 >>
rect 576 38576 83328 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 83328 38576
rect 576 38512 83328 38536
rect 20995 38408 21053 38409
rect 20995 38368 21004 38408
rect 21044 38368 21053 38408
rect 20995 38367 21053 38368
rect 27139 38408 27197 38409
rect 27139 38368 27148 38408
rect 27188 38368 27197 38408
rect 27139 38367 27197 38368
rect 27043 38324 27101 38325
rect 27043 38284 27052 38324
rect 27092 38284 27101 38324
rect 27043 38283 27101 38284
rect 28963 38324 29021 38325
rect 28963 38284 28972 38324
rect 29012 38284 29021 38324
rect 28963 38283 29021 38284
rect 21091 38240 21149 38241
rect 21091 38200 21100 38240
rect 21140 38200 21149 38240
rect 21091 38199 21149 38200
rect 26859 38240 26901 38249
rect 26859 38200 26860 38240
rect 26900 38200 26901 38240
rect 26859 38191 26901 38200
rect 26955 38240 26997 38249
rect 26955 38200 26956 38240
rect 26996 38200 26997 38240
rect 26955 38191 26997 38200
rect 28483 38240 28541 38241
rect 28483 38200 28492 38240
rect 28532 38200 28541 38240
rect 28483 38199 28541 38200
rect 28867 38240 28925 38241
rect 28867 38200 28876 38240
rect 28916 38200 28925 38240
rect 28867 38199 28925 38200
rect 29259 38240 29301 38249
rect 29259 38200 29260 38240
rect 29300 38200 29301 38240
rect 29259 38191 29301 38200
rect 29443 38240 29501 38241
rect 29443 38200 29452 38240
rect 29492 38200 29501 38240
rect 29443 38199 29501 38200
rect 38467 38240 38525 38241
rect 38467 38200 38476 38240
rect 38516 38200 38525 38240
rect 38467 38199 38525 38200
rect 38763 38240 38805 38249
rect 38763 38200 38764 38240
rect 38804 38200 38805 38240
rect 38763 38191 38805 38200
rect 38859 38240 38901 38249
rect 38859 38200 38860 38240
rect 38900 38200 38901 38240
rect 38859 38191 38901 38200
rect 41059 38240 41117 38241
rect 41059 38200 41068 38240
rect 41108 38200 41117 38240
rect 41059 38199 41117 38200
rect 41355 38240 41397 38249
rect 41355 38200 41356 38240
rect 41396 38200 41397 38240
rect 41355 38191 41397 38200
rect 41451 38240 41493 38249
rect 41451 38200 41452 38240
rect 41492 38200 41493 38240
rect 41451 38191 41493 38200
rect 70347 38240 70389 38249
rect 70347 38200 70348 38240
rect 70388 38200 70389 38240
rect 70347 38191 70389 38200
rect 643 38156 701 38157
rect 643 38116 652 38156
rect 692 38116 701 38156
rect 643 38115 701 38116
rect 21763 38156 21821 38157
rect 21763 38116 21772 38156
rect 21812 38116 21821 38156
rect 21763 38115 21821 38116
rect 23203 38156 23261 38157
rect 23203 38116 23212 38156
rect 23252 38116 23261 38156
rect 23203 38115 23261 38116
rect 23587 38156 23645 38157
rect 23587 38116 23596 38156
rect 23636 38116 23645 38156
rect 23587 38115 23645 38116
rect 23971 38156 24029 38157
rect 23971 38116 23980 38156
rect 24020 38116 24029 38156
rect 23971 38115 24029 38116
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 21283 37988 21341 37989
rect 21283 37948 21292 37988
rect 21332 37948 21341 37988
rect 21283 37947 21341 37948
rect 21963 37988 22005 37997
rect 21963 37948 21964 37988
rect 22004 37948 22005 37988
rect 21963 37939 22005 37948
rect 23403 37988 23445 37997
rect 23403 37948 23404 37988
rect 23444 37948 23445 37988
rect 23403 37939 23445 37948
rect 23787 37988 23829 37997
rect 23787 37948 23788 37988
rect 23828 37948 23829 37988
rect 23787 37939 23829 37948
rect 24171 37988 24213 37997
rect 24171 37948 24172 37988
rect 24212 37948 24213 37988
rect 24171 37939 24213 37948
rect 26955 37988 26997 37997
rect 26955 37948 26956 37988
rect 26996 37948 26997 37988
rect 26955 37939 26997 37948
rect 29355 37988 29397 37997
rect 29355 37948 29356 37988
rect 29396 37948 29397 37988
rect 29355 37939 29397 37948
rect 39139 37988 39197 37989
rect 39139 37948 39148 37988
rect 39188 37948 39197 37988
rect 39139 37947 39197 37948
rect 41731 37988 41789 37989
rect 41731 37948 41740 37988
rect 41780 37948 41789 37988
rect 41731 37947 41789 37948
rect 70539 37988 70581 37997
rect 70539 37948 70540 37988
rect 70580 37948 70581 37988
rect 70539 37939 70581 37948
rect 576 37820 83328 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 83328 37820
rect 576 37756 83328 37780
rect 26091 37568 26133 37577
rect 26091 37528 26092 37568
rect 26132 37528 26133 37568
rect 26091 37519 26133 37528
rect 41923 37568 41981 37569
rect 41923 37528 41932 37568
rect 41972 37528 41981 37568
rect 41923 37527 41981 37528
rect 19275 37400 19317 37409
rect 19275 37360 19276 37400
rect 19316 37360 19317 37400
rect 19275 37351 19317 37360
rect 19371 37400 19413 37409
rect 19371 37360 19372 37400
rect 19412 37360 19413 37400
rect 19371 37351 19413 37360
rect 20515 37400 20573 37401
rect 20515 37360 20524 37400
rect 20564 37360 20573 37400
rect 20515 37359 20573 37360
rect 21379 37400 21437 37401
rect 21379 37360 21388 37400
rect 21428 37360 21437 37400
rect 21379 37359 21437 37360
rect 23107 37400 23165 37401
rect 23107 37360 23116 37400
rect 23156 37360 23165 37400
rect 23107 37359 23165 37360
rect 23971 37400 24029 37401
rect 23971 37360 23980 37400
rect 24020 37360 24029 37400
rect 23971 37359 24029 37360
rect 25899 37400 25941 37409
rect 25899 37360 25900 37400
rect 25940 37360 25941 37400
rect 25899 37351 25941 37360
rect 26091 37400 26133 37409
rect 26091 37360 26092 37400
rect 26132 37360 26133 37400
rect 26091 37351 26133 37360
rect 26283 37400 26325 37409
rect 26283 37360 26284 37400
rect 26324 37360 26325 37400
rect 26283 37351 26325 37360
rect 26659 37400 26717 37401
rect 26659 37360 26668 37400
rect 26708 37360 26717 37400
rect 26659 37359 26717 37360
rect 27523 37400 27581 37401
rect 27523 37360 27532 37400
rect 27572 37360 27581 37400
rect 27523 37359 27581 37360
rect 29355 37400 29397 37409
rect 29355 37360 29356 37400
rect 29396 37360 29397 37400
rect 29355 37351 29397 37360
rect 29443 37400 29501 37401
rect 29443 37360 29452 37400
rect 29492 37360 29501 37400
rect 29443 37359 29501 37360
rect 30307 37400 30365 37401
rect 30307 37360 30316 37400
rect 30356 37360 30365 37400
rect 30307 37359 30365 37360
rect 31171 37400 31229 37401
rect 31171 37360 31180 37400
rect 31220 37360 31229 37400
rect 31171 37359 31229 37360
rect 38179 37400 38237 37401
rect 38179 37360 38188 37400
rect 38228 37360 38237 37400
rect 38179 37359 38237 37360
rect 39043 37400 39101 37401
rect 39043 37360 39052 37400
rect 39092 37360 39101 37400
rect 39043 37359 39101 37360
rect 41251 37400 41309 37401
rect 41251 37360 41260 37400
rect 41300 37360 41309 37400
rect 41251 37359 41309 37360
rect 41547 37400 41589 37409
rect 41547 37360 41548 37400
rect 41588 37360 41589 37400
rect 41547 37351 41589 37360
rect 42123 37400 42165 37409
rect 42123 37360 42124 37400
rect 42164 37360 42165 37400
rect 42123 37351 42165 37360
rect 42499 37400 42557 37401
rect 42499 37360 42508 37400
rect 42548 37360 42557 37400
rect 42499 37359 42557 37360
rect 43363 37400 43421 37401
rect 43363 37360 43372 37400
rect 43412 37360 43421 37400
rect 43363 37359 43421 37360
rect 20139 37316 20181 37325
rect 20139 37276 20140 37316
rect 20180 37276 20181 37316
rect 20139 37267 20181 37276
rect 22731 37316 22773 37325
rect 22731 37276 22732 37316
rect 22772 37276 22773 37316
rect 22731 37267 22773 37276
rect 29931 37316 29973 37325
rect 29931 37276 29932 37316
rect 29972 37276 29973 37316
rect 29931 37267 29973 37276
rect 37803 37316 37845 37325
rect 37803 37276 37804 37316
rect 37844 37276 37845 37316
rect 37803 37267 37845 37276
rect 41643 37316 41685 37325
rect 41643 37276 41644 37316
rect 41684 37276 41685 37316
rect 41643 37267 41685 37276
rect 19555 37232 19613 37233
rect 19555 37192 19564 37232
rect 19604 37192 19613 37232
rect 19555 37191 19613 37192
rect 22531 37232 22589 37233
rect 22531 37192 22540 37232
rect 22580 37192 22589 37232
rect 22531 37191 22589 37192
rect 25123 37232 25181 37233
rect 25123 37192 25132 37232
rect 25172 37192 25181 37232
rect 25123 37191 25181 37192
rect 28675 37232 28733 37233
rect 28675 37192 28684 37232
rect 28724 37192 28733 37232
rect 28675 37191 28733 37192
rect 29739 37232 29781 37241
rect 29739 37192 29740 37232
rect 29780 37192 29781 37232
rect 29739 37183 29781 37192
rect 32323 37232 32381 37233
rect 32323 37192 32332 37232
rect 32372 37192 32381 37232
rect 32323 37191 32381 37192
rect 40195 37232 40253 37233
rect 40195 37192 40204 37232
rect 40244 37192 40253 37232
rect 40195 37191 40253 37192
rect 44515 37232 44573 37233
rect 44515 37192 44524 37232
rect 44564 37192 44573 37232
rect 44515 37191 44573 37192
rect 576 37064 83328 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 83328 37064
rect 576 37000 83328 37024
rect 21771 36954 21813 36963
rect 21771 36914 21772 36954
rect 21812 36914 21813 36954
rect 21771 36905 21813 36914
rect 20619 36896 20661 36905
rect 20619 36856 20620 36896
rect 20660 36856 20661 36896
rect 20619 36847 20661 36856
rect 22635 36896 22677 36905
rect 22635 36856 22636 36896
rect 22676 36856 22677 36896
rect 22635 36847 22677 36856
rect 24355 36896 24413 36897
rect 24355 36856 24364 36896
rect 24404 36856 24413 36896
rect 24355 36855 24413 36856
rect 25219 36896 25277 36897
rect 25219 36856 25228 36896
rect 25268 36856 25277 36896
rect 25219 36855 25277 36856
rect 25987 36896 26045 36897
rect 25987 36856 25996 36896
rect 26036 36856 26045 36896
rect 25987 36855 26045 36856
rect 26947 36896 27005 36897
rect 26947 36856 26956 36896
rect 26996 36856 27005 36896
rect 26947 36855 27005 36856
rect 27243 36896 27285 36905
rect 27243 36856 27244 36896
rect 27284 36856 27285 36896
rect 27243 36847 27285 36856
rect 27619 36896 27677 36897
rect 27619 36856 27628 36896
rect 27668 36856 27677 36896
rect 27619 36855 27677 36856
rect 31459 36896 31517 36897
rect 31459 36856 31468 36896
rect 31508 36856 31517 36896
rect 31459 36855 31517 36856
rect 43459 36896 43517 36897
rect 43459 36856 43468 36896
rect 43508 36856 43517 36896
rect 43459 36855 43517 36856
rect 24643 36812 24701 36813
rect 24643 36772 24652 36812
rect 24692 36772 24701 36812
rect 24643 36771 24701 36772
rect 27907 36812 27965 36813
rect 27907 36772 27916 36812
rect 27956 36772 27965 36812
rect 27907 36771 27965 36772
rect 29067 36812 29109 36821
rect 29067 36772 29068 36812
rect 29108 36772 29109 36812
rect 29067 36763 29109 36772
rect 41067 36812 41109 36821
rect 41067 36772 41068 36812
rect 41108 36772 41109 36812
rect 41067 36763 41109 36772
rect 17835 36728 17877 36737
rect 17835 36688 17836 36728
rect 17876 36688 17877 36728
rect 17835 36679 17877 36688
rect 18211 36728 18269 36729
rect 18211 36688 18220 36728
rect 18260 36688 18269 36728
rect 18211 36687 18269 36688
rect 19075 36728 19133 36729
rect 19075 36688 19084 36728
rect 19124 36688 19133 36728
rect 19075 36687 19133 36688
rect 20427 36728 20469 36737
rect 20427 36688 20428 36728
rect 20468 36688 20469 36728
rect 20427 36679 20469 36688
rect 20715 36728 20757 36737
rect 20715 36688 20716 36728
rect 20756 36688 20757 36728
rect 20715 36679 20757 36688
rect 20899 36728 20957 36729
rect 20899 36688 20908 36728
rect 20948 36688 20957 36728
rect 20899 36687 20957 36688
rect 21579 36728 21621 36737
rect 21579 36688 21580 36728
rect 21620 36688 21621 36728
rect 21579 36679 21621 36688
rect 21667 36728 21725 36729
rect 21667 36688 21676 36728
rect 21716 36688 21725 36728
rect 21667 36687 21725 36688
rect 22251 36728 22293 36737
rect 22251 36688 22252 36728
rect 22292 36688 22293 36728
rect 22251 36679 22293 36688
rect 22339 36728 22397 36729
rect 22339 36688 22348 36728
rect 22388 36688 22397 36728
rect 22339 36687 22397 36688
rect 22915 36728 22973 36729
rect 22915 36688 22924 36728
rect 22964 36688 22973 36728
rect 22915 36687 22973 36688
rect 23019 36728 23061 36737
rect 23019 36688 23020 36728
rect 23060 36688 23061 36728
rect 23019 36679 23061 36688
rect 23203 36728 23261 36729
rect 23203 36688 23212 36728
rect 23252 36688 23261 36728
rect 23203 36687 23261 36688
rect 23307 36728 23349 36737
rect 23307 36688 23308 36728
rect 23348 36688 23349 36728
rect 23307 36679 23349 36688
rect 23491 36728 23549 36729
rect 23491 36688 23500 36728
rect 23540 36688 23549 36728
rect 23491 36687 23549 36688
rect 23691 36728 23733 36737
rect 23691 36688 23692 36728
rect 23732 36688 23733 36728
rect 23691 36679 23733 36688
rect 23883 36728 23925 36737
rect 23883 36688 23884 36728
rect 23924 36688 23925 36728
rect 23883 36679 23925 36688
rect 23971 36728 24029 36729
rect 23971 36688 23980 36728
rect 24020 36688 24029 36728
rect 23971 36687 24029 36688
rect 24451 36728 24509 36729
rect 24451 36688 24460 36728
rect 24500 36688 24509 36728
rect 24451 36687 24509 36688
rect 25227 36728 25269 36737
rect 25227 36688 25228 36728
rect 25268 36688 25269 36728
rect 25227 36679 25269 36688
rect 25323 36728 25365 36737
rect 25323 36688 25324 36728
rect 25364 36688 25365 36728
rect 25323 36679 25365 36688
rect 25899 36728 25941 36737
rect 25899 36688 25900 36728
rect 25940 36688 25941 36728
rect 25899 36679 25941 36688
rect 26091 36728 26133 36737
rect 26091 36688 26092 36728
rect 26132 36688 26133 36728
rect 26091 36679 26133 36688
rect 26179 36728 26237 36729
rect 26179 36688 26188 36728
rect 26228 36688 26237 36728
rect 26179 36687 26237 36688
rect 26475 36728 26517 36737
rect 26475 36688 26476 36728
rect 26516 36688 26517 36728
rect 26475 36679 26517 36688
rect 26571 36728 26613 36737
rect 26571 36688 26572 36728
rect 26612 36688 26613 36728
rect 26571 36679 26613 36688
rect 26667 36728 26709 36737
rect 26667 36688 26668 36728
rect 26708 36688 26709 36728
rect 26667 36679 26709 36688
rect 26763 36728 26805 36737
rect 26763 36688 26764 36728
rect 26804 36688 26805 36728
rect 26763 36679 26805 36688
rect 27147 36728 27189 36737
rect 27147 36688 27148 36728
rect 27188 36688 27189 36728
rect 27147 36679 27189 36688
rect 27339 36728 27381 36737
rect 27339 36688 27340 36728
rect 27380 36688 27381 36728
rect 27339 36679 27381 36688
rect 27435 36728 27477 36737
rect 27435 36688 27436 36728
rect 27476 36688 27477 36728
rect 27435 36679 27477 36688
rect 27715 36728 27773 36729
rect 27715 36688 27724 36728
rect 27764 36688 27773 36728
rect 27715 36687 27773 36688
rect 29443 36728 29501 36729
rect 29443 36688 29452 36728
rect 29492 36688 29501 36728
rect 29443 36687 29501 36688
rect 30307 36728 30365 36729
rect 30307 36688 30316 36728
rect 30356 36688 30365 36728
rect 30307 36687 30365 36688
rect 32427 36728 32469 36737
rect 32427 36688 32428 36728
rect 32468 36688 32469 36728
rect 32427 36679 32469 36688
rect 32803 36728 32861 36729
rect 32803 36688 32812 36728
rect 32852 36688 32861 36728
rect 32803 36687 32861 36688
rect 33667 36728 33725 36729
rect 33667 36688 33676 36728
rect 33716 36688 33725 36728
rect 33667 36687 33725 36688
rect 35107 36728 35165 36729
rect 35107 36688 35116 36728
rect 35156 36688 35165 36728
rect 35107 36687 35165 36688
rect 35403 36728 35445 36737
rect 35403 36688 35404 36728
rect 35444 36688 35445 36728
rect 35403 36679 35445 36688
rect 35499 36728 35541 36737
rect 35499 36688 35500 36728
rect 35540 36688 35541 36728
rect 35499 36679 35541 36688
rect 38475 36728 38517 36737
rect 38475 36688 38476 36728
rect 38516 36688 38517 36728
rect 38475 36679 38517 36688
rect 38851 36728 38909 36729
rect 38851 36688 38860 36728
rect 38900 36688 38909 36728
rect 38851 36687 38909 36688
rect 39715 36728 39773 36729
rect 39715 36688 39724 36728
rect 39764 36688 39773 36728
rect 39715 36687 39773 36688
rect 41443 36728 41501 36729
rect 41443 36688 41452 36728
rect 41492 36688 41501 36728
rect 41443 36687 41501 36688
rect 42307 36728 42365 36729
rect 42307 36688 42316 36728
rect 42356 36688 42365 36728
rect 42307 36687 42365 36688
rect 20235 36644 20277 36653
rect 20235 36604 20236 36644
rect 20276 36604 20277 36644
rect 20235 36595 20277 36604
rect 44899 36644 44957 36645
rect 44899 36604 44908 36644
rect 44948 36604 44957 36644
rect 44899 36603 44957 36604
rect 45283 36644 45341 36645
rect 45283 36604 45292 36644
rect 45332 36604 45341 36644
rect 45283 36603 45341 36604
rect 21291 36560 21333 36569
rect 21291 36520 21292 36560
rect 21332 36520 21333 36560
rect 21291 36511 21333 36520
rect 23499 36560 23541 36569
rect 23499 36520 23500 36560
rect 23540 36520 23541 36560
rect 23499 36511 23541 36520
rect 21003 36476 21045 36485
rect 21003 36436 21004 36476
rect 21044 36436 21045 36476
rect 21003 36427 21045 36436
rect 23691 36476 23733 36485
rect 23691 36436 23692 36476
rect 23732 36436 23733 36476
rect 23691 36427 23733 36436
rect 25515 36476 25557 36485
rect 25515 36436 25516 36476
rect 25556 36436 25557 36476
rect 25515 36427 25557 36436
rect 34819 36476 34877 36477
rect 34819 36436 34828 36476
rect 34868 36436 34877 36476
rect 34819 36435 34877 36436
rect 35779 36476 35837 36477
rect 35779 36436 35788 36476
rect 35828 36436 35837 36476
rect 35779 36435 35837 36436
rect 40867 36476 40925 36477
rect 40867 36436 40876 36476
rect 40916 36436 40925 36476
rect 40867 36435 40925 36436
rect 45099 36476 45141 36485
rect 45099 36436 45100 36476
rect 45140 36436 45141 36476
rect 45099 36427 45141 36436
rect 45483 36476 45525 36485
rect 45483 36436 45484 36476
rect 45524 36436 45525 36476
rect 45483 36427 45525 36436
rect 576 36308 83328 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 83328 36308
rect 576 36244 83328 36268
rect 18891 36140 18933 36149
rect 18891 36100 18892 36140
rect 18932 36100 18933 36140
rect 18891 36091 18933 36100
rect 21867 36140 21909 36149
rect 21867 36100 21868 36140
rect 21908 36100 21909 36140
rect 21867 36091 21909 36100
rect 24835 36140 24893 36141
rect 24835 36100 24844 36140
rect 24884 36100 24893 36140
rect 24835 36099 24893 36100
rect 28003 36140 28061 36141
rect 28003 36100 28012 36140
rect 28052 36100 28061 36140
rect 28003 36099 28061 36100
rect 32227 36140 32285 36141
rect 32227 36100 32236 36140
rect 32276 36100 32285 36140
rect 32227 36099 32285 36100
rect 39139 36140 39197 36141
rect 39139 36100 39148 36140
rect 39188 36100 39197 36140
rect 39139 36099 39197 36100
rect 14851 36056 14909 36057
rect 14851 36016 14860 36056
rect 14900 36016 14909 36056
rect 14851 36015 14909 36016
rect 20419 36056 20477 36057
rect 20419 36016 20428 36056
rect 20468 36016 20477 36056
rect 20419 36015 20477 36016
rect 40195 36056 40253 36057
rect 40195 36016 40204 36056
rect 40244 36016 40253 36056
rect 40195 36015 40253 36016
rect 44227 36056 44285 36057
rect 44227 36016 44236 36056
rect 44276 36016 44285 36056
rect 44227 36015 44285 36016
rect 47979 36056 48021 36065
rect 47979 36016 47980 36056
rect 48020 36016 48021 36056
rect 47979 36007 48021 36016
rect 52963 36056 53021 36057
rect 52963 36016 52972 36056
rect 53012 36016 53021 36056
rect 52963 36015 53021 36016
rect 53923 36056 53981 36057
rect 53923 36016 53932 36056
rect 53972 36016 53981 36056
rect 53923 36015 53981 36016
rect 13699 35972 13757 35973
rect 13699 35932 13708 35972
rect 13748 35932 13757 35972
rect 13699 35931 13757 35932
rect 20611 35972 20669 35973
rect 20611 35932 20620 35972
rect 20660 35932 20669 35972
rect 20611 35931 20669 35932
rect 20995 35972 21053 35973
rect 20995 35932 21004 35972
rect 21044 35932 21053 35972
rect 20995 35931 21053 35932
rect 31075 35972 31133 35973
rect 31075 35932 31084 35972
rect 31124 35932 31133 35972
rect 31075 35931 31133 35932
rect 41347 35972 41405 35973
rect 41347 35932 41356 35972
rect 41396 35932 41405 35972
rect 41347 35931 41405 35932
rect 14179 35888 14237 35889
rect 14179 35848 14188 35888
rect 14228 35848 14237 35888
rect 14179 35847 14237 35848
rect 14475 35888 14517 35897
rect 14475 35848 14476 35888
rect 14516 35848 14517 35888
rect 14475 35839 14517 35848
rect 15243 35888 15285 35897
rect 15243 35848 15244 35888
rect 15284 35848 15285 35888
rect 15243 35839 15285 35848
rect 15619 35888 15677 35889
rect 15619 35848 15628 35888
rect 15668 35848 15677 35888
rect 15619 35847 15677 35848
rect 16483 35888 16541 35889
rect 16483 35848 16492 35888
rect 16532 35848 16541 35888
rect 16483 35847 16541 35848
rect 19179 35888 19221 35897
rect 19179 35848 19180 35888
rect 19220 35848 19221 35888
rect 19179 35839 19221 35848
rect 19267 35888 19325 35889
rect 19267 35848 19276 35888
rect 19316 35848 19325 35888
rect 19267 35847 19325 35848
rect 19747 35888 19805 35889
rect 19747 35848 19756 35888
rect 19796 35848 19805 35888
rect 19747 35847 19805 35848
rect 20043 35888 20085 35897
rect 20043 35848 20044 35888
rect 20084 35848 20085 35888
rect 20043 35839 20085 35848
rect 21571 35888 21629 35889
rect 21571 35848 21580 35888
rect 21620 35848 21629 35888
rect 21571 35847 21629 35848
rect 21675 35888 21717 35897
rect 21675 35848 21676 35888
rect 21716 35848 21717 35888
rect 21675 35839 21717 35848
rect 21859 35888 21917 35889
rect 21859 35848 21868 35888
rect 21908 35848 21917 35888
rect 21859 35847 21917 35848
rect 22443 35888 22485 35897
rect 22443 35848 22444 35888
rect 22484 35848 22485 35888
rect 22443 35839 22485 35848
rect 22819 35888 22877 35889
rect 22819 35848 22828 35888
rect 22868 35848 22877 35888
rect 22819 35847 22877 35848
rect 23683 35888 23741 35889
rect 23683 35848 23692 35888
rect 23732 35848 23741 35888
rect 23683 35847 23741 35848
rect 25987 35888 26045 35889
rect 25987 35848 25996 35888
rect 26036 35848 26045 35888
rect 25987 35847 26045 35848
rect 26851 35888 26909 35889
rect 26851 35848 26860 35888
rect 26900 35848 26909 35888
rect 26851 35847 26909 35848
rect 31555 35888 31613 35889
rect 31555 35848 31564 35888
rect 31604 35848 31613 35888
rect 31555 35847 31613 35848
rect 31851 35888 31893 35897
rect 31851 35848 31852 35888
rect 31892 35848 31893 35888
rect 31851 35839 31893 35848
rect 34435 35888 34493 35889
rect 34435 35848 34444 35888
rect 34484 35848 34493 35888
rect 34435 35847 34493 35848
rect 35779 35888 35837 35889
rect 35779 35848 35788 35888
rect 35828 35848 35837 35888
rect 35779 35847 35837 35848
rect 36643 35888 36701 35889
rect 36643 35848 36652 35888
rect 36692 35848 36701 35888
rect 36643 35847 36701 35848
rect 38467 35888 38525 35889
rect 38467 35848 38476 35888
rect 38516 35848 38525 35888
rect 38467 35847 38525 35848
rect 38763 35888 38805 35897
rect 38763 35848 38764 35888
rect 38804 35848 38805 35888
rect 38763 35839 38805 35848
rect 38859 35888 38901 35897
rect 38859 35848 38860 35888
rect 38900 35848 38901 35888
rect 38859 35839 38901 35848
rect 39523 35888 39581 35889
rect 39523 35848 39532 35888
rect 39572 35848 39581 35888
rect 39523 35847 39581 35848
rect 39819 35888 39861 35897
rect 39819 35848 39820 35888
rect 39860 35848 39861 35888
rect 39819 35839 39861 35848
rect 39915 35888 39957 35897
rect 39915 35848 39916 35888
rect 39956 35848 39957 35888
rect 39915 35839 39957 35848
rect 41827 35888 41885 35889
rect 41827 35848 41836 35888
rect 41876 35848 41885 35888
rect 41827 35847 41885 35848
rect 42123 35888 42165 35897
rect 42123 35848 42124 35888
rect 42164 35848 42165 35888
rect 42123 35839 42165 35848
rect 42219 35888 42261 35897
rect 42219 35848 42220 35888
rect 42260 35848 42261 35888
rect 42219 35839 42261 35848
rect 43555 35888 43613 35889
rect 43555 35848 43564 35888
rect 43604 35848 43613 35888
rect 43555 35847 43613 35848
rect 43851 35888 43893 35897
rect 43851 35848 43852 35888
rect 43892 35848 43893 35888
rect 43851 35839 43893 35848
rect 44427 35888 44469 35897
rect 44427 35848 44428 35888
rect 44468 35848 44469 35888
rect 44427 35839 44469 35848
rect 44803 35888 44861 35889
rect 44803 35848 44812 35888
rect 44852 35848 44861 35888
rect 44803 35847 44861 35848
rect 45667 35888 45725 35889
rect 45667 35848 45676 35888
rect 45716 35848 45725 35888
rect 45667 35847 45725 35848
rect 49507 35888 49565 35889
rect 49507 35848 49516 35888
rect 49556 35848 49565 35888
rect 49507 35847 49565 35848
rect 52291 35888 52349 35889
rect 52291 35848 52300 35888
rect 52340 35848 52349 35888
rect 52291 35847 52349 35848
rect 52587 35888 52629 35897
rect 52587 35848 52588 35888
rect 52628 35848 52629 35888
rect 52587 35839 52629 35848
rect 53251 35888 53309 35889
rect 53251 35848 53260 35888
rect 53300 35848 53309 35888
rect 53251 35847 53309 35848
rect 53547 35888 53589 35897
rect 53547 35848 53548 35888
rect 53588 35848 53589 35888
rect 53547 35839 53589 35848
rect 72267 35888 72309 35897
rect 72267 35848 72268 35888
rect 72308 35848 72309 35888
rect 72267 35839 72309 35848
rect 14571 35804 14613 35813
rect 14571 35764 14572 35804
rect 14612 35764 14613 35804
rect 14571 35755 14613 35764
rect 20139 35804 20181 35813
rect 20139 35764 20140 35804
rect 20180 35764 20181 35804
rect 20139 35755 20181 35764
rect 25611 35804 25653 35813
rect 25611 35764 25612 35804
rect 25652 35764 25653 35804
rect 25611 35755 25653 35764
rect 31947 35804 31989 35813
rect 31947 35764 31948 35804
rect 31988 35764 31989 35804
rect 31947 35755 31989 35764
rect 35403 35804 35445 35813
rect 35403 35764 35404 35804
rect 35444 35764 35445 35804
rect 35403 35755 35445 35764
rect 43947 35804 43989 35813
rect 43947 35764 43948 35804
rect 43988 35764 43989 35804
rect 43947 35755 43989 35764
rect 52683 35804 52725 35813
rect 52683 35764 52684 35804
rect 52724 35764 52725 35804
rect 52683 35755 52725 35764
rect 53643 35804 53685 35813
rect 53643 35764 53644 35804
rect 53684 35764 53685 35804
rect 53643 35755 53685 35764
rect 13899 35720 13941 35729
rect 13899 35680 13900 35720
rect 13940 35680 13941 35720
rect 13899 35671 13941 35680
rect 17635 35720 17693 35721
rect 17635 35680 17644 35720
rect 17684 35680 17693 35720
rect 17635 35679 17693 35680
rect 19371 35716 19413 35725
rect 19371 35676 19372 35716
rect 19412 35676 19413 35716
rect 19371 35667 19413 35676
rect 20811 35720 20853 35729
rect 20811 35680 20812 35720
rect 20852 35680 20853 35720
rect 20811 35671 20853 35680
rect 21195 35720 21237 35729
rect 21195 35680 21196 35720
rect 21236 35680 21237 35720
rect 21195 35671 21237 35680
rect 31275 35720 31317 35729
rect 31275 35680 31276 35720
rect 31316 35680 31317 35720
rect 31275 35671 31317 35680
rect 32907 35720 32949 35729
rect 32907 35680 32908 35720
rect 32948 35680 32949 35720
rect 32907 35671 32949 35680
rect 37795 35720 37853 35721
rect 37795 35680 37804 35720
rect 37844 35680 37853 35720
rect 37795 35679 37853 35680
rect 41547 35720 41589 35729
rect 41547 35680 41548 35720
rect 41588 35680 41589 35720
rect 46819 35720 46877 35721
rect 41547 35671 41589 35680
rect 42507 35678 42549 35687
rect 46819 35680 46828 35720
rect 46868 35680 46877 35720
rect 46819 35679 46877 35680
rect 72651 35720 72693 35729
rect 72651 35680 72652 35720
rect 72692 35680 72693 35720
rect 42507 35638 42508 35678
rect 42548 35638 42549 35678
rect 72651 35671 72693 35680
rect 42507 35629 42549 35638
rect 576 35552 83328 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 83328 35552
rect 576 35488 83328 35512
rect 17451 35384 17493 35393
rect 17451 35344 17452 35384
rect 17492 35344 17493 35384
rect 17451 35335 17493 35344
rect 21571 35384 21629 35385
rect 21571 35344 21580 35384
rect 21620 35344 21629 35384
rect 21571 35343 21629 35344
rect 27243 35384 27285 35393
rect 27243 35344 27244 35384
rect 27284 35344 27285 35384
rect 27243 35335 27285 35344
rect 27723 35384 27765 35393
rect 27723 35344 27724 35384
rect 27764 35344 27765 35384
rect 27723 35335 27765 35344
rect 32227 35384 32285 35385
rect 32227 35344 32236 35384
rect 32276 35344 32285 35384
rect 32227 35343 32285 35344
rect 43555 35384 43613 35385
rect 43555 35344 43564 35384
rect 43604 35344 43613 35384
rect 43555 35343 43613 35344
rect 18699 35300 18741 35309
rect 18699 35260 18700 35300
rect 18740 35260 18741 35300
rect 18699 35251 18741 35260
rect 28395 35300 28437 35309
rect 28395 35260 28396 35300
rect 28436 35260 28437 35300
rect 28395 35251 28437 35260
rect 29355 35300 29397 35309
rect 29355 35260 29356 35300
rect 29396 35260 29397 35300
rect 29355 35251 29397 35260
rect 44043 35300 44085 35309
rect 44043 35260 44044 35300
rect 44084 35260 44085 35300
rect 44043 35251 44085 35260
rect 53163 35300 53205 35309
rect 53163 35260 53164 35300
rect 53204 35260 53205 35300
rect 53163 35251 53205 35260
rect 13411 35216 13469 35217
rect 13411 35176 13420 35216
rect 13460 35176 13469 35216
rect 13411 35175 13469 35176
rect 13707 35216 13749 35225
rect 13707 35176 13708 35216
rect 13748 35176 13749 35216
rect 13707 35167 13749 35176
rect 13803 35216 13845 35225
rect 13803 35176 13804 35216
rect 13844 35176 13845 35216
rect 13803 35167 13845 35176
rect 14283 35216 14325 35225
rect 14283 35176 14284 35216
rect 14324 35176 14325 35216
rect 14283 35167 14325 35176
rect 14659 35216 14717 35217
rect 14659 35176 14668 35216
rect 14708 35176 14717 35216
rect 14659 35175 14717 35176
rect 15523 35216 15581 35217
rect 15523 35176 15532 35216
rect 15572 35176 15581 35216
rect 15523 35175 15581 35176
rect 17067 35216 17109 35225
rect 17067 35176 17068 35216
rect 17108 35176 17109 35216
rect 17067 35167 17109 35176
rect 18307 35216 18365 35217
rect 18307 35176 18316 35216
rect 18356 35176 18365 35216
rect 18307 35175 18365 35176
rect 18603 35216 18645 35225
rect 18603 35176 18604 35216
rect 18644 35176 18645 35216
rect 18603 35167 18645 35176
rect 19179 35216 19221 35225
rect 19179 35176 19180 35216
rect 19220 35176 19221 35216
rect 19179 35167 19221 35176
rect 19555 35216 19613 35217
rect 19555 35176 19564 35216
rect 19604 35176 19613 35216
rect 19555 35175 19613 35176
rect 20419 35216 20477 35217
rect 20419 35176 20428 35216
rect 20468 35176 20477 35216
rect 20419 35175 20477 35176
rect 24459 35216 24501 35225
rect 24459 35176 24460 35216
rect 24500 35176 24501 35216
rect 24459 35167 24501 35176
rect 25707 35216 25749 35225
rect 25707 35176 25708 35216
rect 25748 35176 25749 35216
rect 25707 35167 25749 35176
rect 26755 35216 26813 35217
rect 26755 35176 26764 35216
rect 26804 35176 26813 35216
rect 26755 35175 26813 35176
rect 27043 35216 27101 35217
rect 27043 35176 27052 35216
rect 27092 35176 27101 35216
rect 27043 35175 27101 35176
rect 28003 35216 28061 35217
rect 28003 35176 28012 35216
rect 28052 35176 28061 35216
rect 28003 35175 28061 35176
rect 28299 35216 28341 35225
rect 28299 35176 28300 35216
rect 28340 35176 28341 35216
rect 28299 35167 28341 35176
rect 28963 35216 29021 35217
rect 28963 35176 28972 35216
rect 29012 35176 29021 35216
rect 28963 35175 29021 35176
rect 29259 35216 29301 35225
rect 29259 35176 29260 35216
rect 29300 35176 29301 35216
rect 29259 35167 29301 35176
rect 29835 35216 29877 35225
rect 29835 35176 29836 35216
rect 29876 35176 29877 35216
rect 29835 35167 29877 35176
rect 30211 35216 30269 35217
rect 30211 35176 30220 35216
rect 30260 35176 30269 35216
rect 30211 35175 30269 35176
rect 31075 35216 31133 35217
rect 31075 35176 31084 35216
rect 31124 35176 31133 35216
rect 31075 35175 31133 35176
rect 33475 35216 33533 35217
rect 33475 35176 33484 35216
rect 33524 35176 33533 35216
rect 33475 35175 33533 35176
rect 34635 35216 34677 35225
rect 34635 35176 34636 35216
rect 34676 35176 34677 35216
rect 34635 35167 34677 35176
rect 35011 35216 35069 35217
rect 35011 35176 35020 35216
rect 35060 35176 35069 35216
rect 35011 35175 35069 35176
rect 35875 35216 35933 35217
rect 35875 35176 35884 35216
rect 35924 35176 35933 35216
rect 35875 35175 35933 35176
rect 37611 35216 37653 35225
rect 37611 35176 37612 35216
rect 37652 35176 37653 35216
rect 37611 35167 37653 35176
rect 38755 35216 38813 35217
rect 38755 35176 38764 35216
rect 38804 35176 38813 35216
rect 38755 35175 38813 35176
rect 39051 35216 39093 35225
rect 39051 35176 39052 35216
rect 39092 35176 39093 35216
rect 39051 35167 39093 35176
rect 39147 35216 39189 35225
rect 39147 35176 39148 35216
rect 39188 35176 39189 35216
rect 39147 35167 39189 35176
rect 40395 35216 40437 35225
rect 40395 35176 40396 35216
rect 40436 35176 40437 35216
rect 40395 35167 40437 35176
rect 40587 35216 40629 35225
rect 40587 35176 40588 35216
rect 40628 35176 40629 35216
rect 40587 35167 40629 35176
rect 40779 35216 40821 35225
rect 40779 35176 40780 35216
rect 40820 35176 40821 35216
rect 40779 35167 40821 35176
rect 41155 35216 41213 35217
rect 41155 35176 41164 35216
rect 41204 35176 41213 35216
rect 41155 35175 41213 35176
rect 42019 35216 42077 35217
rect 42019 35176 42028 35216
rect 42068 35176 42077 35216
rect 42019 35175 42077 35176
rect 43467 35216 43509 35225
rect 43467 35176 43468 35216
rect 43508 35176 43509 35216
rect 43467 35167 43509 35176
rect 43659 35216 43701 35225
rect 43659 35176 43660 35216
rect 43700 35176 43701 35216
rect 43659 35167 43701 35176
rect 43747 35216 43805 35217
rect 43747 35176 43756 35216
rect 43796 35176 43805 35216
rect 43747 35175 43805 35176
rect 44419 35216 44477 35217
rect 44419 35176 44428 35216
rect 44468 35176 44477 35216
rect 44419 35175 44477 35176
rect 45283 35216 45341 35217
rect 45283 35176 45292 35216
rect 45332 35176 45341 35216
rect 45283 35175 45341 35176
rect 46723 35216 46781 35217
rect 46723 35176 46732 35216
rect 46772 35176 46781 35216
rect 46723 35175 46781 35176
rect 47019 35216 47061 35225
rect 47019 35176 47020 35216
rect 47060 35176 47061 35216
rect 47019 35167 47061 35176
rect 47115 35216 47157 35225
rect 47115 35176 47116 35216
rect 47156 35176 47157 35216
rect 47115 35167 47157 35176
rect 47979 35216 48021 35225
rect 47979 35176 47980 35216
rect 48020 35176 48021 35216
rect 47979 35167 48021 35176
rect 48355 35216 48413 35217
rect 48355 35176 48364 35216
rect 48404 35176 48413 35216
rect 48355 35175 48413 35176
rect 49219 35216 49277 35217
rect 49219 35176 49228 35216
rect 49268 35176 49277 35216
rect 49219 35175 49277 35176
rect 50571 35216 50613 35225
rect 50571 35176 50572 35216
rect 50612 35176 50613 35216
rect 50571 35167 50613 35176
rect 50947 35216 51005 35217
rect 50947 35176 50956 35216
rect 50996 35176 51005 35216
rect 50947 35175 51005 35176
rect 51811 35216 51869 35217
rect 51811 35176 51820 35216
rect 51860 35176 51869 35216
rect 51811 35175 51869 35176
rect 53539 35216 53597 35217
rect 53539 35176 53548 35216
rect 53588 35176 53597 35216
rect 53539 35175 53597 35176
rect 54403 35216 54461 35217
rect 54403 35176 54412 35216
rect 54452 35176 54461 35216
rect 54403 35175 54461 35176
rect 12259 35132 12317 35133
rect 12259 35092 12268 35132
rect 12308 35092 12317 35132
rect 12259 35091 12317 35092
rect 27523 35132 27581 35133
rect 27523 35092 27532 35132
rect 27572 35092 27581 35132
rect 27523 35091 27581 35092
rect 47587 35132 47645 35133
rect 47587 35092 47596 35132
rect 47636 35092 47645 35132
rect 47587 35091 47645 35092
rect 14083 35048 14141 35049
rect 14083 35008 14092 35048
rect 14132 35008 14141 35048
rect 14083 35007 14141 35008
rect 18979 35048 19037 35049
rect 18979 35008 18988 35048
rect 19028 35008 19037 35048
rect 18979 35007 19037 35008
rect 29635 35048 29693 35049
rect 29635 35008 29644 35048
rect 29684 35008 29693 35048
rect 29635 35007 29693 35008
rect 12459 34964 12501 34973
rect 12459 34924 12460 34964
rect 12500 34924 12501 34964
rect 12459 34915 12501 34924
rect 16675 34964 16733 34965
rect 16675 34924 16684 34964
rect 16724 34924 16733 34964
rect 16675 34923 16733 34924
rect 17643 34964 17685 34973
rect 17643 34924 17644 34964
rect 17684 34924 17685 34964
rect 17643 34915 17685 34924
rect 24843 34964 24885 34973
rect 24843 34924 24844 34964
rect 24884 34924 24885 34964
rect 24843 34915 24885 34924
rect 26091 34964 26133 34973
rect 26091 34924 26092 34964
rect 26132 34924 26133 34964
rect 26091 34915 26133 34924
rect 28675 34964 28733 34965
rect 28675 34924 28684 34964
rect 28724 34924 28733 34964
rect 28675 34923 28733 34924
rect 32227 34964 32285 34965
rect 32227 34924 32236 34964
rect 32276 34924 32285 34964
rect 32227 34923 32285 34924
rect 33771 34964 33813 34973
rect 33771 34924 33772 34964
rect 33812 34924 33813 34964
rect 33771 34915 33813 34924
rect 37027 34964 37085 34965
rect 37027 34924 37036 34964
rect 37076 34924 37085 34964
rect 37027 34923 37085 34924
rect 37803 34964 37845 34973
rect 37803 34924 37804 34964
rect 37844 34924 37845 34964
rect 37803 34915 37845 34924
rect 39427 34964 39485 34965
rect 39427 34924 39436 34964
rect 39476 34924 39485 34964
rect 39427 34923 39485 34924
rect 40587 34964 40629 34973
rect 40587 34924 40588 34964
rect 40628 34924 40629 34964
rect 40587 34915 40629 34924
rect 43171 34964 43229 34965
rect 43171 34924 43180 34964
rect 43220 34924 43229 34964
rect 43171 34923 43229 34924
rect 46435 34964 46493 34965
rect 46435 34924 46444 34964
rect 46484 34924 46493 34964
rect 46435 34923 46493 34924
rect 47395 34964 47453 34965
rect 47395 34924 47404 34964
rect 47444 34924 47453 34964
rect 47395 34923 47453 34924
rect 47787 34964 47829 34973
rect 47787 34924 47788 34964
rect 47828 34924 47829 34964
rect 47787 34915 47829 34924
rect 50371 34964 50429 34965
rect 50371 34924 50380 34964
rect 50420 34924 50429 34964
rect 50371 34923 50429 34924
rect 52963 34964 53021 34965
rect 52963 34924 52972 34964
rect 53012 34924 53021 34964
rect 52963 34923 53021 34924
rect 55555 34964 55613 34965
rect 55555 34924 55564 34964
rect 55604 34924 55613 34964
rect 55555 34923 55613 34924
rect 576 34796 83328 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 83328 34796
rect 576 34732 83328 34756
rect 20331 34628 20373 34637
rect 20331 34588 20332 34628
rect 20372 34588 20373 34628
rect 20331 34579 20373 34588
rect 35491 34628 35549 34629
rect 35491 34588 35500 34628
rect 35540 34588 35549 34628
rect 35491 34587 35549 34588
rect 47203 34628 47261 34629
rect 47203 34588 47212 34628
rect 47252 34588 47261 34628
rect 47203 34587 47261 34588
rect 50755 34628 50813 34629
rect 50755 34588 50764 34628
rect 50804 34588 50813 34628
rect 50755 34587 50813 34588
rect 51915 34628 51957 34637
rect 51915 34588 51916 34628
rect 51956 34588 51957 34628
rect 51915 34579 51957 34588
rect 11587 34544 11645 34545
rect 11587 34504 11596 34544
rect 11636 34504 11645 34544
rect 11587 34503 11645 34504
rect 16291 34544 16349 34545
rect 16291 34504 16300 34544
rect 16340 34504 16349 34544
rect 16291 34503 16349 34504
rect 23395 34544 23453 34545
rect 23395 34504 23404 34544
rect 23444 34504 23453 34544
rect 23395 34503 23453 34504
rect 24451 34544 24509 34545
rect 24451 34504 24460 34544
rect 24500 34504 24509 34544
rect 24451 34503 24509 34504
rect 31939 34544 31997 34545
rect 31939 34504 31948 34544
rect 31988 34504 31997 34544
rect 31939 34503 31997 34504
rect 42891 34544 42933 34553
rect 42891 34504 42892 34544
rect 42932 34504 42933 34544
rect 42891 34495 42933 34504
rect 43371 34544 43413 34553
rect 43371 34504 43372 34544
rect 43412 34504 43413 34544
rect 43371 34495 43413 34504
rect 49795 34544 49853 34545
rect 49795 34504 49804 34544
rect 49844 34504 49853 34544
rect 49795 34503 49853 34504
rect 18891 34460 18933 34469
rect 18891 34420 18892 34460
rect 18932 34420 18933 34460
rect 18891 34411 18933 34420
rect 27051 34460 27093 34469
rect 27051 34420 27052 34460
rect 27092 34420 27093 34460
rect 27051 34411 27093 34420
rect 30411 34460 30453 34469
rect 30411 34420 30412 34460
rect 30452 34420 30453 34460
rect 30411 34411 30453 34420
rect 7371 34376 7413 34385
rect 7371 34336 7372 34376
rect 7412 34336 7413 34376
rect 7371 34327 7413 34336
rect 10915 34376 10973 34377
rect 10915 34336 10924 34376
rect 10964 34336 10973 34376
rect 10915 34335 10973 34336
rect 11211 34376 11253 34385
rect 11211 34336 11212 34376
rect 11252 34336 11253 34376
rect 11211 34327 11253 34336
rect 11787 34376 11829 34385
rect 11787 34336 11788 34376
rect 11828 34336 11829 34376
rect 11787 34327 11829 34336
rect 12163 34376 12221 34377
rect 12163 34336 12172 34376
rect 12212 34336 12221 34376
rect 12163 34335 12221 34336
rect 13027 34376 13085 34377
rect 13027 34336 13036 34376
rect 13076 34336 13085 34376
rect 13027 34335 13085 34336
rect 15235 34376 15293 34377
rect 15235 34336 15244 34376
rect 15284 34336 15293 34376
rect 15235 34335 15293 34336
rect 15619 34376 15677 34377
rect 15619 34336 15628 34376
rect 15668 34336 15677 34376
rect 15619 34335 15677 34336
rect 15915 34376 15957 34385
rect 15915 34336 15916 34376
rect 15956 34336 15957 34376
rect 15915 34327 15957 34336
rect 16011 34376 16053 34385
rect 16011 34336 16012 34376
rect 16052 34336 16053 34376
rect 16011 34327 16053 34336
rect 16491 34376 16533 34385
rect 16491 34336 16492 34376
rect 16532 34336 16533 34376
rect 16491 34327 16533 34336
rect 16867 34376 16925 34377
rect 16867 34336 16876 34376
rect 16916 34336 16925 34376
rect 16867 34335 16925 34336
rect 17731 34376 17789 34377
rect 17731 34336 17740 34376
rect 17780 34336 17789 34376
rect 17731 34335 17789 34336
rect 19843 34376 19901 34377
rect 19843 34336 19852 34376
rect 19892 34336 19901 34376
rect 19843 34335 19901 34336
rect 20803 34376 20861 34377
rect 20803 34336 20812 34376
rect 20852 34336 20861 34376
rect 20803 34335 20861 34336
rect 21003 34376 21045 34385
rect 21003 34336 21004 34376
rect 21044 34336 21045 34376
rect 21003 34327 21045 34336
rect 21379 34376 21437 34377
rect 21379 34336 21388 34376
rect 21428 34336 21437 34376
rect 21379 34335 21437 34336
rect 22243 34376 22301 34377
rect 22243 34336 22252 34376
rect 22292 34336 22301 34376
rect 22243 34335 22301 34336
rect 23779 34376 23837 34377
rect 23779 34336 23788 34376
rect 23828 34336 23837 34376
rect 23779 34335 23837 34336
rect 24075 34376 24117 34385
rect 24075 34336 24076 34376
rect 24116 34336 24117 34376
rect 24075 34327 24117 34336
rect 24651 34376 24693 34385
rect 24651 34336 24652 34376
rect 24692 34336 24693 34376
rect 24651 34327 24693 34336
rect 25027 34376 25085 34377
rect 25027 34336 25036 34376
rect 25076 34336 25085 34376
rect 25027 34335 25085 34336
rect 25891 34376 25949 34377
rect 25891 34336 25900 34376
rect 25940 34336 25949 34376
rect 25891 34335 25949 34336
rect 28011 34376 28053 34385
rect 28011 34336 28012 34376
rect 28052 34336 28053 34376
rect 28011 34327 28053 34336
rect 28387 34376 28445 34377
rect 28387 34336 28396 34376
rect 28436 34336 28445 34376
rect 28387 34335 28445 34336
rect 29251 34376 29309 34377
rect 29251 34336 29260 34376
rect 29300 34336 29309 34376
rect 29251 34335 29309 34336
rect 31267 34376 31325 34377
rect 31267 34336 31276 34376
rect 31316 34336 31325 34376
rect 31267 34335 31325 34336
rect 31563 34376 31605 34385
rect 31563 34336 31564 34376
rect 31604 34336 31605 34376
rect 31563 34327 31605 34336
rect 32139 34376 32181 34385
rect 32139 34336 32140 34376
rect 32180 34336 32181 34376
rect 32139 34327 32181 34336
rect 32515 34376 32573 34377
rect 32515 34336 32524 34376
rect 32564 34336 32573 34376
rect 32515 34335 32573 34336
rect 33379 34376 33437 34377
rect 33379 34336 33388 34376
rect 33428 34336 33437 34376
rect 33379 34335 33437 34336
rect 34819 34376 34877 34377
rect 34819 34336 34828 34376
rect 34868 34336 34877 34376
rect 34819 34335 34877 34336
rect 35115 34376 35157 34385
rect 35115 34336 35116 34376
rect 35156 34336 35157 34376
rect 35115 34327 35157 34336
rect 37323 34376 37365 34385
rect 37323 34336 37324 34376
rect 37364 34336 37365 34376
rect 37323 34327 37365 34336
rect 37699 34376 37757 34377
rect 37699 34336 37708 34376
rect 37748 34336 37757 34376
rect 37699 34335 37757 34336
rect 38563 34376 38621 34377
rect 38563 34336 38572 34376
rect 38612 34336 38621 34376
rect 38563 34335 38621 34336
rect 41067 34376 41109 34385
rect 41067 34336 41068 34376
rect 41108 34336 41109 34376
rect 41067 34327 41109 34336
rect 41259 34376 41301 34385
rect 41259 34336 41260 34376
rect 41300 34336 41301 34376
rect 41259 34327 41301 34336
rect 41347 34376 41405 34377
rect 41347 34336 41356 34376
rect 41396 34336 41405 34376
rect 41347 34335 41405 34336
rect 41643 34376 41685 34385
rect 41643 34336 41644 34376
rect 41684 34336 41685 34376
rect 41643 34327 41685 34336
rect 41835 34376 41877 34385
rect 41835 34336 41836 34376
rect 41876 34336 41877 34376
rect 41835 34327 41877 34336
rect 42211 34376 42269 34377
rect 42211 34336 42220 34376
rect 42260 34336 42269 34376
rect 42211 34335 42269 34336
rect 42699 34376 42741 34385
rect 42699 34336 42700 34376
rect 42740 34336 42741 34376
rect 42699 34327 42741 34336
rect 42891 34376 42933 34385
rect 42891 34336 42892 34376
rect 42932 34336 42933 34376
rect 42891 34327 42933 34336
rect 43755 34376 43797 34385
rect 43755 34336 43756 34376
rect 43796 34336 43797 34376
rect 43755 34327 43797 34336
rect 45187 34376 45245 34377
rect 45187 34336 45196 34376
rect 45236 34336 45245 34376
rect 45187 34335 45245 34336
rect 46531 34376 46589 34377
rect 46531 34336 46540 34376
rect 46580 34336 46589 34376
rect 46531 34335 46589 34336
rect 46827 34376 46869 34385
rect 46827 34336 46828 34376
rect 46868 34336 46869 34376
rect 46827 34327 46869 34336
rect 46923 34376 46965 34385
rect 46923 34336 46924 34376
rect 46964 34336 46965 34376
rect 46923 34327 46965 34336
rect 47403 34376 47445 34385
rect 47403 34336 47404 34376
rect 47444 34336 47445 34376
rect 47403 34327 47445 34336
rect 47779 34376 47837 34377
rect 47779 34336 47788 34376
rect 47828 34336 47837 34376
rect 47779 34335 47837 34336
rect 48643 34376 48701 34377
rect 48643 34336 48652 34376
rect 48692 34336 48701 34376
rect 48643 34335 48701 34336
rect 50083 34376 50141 34377
rect 50083 34336 50092 34376
rect 50132 34336 50141 34376
rect 50083 34335 50141 34336
rect 50379 34376 50421 34385
rect 50379 34336 50380 34376
rect 50420 34336 50421 34376
rect 50379 34327 50421 34336
rect 51531 34376 51573 34385
rect 51531 34336 51532 34376
rect 51572 34336 51573 34376
rect 51531 34327 51573 34336
rect 52779 34376 52821 34385
rect 52779 34336 52780 34376
rect 52820 34336 52821 34376
rect 52779 34327 52821 34336
rect 53635 34376 53693 34377
rect 53635 34336 53644 34376
rect 53684 34336 53693 34376
rect 53635 34335 53693 34336
rect 54123 34376 54165 34385
rect 54123 34336 54124 34376
rect 54164 34336 54165 34376
rect 54123 34327 54165 34336
rect 54499 34376 54557 34377
rect 54499 34336 54508 34376
rect 54548 34336 54557 34376
rect 54499 34335 54557 34336
rect 55363 34376 55421 34377
rect 55363 34336 55372 34376
rect 55412 34336 55421 34376
rect 55363 34335 55421 34336
rect 61507 34376 61565 34377
rect 61507 34336 61516 34376
rect 61556 34336 61565 34376
rect 61507 34335 61565 34336
rect 62467 34376 62525 34377
rect 62467 34336 62476 34376
rect 62516 34336 62525 34376
rect 62467 34335 62525 34336
rect 63339 34376 63381 34385
rect 63339 34336 63340 34376
rect 63380 34336 63381 34376
rect 63339 34327 63381 34336
rect 64675 34376 64733 34377
rect 64675 34336 64684 34376
rect 64724 34336 64733 34376
rect 64675 34335 64733 34336
rect 65923 34376 65981 34377
rect 65923 34336 65932 34376
rect 65972 34336 65981 34376
rect 65923 34335 65981 34336
rect 66883 34376 66941 34377
rect 66883 34336 66892 34376
rect 66932 34336 66941 34376
rect 66883 34335 66941 34336
rect 81187 34376 81245 34377
rect 81187 34336 81196 34376
rect 81236 34336 81245 34376
rect 81187 34335 81245 34336
rect 82051 34376 82109 34377
rect 82051 34336 82060 34376
rect 82100 34336 82109 34376
rect 82051 34335 82109 34336
rect 11307 34292 11349 34301
rect 11307 34252 11308 34292
rect 11348 34252 11349 34292
rect 11307 34243 11349 34252
rect 24171 34292 24213 34301
rect 24171 34252 24172 34292
rect 24212 34252 24213 34292
rect 24171 34243 24213 34252
rect 31659 34292 31701 34301
rect 31659 34252 31660 34292
rect 31700 34252 31701 34292
rect 31659 34243 31701 34252
rect 35211 34292 35253 34301
rect 35211 34252 35212 34292
rect 35252 34252 35253 34292
rect 35211 34243 35253 34252
rect 41163 34292 41205 34301
rect 41163 34252 41164 34292
rect 41204 34252 41205 34292
rect 41163 34243 41205 34252
rect 50475 34292 50517 34301
rect 50475 34252 50476 34292
rect 50516 34252 50517 34292
rect 50475 34243 50517 34252
rect 80811 34292 80853 34301
rect 80811 34252 80812 34292
rect 80852 34252 80853 34292
rect 80811 34243 80853 34252
rect 7755 34208 7797 34217
rect 7755 34168 7756 34208
rect 7796 34168 7797 34208
rect 7755 34159 7797 34168
rect 14179 34208 14237 34209
rect 14179 34168 14188 34208
rect 14228 34168 14237 34208
rect 14179 34167 14237 34168
rect 34531 34208 34589 34209
rect 34531 34168 34540 34208
rect 34580 34168 34589 34208
rect 34531 34167 34589 34168
rect 39715 34208 39773 34209
rect 39715 34168 39724 34208
rect 39764 34168 39773 34208
rect 39715 34167 39773 34168
rect 41739 34208 41781 34217
rect 41739 34168 41740 34208
rect 41780 34168 41781 34208
rect 41739 34159 41781 34168
rect 42315 34208 42357 34217
rect 42315 34168 42316 34208
rect 42356 34168 42357 34208
rect 42315 34159 42357 34168
rect 56515 34208 56573 34209
rect 56515 34168 56524 34208
rect 56564 34168 56573 34208
rect 56515 34167 56573 34168
rect 83203 34208 83261 34209
rect 83203 34168 83212 34208
rect 83252 34168 83261 34208
rect 83203 34167 83261 34168
rect 576 34040 83328 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 83328 34040
rect 576 33976 83328 34000
rect 80139 33788 80181 33797
rect 80139 33748 80140 33788
rect 80180 33748 80181 33788
rect 80139 33739 80181 33748
rect 79747 33704 79805 33705
rect 79747 33664 79756 33704
rect 79796 33664 79805 33704
rect 79747 33663 79805 33664
rect 80043 33704 80085 33713
rect 80043 33664 80044 33704
rect 80084 33664 80085 33704
rect 80043 33655 80085 33664
rect 80707 33704 80765 33705
rect 80707 33664 80716 33704
rect 80756 33664 80765 33704
rect 80707 33663 80765 33664
rect 81003 33704 81045 33713
rect 81003 33664 81004 33704
rect 81044 33664 81045 33704
rect 81003 33655 81045 33664
rect 81099 33704 81141 33713
rect 81099 33664 81100 33704
rect 81140 33664 81141 33704
rect 81099 33655 81141 33664
rect 81763 33620 81821 33621
rect 81763 33580 81772 33620
rect 81812 33580 81821 33620
rect 81763 33579 81821 33580
rect 80419 33536 80477 33537
rect 80419 33496 80428 33536
rect 80468 33496 80477 33536
rect 80419 33495 80477 33496
rect 81379 33452 81437 33453
rect 81379 33412 81388 33452
rect 81428 33412 81437 33452
rect 81379 33411 81437 33412
rect 81963 33452 82005 33461
rect 81963 33412 81964 33452
rect 82004 33412 82005 33452
rect 81963 33403 82005 33412
rect 576 33284 5952 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 5952 33284
rect 576 33220 5952 33244
rect 74016 33284 83328 33308
rect 74016 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 83328 33284
rect 74016 33220 83328 33244
rect 5643 33116 5685 33125
rect 5643 33076 5644 33116
rect 5684 33076 5685 33116
rect 5643 33067 5685 33076
rect 5443 32948 5501 32949
rect 5443 32908 5452 32948
rect 5492 32908 5501 32948
rect 5443 32907 5501 32908
rect 80419 32948 80477 32949
rect 80419 32908 80428 32948
rect 80468 32908 80477 32948
rect 80419 32907 80477 32908
rect 80811 32864 80853 32873
rect 80811 32824 80812 32864
rect 80852 32824 80853 32864
rect 80811 32815 80853 32824
rect 81187 32864 81245 32865
rect 81187 32824 81196 32864
rect 81236 32824 81245 32864
rect 81187 32823 81245 32824
rect 82051 32864 82109 32865
rect 82051 32824 82060 32864
rect 82100 32824 82109 32864
rect 82051 32823 82109 32824
rect 5643 32696 5685 32705
rect 5643 32656 5644 32696
rect 5684 32656 5685 32696
rect 5643 32647 5685 32656
rect 80619 32696 80661 32705
rect 80619 32656 80620 32696
rect 80660 32656 80661 32696
rect 80619 32647 80661 32656
rect 83203 32696 83261 32697
rect 83203 32656 83212 32696
rect 83252 32656 83261 32696
rect 83203 32655 83261 32656
rect 576 32528 5952 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 5952 32528
rect 576 32464 5952 32488
rect 74016 32528 83328 32552
rect 74016 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 83328 32528
rect 74016 32464 83328 32488
rect 83203 32360 83261 32361
rect 83203 32320 83212 32360
rect 83252 32320 83261 32360
rect 83203 32319 83261 32320
rect 4971 32192 5013 32201
rect 4971 32152 4972 32192
rect 5012 32152 5013 32192
rect 4971 32143 5013 32152
rect 80811 32192 80853 32201
rect 80811 32152 80812 32192
rect 80852 32152 80853 32192
rect 80811 32143 80853 32152
rect 81187 32192 81245 32193
rect 81187 32152 81196 32192
rect 81236 32152 81245 32192
rect 81187 32151 81245 32152
rect 82051 32192 82109 32193
rect 82051 32152 82060 32192
rect 82100 32152 82109 32192
rect 82051 32151 82109 32152
rect 4387 32108 4445 32109
rect 4387 32068 4396 32108
rect 4436 32068 4445 32108
rect 4387 32067 4445 32068
rect 4587 31940 4629 31949
rect 4587 31900 4588 31940
rect 4628 31900 4629 31940
rect 4587 31891 4629 31900
rect 5163 31940 5205 31949
rect 5163 31900 5164 31940
rect 5204 31900 5205 31940
rect 5163 31891 5205 31900
rect 576 31772 5952 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 5952 31772
rect 576 31708 5952 31732
rect 74016 31772 83328 31796
rect 74016 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 83328 31772
rect 74016 31708 83328 31732
rect 81379 31604 81437 31605
rect 81379 31564 81388 31604
rect 81428 31564 81437 31604
rect 81379 31563 81437 31564
rect 5835 31436 5877 31445
rect 5835 31396 5836 31436
rect 5876 31396 5877 31436
rect 5835 31387 5877 31396
rect 81667 31436 81725 31437
rect 81667 31396 81676 31436
rect 81716 31396 81725 31436
rect 81667 31395 81725 31396
rect 3811 31352 3869 31353
rect 3811 31312 3820 31352
rect 3860 31312 3869 31352
rect 3811 31311 3869 31312
rect 4675 31352 4733 31353
rect 4675 31312 4684 31352
rect 4724 31312 4733 31352
rect 4675 31311 4733 31312
rect 80707 31352 80765 31353
rect 80707 31312 80716 31352
rect 80756 31312 80765 31352
rect 80707 31311 80765 31312
rect 81003 31352 81045 31361
rect 81003 31312 81004 31352
rect 81044 31312 81045 31352
rect 81003 31303 81045 31312
rect 81099 31352 81141 31361
rect 81099 31312 81100 31352
rect 81140 31312 81141 31352
rect 81099 31303 81141 31312
rect 3435 31268 3477 31277
rect 3435 31228 3436 31268
rect 3476 31228 3477 31268
rect 3435 31219 3477 31228
rect 81867 31184 81909 31193
rect 81867 31144 81868 31184
rect 81908 31144 81909 31184
rect 81867 31135 81909 31144
rect 576 31016 5952 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 5952 31016
rect 576 30952 5952 30976
rect 74016 31016 83328 31040
rect 74016 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 83328 31016
rect 74016 30952 83328 30976
rect 83203 30848 83261 30849
rect 83203 30808 83212 30848
rect 83252 30808 83261 30848
rect 83203 30807 83261 30808
rect 4875 30764 4917 30773
rect 4875 30724 4876 30764
rect 4916 30724 4917 30764
rect 4875 30715 4917 30724
rect 4483 30680 4541 30681
rect 4483 30640 4492 30680
rect 4532 30640 4541 30680
rect 4483 30639 4541 30640
rect 4779 30680 4821 30689
rect 4779 30640 4780 30680
rect 4820 30640 4821 30680
rect 4779 30631 4821 30640
rect 80811 30680 80853 30689
rect 80811 30640 80812 30680
rect 80852 30640 80853 30680
rect 80811 30631 80853 30640
rect 81187 30680 81245 30681
rect 81187 30640 81196 30680
rect 81236 30640 81245 30680
rect 81187 30639 81245 30640
rect 82051 30680 82109 30681
rect 82051 30640 82060 30680
rect 82100 30640 82109 30680
rect 82051 30639 82109 30640
rect 79939 30596 79997 30597
rect 79939 30556 79948 30596
rect 79988 30556 79997 30596
rect 79939 30555 79997 30556
rect 5155 30512 5213 30513
rect 5155 30472 5164 30512
rect 5204 30472 5213 30512
rect 5155 30471 5213 30472
rect 80139 30428 80181 30437
rect 80139 30388 80140 30428
rect 80180 30388 80181 30428
rect 80139 30379 80181 30388
rect 83203 30428 83261 30429
rect 83203 30388 83212 30428
rect 83252 30388 83261 30428
rect 83203 30387 83261 30388
rect 576 30260 5952 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 5952 30260
rect 576 30196 5952 30220
rect 74016 30260 83328 30284
rect 74016 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 83328 30260
rect 74016 30196 83328 30220
rect 82435 30092 82493 30093
rect 82435 30052 82444 30092
rect 82484 30052 82493 30092
rect 82435 30051 82493 30052
rect 79843 30008 79901 30009
rect 79843 29968 79852 30008
rect 79892 29968 79901 30008
rect 79843 29967 79901 29968
rect 79171 29840 79229 29841
rect 79171 29800 79180 29840
rect 79220 29800 79229 29840
rect 79171 29799 79229 29800
rect 79467 29840 79509 29849
rect 79467 29800 79468 29840
rect 79508 29800 79509 29840
rect 79467 29791 79509 29800
rect 79563 29840 79605 29849
rect 79563 29800 79564 29840
rect 79604 29800 79605 29840
rect 79563 29791 79605 29800
rect 80043 29840 80085 29849
rect 80043 29800 80044 29840
rect 80084 29800 80085 29840
rect 80043 29791 80085 29800
rect 80419 29840 80477 29841
rect 80419 29800 80428 29840
rect 80468 29800 80477 29840
rect 80419 29799 80477 29800
rect 81283 29840 81341 29841
rect 81283 29800 81292 29840
rect 81332 29800 81341 29840
rect 81283 29799 81341 29800
rect 576 29504 5952 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 5952 29504
rect 576 29440 5952 29464
rect 74016 29504 83328 29528
rect 74016 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 83328 29504
rect 74016 29440 83328 29464
rect 80427 29252 80469 29261
rect 80427 29212 80428 29252
rect 80468 29212 80469 29252
rect 80427 29203 80469 29212
rect 80035 29168 80093 29169
rect 80035 29128 80044 29168
rect 80084 29128 80093 29168
rect 80035 29127 80093 29128
rect 80331 29168 80373 29177
rect 80331 29128 80332 29168
rect 80372 29128 80373 29168
rect 80331 29119 80373 29128
rect 80995 29168 81053 29169
rect 80995 29128 81004 29168
rect 81044 29128 81053 29168
rect 80995 29127 81053 29128
rect 81291 29168 81333 29177
rect 81291 29128 81292 29168
rect 81332 29128 81333 29168
rect 81291 29119 81333 29128
rect 81387 29168 81429 29177
rect 81387 29128 81388 29168
rect 81428 29128 81429 29168
rect 81387 29119 81429 29128
rect 80707 29000 80765 29001
rect 80707 28960 80716 29000
rect 80756 28960 80765 29000
rect 80707 28959 80765 28960
rect 81667 28916 81725 28917
rect 81667 28876 81676 28916
rect 81716 28876 81725 28916
rect 81667 28875 81725 28876
rect 576 28748 5952 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 5952 28748
rect 576 28684 5952 28708
rect 74016 28748 83328 28772
rect 74016 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 83328 28748
rect 74016 28684 83328 28708
rect 82627 28580 82685 28581
rect 82627 28540 82636 28580
rect 82676 28540 82685 28580
rect 82627 28539 82685 28540
rect 80035 28496 80093 28497
rect 80035 28456 80044 28496
rect 80084 28456 80093 28496
rect 80035 28455 80093 28456
rect 74763 28328 74805 28337
rect 74763 28288 74764 28328
rect 74804 28288 74805 28328
rect 74763 28279 74805 28288
rect 76099 28328 76157 28329
rect 76099 28288 76108 28328
rect 76148 28288 76157 28328
rect 76099 28287 76157 28288
rect 79363 28328 79421 28329
rect 79363 28288 79372 28328
rect 79412 28288 79421 28328
rect 79363 28287 79421 28288
rect 79659 28328 79701 28337
rect 79659 28288 79660 28328
rect 79700 28288 79701 28328
rect 79659 28279 79701 28288
rect 79755 28328 79797 28337
rect 79755 28288 79756 28328
rect 79796 28288 79797 28328
rect 79755 28279 79797 28288
rect 80235 28328 80277 28337
rect 80235 28288 80236 28328
rect 80276 28288 80277 28328
rect 80235 28279 80277 28288
rect 80611 28328 80669 28329
rect 80611 28288 80620 28328
rect 80660 28288 80669 28328
rect 80611 28287 80669 28288
rect 81475 28328 81533 28329
rect 81475 28288 81484 28328
rect 81524 28288 81533 28328
rect 81475 28287 81533 28288
rect 82627 28160 82685 28161
rect 82627 28120 82636 28160
rect 82676 28120 82685 28160
rect 82627 28119 82685 28120
rect 576 27992 5952 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 5952 27992
rect 576 27928 5952 27952
rect 74016 27992 83328 28016
rect 74016 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 83328 27992
rect 74016 27928 83328 27952
rect 83203 27824 83261 27825
rect 83203 27784 83212 27824
rect 83252 27784 83261 27824
rect 83203 27783 83261 27784
rect 80811 27740 80853 27749
rect 80811 27700 80812 27740
rect 80852 27700 80853 27740
rect 80811 27691 80853 27700
rect 3435 27656 3477 27665
rect 3435 27616 3436 27656
rect 3476 27616 3477 27656
rect 3435 27607 3477 27616
rect 3811 27656 3869 27657
rect 3811 27616 3820 27656
rect 3860 27616 3869 27656
rect 3811 27615 3869 27616
rect 4675 27656 4733 27657
rect 4675 27616 4684 27656
rect 4724 27616 4733 27656
rect 4675 27615 4733 27616
rect 81187 27656 81245 27657
rect 81187 27616 81196 27656
rect 81236 27616 81245 27656
rect 81187 27615 81245 27616
rect 82051 27656 82109 27657
rect 82051 27616 82060 27656
rect 82100 27616 82109 27656
rect 82051 27615 82109 27616
rect 5827 27404 5885 27405
rect 5827 27364 5836 27404
rect 5876 27364 5885 27404
rect 5827 27363 5885 27364
rect 576 27236 5952 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 5952 27236
rect 576 27172 5952 27196
rect 74016 27236 83328 27260
rect 74016 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 83328 27236
rect 74016 27172 83328 27196
rect 5155 27068 5213 27069
rect 5155 27028 5164 27068
rect 5204 27028 5213 27068
rect 5155 27027 5213 27028
rect 82819 27068 82877 27069
rect 82819 27028 82828 27068
rect 82868 27028 82877 27068
rect 82819 27027 82877 27028
rect 4483 26816 4541 26817
rect 4483 26776 4492 26816
rect 4532 26776 4541 26816
rect 4483 26775 4541 26776
rect 4779 26816 4821 26825
rect 4779 26776 4780 26816
rect 4820 26776 4821 26816
rect 4779 26767 4821 26776
rect 80803 26816 80861 26817
rect 80803 26776 80812 26816
rect 80852 26776 80861 26816
rect 80803 26775 80861 26776
rect 81667 26816 81725 26817
rect 81667 26776 81676 26816
rect 81716 26776 81725 26816
rect 81667 26775 81725 26776
rect 4875 26732 4917 26741
rect 4875 26692 4876 26732
rect 4916 26692 4917 26732
rect 4875 26683 4917 26692
rect 80427 26732 80469 26741
rect 80427 26692 80428 26732
rect 80468 26692 80469 26732
rect 80427 26683 80469 26692
rect 576 26480 5952 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 5952 26480
rect 576 26416 5952 26440
rect 74016 26480 83328 26504
rect 74016 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 83328 26480
rect 74016 26416 83328 26440
rect 80619 26228 80661 26237
rect 80619 26188 80620 26228
rect 80660 26188 80661 26228
rect 80619 26179 80661 26188
rect 80227 26144 80285 26145
rect 80227 26104 80236 26144
rect 80276 26104 80285 26144
rect 80227 26103 80285 26104
rect 80523 26144 80565 26153
rect 80523 26104 80524 26144
rect 80564 26104 80565 26144
rect 80523 26095 80565 26104
rect 81283 26144 81341 26145
rect 81283 26104 81292 26144
rect 81332 26104 81341 26144
rect 81283 26103 81341 26104
rect 81579 26144 81621 26153
rect 81579 26104 81580 26144
rect 81620 26104 81621 26144
rect 81579 26095 81621 26104
rect 81675 26144 81717 26153
rect 81675 26104 81676 26144
rect 81716 26104 81717 26144
rect 81675 26095 81717 26104
rect 80899 25976 80957 25977
rect 80899 25936 80908 25976
rect 80948 25936 80957 25976
rect 80899 25935 80957 25936
rect 81955 25892 82013 25893
rect 81955 25852 81964 25892
rect 82004 25852 82013 25892
rect 81955 25851 82013 25852
rect 576 25724 5952 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 5952 25724
rect 576 25660 5952 25684
rect 74016 25724 83328 25748
rect 74016 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 83328 25724
rect 74016 25660 83328 25684
rect 5827 25556 5885 25557
rect 5827 25516 5836 25556
rect 5876 25516 5885 25556
rect 5827 25515 5885 25516
rect 83203 25556 83261 25557
rect 83203 25516 83212 25556
rect 83252 25516 83261 25556
rect 83203 25515 83261 25516
rect 80611 25472 80669 25473
rect 80611 25432 80620 25472
rect 80660 25432 80669 25472
rect 80611 25431 80669 25432
rect 643 25388 701 25389
rect 643 25348 652 25388
rect 692 25348 701 25388
rect 643 25347 701 25348
rect 3811 25304 3869 25305
rect 3811 25264 3820 25304
rect 3860 25264 3869 25304
rect 3811 25263 3869 25264
rect 4675 25304 4733 25305
rect 4675 25264 4684 25304
rect 4724 25264 4733 25304
rect 4675 25263 4733 25264
rect 79939 25304 79997 25305
rect 79939 25264 79948 25304
rect 79988 25264 79997 25304
rect 79939 25263 79997 25264
rect 80235 25304 80277 25313
rect 80235 25264 80236 25304
rect 80276 25264 80277 25304
rect 80235 25255 80277 25264
rect 80811 25304 80853 25313
rect 80811 25264 80812 25304
rect 80852 25264 80853 25304
rect 80811 25255 80853 25264
rect 81187 25304 81245 25305
rect 81187 25264 81196 25304
rect 81236 25264 81245 25304
rect 81187 25263 81245 25264
rect 82051 25304 82109 25305
rect 82051 25264 82060 25304
rect 82100 25264 82109 25304
rect 82051 25263 82109 25264
rect 3435 25220 3477 25229
rect 3435 25180 3436 25220
rect 3476 25180 3477 25220
rect 3435 25171 3477 25180
rect 80331 25220 80373 25229
rect 80331 25180 80332 25220
rect 80372 25180 80373 25220
rect 80331 25171 80373 25180
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 5827 25136 5885 25137
rect 5827 25096 5836 25136
rect 5876 25096 5885 25136
rect 5827 25095 5885 25096
rect 576 24968 5952 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 5952 24968
rect 576 24904 5952 24928
rect 74016 24968 83328 24992
rect 74016 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 83328 24968
rect 74016 24904 83328 24928
rect 5067 24842 5109 24851
rect 5067 24802 5068 24842
rect 5108 24802 5109 24842
rect 5067 24793 5109 24802
rect 4779 24716 4821 24725
rect 4779 24676 4780 24716
rect 4820 24676 4821 24716
rect 4779 24667 4821 24676
rect 80523 24716 80565 24725
rect 80523 24676 80524 24716
rect 80564 24676 80565 24716
rect 80523 24667 80565 24676
rect 4387 24632 4445 24633
rect 4387 24592 4396 24632
rect 4436 24592 4445 24632
rect 4387 24591 4445 24592
rect 4683 24632 4725 24641
rect 4683 24592 4684 24632
rect 4724 24592 4725 24632
rect 4683 24583 4725 24592
rect 74083 24632 74141 24633
rect 74083 24592 74092 24632
rect 74132 24592 74141 24632
rect 74083 24591 74141 24592
rect 80899 24632 80957 24633
rect 80899 24592 80908 24632
rect 80948 24592 80957 24632
rect 80899 24591 80957 24592
rect 81763 24632 81821 24633
rect 81763 24592 81772 24632
rect 81812 24592 81821 24632
rect 81763 24591 81821 24592
rect 643 24548 701 24549
rect 643 24508 652 24548
rect 692 24508 701 24548
rect 643 24507 701 24508
rect 82923 24548 82965 24557
rect 82923 24508 82924 24548
rect 82964 24508 82965 24548
rect 82923 24499 82965 24508
rect 843 24464 885 24473
rect 843 24424 844 24464
rect 884 24424 885 24464
rect 843 24415 885 24424
rect 576 24212 5952 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 5952 24212
rect 576 24148 5952 24172
rect 74016 24212 83328 24236
rect 74016 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 83328 24212
rect 74016 24148 83328 24172
rect 843 24044 885 24053
rect 843 24004 844 24044
rect 884 24004 885 24044
rect 843 23995 885 24004
rect 643 23876 701 23877
rect 643 23836 652 23876
rect 692 23836 701 23876
rect 643 23835 701 23836
rect 74179 23792 74237 23793
rect 74179 23752 74188 23792
rect 74228 23752 74237 23792
rect 74179 23751 74237 23752
rect 74667 23624 74709 23633
rect 74667 23584 74668 23624
rect 74708 23584 74709 23624
rect 74667 23575 74709 23584
rect 576 23456 5952 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 5952 23456
rect 576 23392 5952 23416
rect 74016 23456 83328 23480
rect 74016 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 83328 23456
rect 74016 23392 83328 23416
rect 843 23288 885 23297
rect 843 23248 844 23288
rect 884 23248 885 23288
rect 843 23239 885 23248
rect 3435 23120 3477 23129
rect 3435 23080 3436 23120
rect 3476 23080 3477 23120
rect 3435 23071 3477 23080
rect 3811 23120 3869 23121
rect 3811 23080 3820 23120
rect 3860 23080 3869 23120
rect 3811 23079 3869 23080
rect 4675 23120 4733 23121
rect 4675 23080 4684 23120
rect 4724 23080 4733 23120
rect 4675 23079 4733 23080
rect 74179 23120 74237 23121
rect 74179 23080 74188 23120
rect 74228 23080 74237 23120
rect 74179 23079 74237 23080
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 5827 22868 5885 22869
rect 5827 22828 5836 22868
rect 5876 22828 5885 22868
rect 5827 22827 5885 22828
rect 74475 22868 74517 22877
rect 74475 22828 74476 22868
rect 74516 22828 74517 22868
rect 74475 22819 74517 22828
rect 576 22700 5952 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 5952 22700
rect 576 22636 5952 22660
rect 74016 22700 83328 22724
rect 74016 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 83328 22700
rect 74016 22636 83328 22660
rect 4387 22532 4445 22533
rect 4387 22492 4396 22532
rect 4436 22492 4445 22532
rect 4387 22491 4445 22492
rect 3715 22280 3773 22281
rect 3715 22240 3724 22280
rect 3764 22240 3773 22280
rect 3715 22239 3773 22240
rect 4011 22280 4053 22289
rect 4011 22240 4012 22280
rect 4052 22240 4053 22280
rect 4011 22231 4053 22240
rect 4107 22280 4149 22289
rect 4107 22240 4108 22280
rect 4148 22240 4149 22280
rect 4107 22231 4149 22240
rect 835 22112 893 22113
rect 835 22072 844 22112
rect 884 22072 893 22112
rect 835 22071 893 22072
rect 576 21944 5952 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 5952 21944
rect 576 21880 5952 21904
rect 74016 21944 99360 21968
rect 74016 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 74016 21880 99360 21904
rect 3435 21608 3477 21617
rect 3435 21568 3436 21608
rect 3476 21568 3477 21608
rect 3435 21559 3477 21568
rect 3811 21608 3869 21609
rect 3811 21568 3820 21608
rect 3860 21568 3869 21608
rect 3811 21567 3869 21568
rect 4675 21608 4733 21609
rect 4675 21568 4684 21608
rect 4724 21568 4733 21608
rect 4675 21567 4733 21568
rect 82731 21608 82773 21617
rect 82731 21568 82732 21608
rect 82772 21568 82773 21608
rect 82731 21559 82773 21568
rect 83107 21608 83165 21609
rect 83107 21568 83116 21608
rect 83156 21568 83165 21608
rect 83107 21567 83165 21568
rect 83971 21608 84029 21609
rect 83971 21568 83980 21608
rect 84020 21568 84029 21608
rect 83971 21567 84029 21568
rect 5835 21524 5877 21533
rect 5835 21484 5836 21524
rect 5876 21484 5877 21524
rect 5835 21475 5877 21484
rect 85123 21356 85181 21357
rect 85123 21316 85132 21356
rect 85172 21316 85181 21356
rect 85123 21315 85181 21316
rect 576 21188 5952 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 5952 21188
rect 576 21124 5952 21148
rect 74016 21188 99360 21212
rect 74016 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 74016 21124 99360 21148
rect 82339 21020 82397 21021
rect 82339 20980 82348 21020
rect 82388 20980 82397 21020
rect 82339 20979 82397 20980
rect 2755 20936 2813 20937
rect 2755 20896 2764 20936
rect 2804 20896 2813 20936
rect 2755 20895 2813 20896
rect 2083 20768 2141 20769
rect 2083 20728 2092 20768
rect 2132 20728 2141 20768
rect 2083 20727 2141 20728
rect 2379 20768 2421 20777
rect 2379 20728 2380 20768
rect 2420 20728 2421 20768
rect 2379 20719 2421 20728
rect 2955 20768 2997 20777
rect 2955 20728 2956 20768
rect 2996 20728 2997 20768
rect 2955 20719 2997 20728
rect 3331 20768 3389 20769
rect 3331 20728 3340 20768
rect 3380 20728 3389 20768
rect 3331 20727 3389 20728
rect 4195 20768 4253 20769
rect 4195 20728 4204 20768
rect 4244 20728 4253 20768
rect 4195 20727 4253 20728
rect 81667 20768 81725 20769
rect 81667 20728 81676 20768
rect 81716 20728 81725 20768
rect 81667 20727 81725 20728
rect 81963 20768 82005 20777
rect 81963 20728 81964 20768
rect 82004 20728 82005 20768
rect 81963 20719 82005 20728
rect 82059 20768 82101 20777
rect 82059 20728 82060 20768
rect 82100 20728 82101 20768
rect 82059 20719 82101 20728
rect 2475 20684 2517 20693
rect 2475 20644 2476 20684
rect 2516 20644 2517 20684
rect 2475 20635 2517 20644
rect 835 20600 893 20601
rect 835 20560 844 20600
rect 884 20560 893 20600
rect 835 20559 893 20560
rect 5347 20600 5405 20601
rect 5347 20560 5356 20600
rect 5396 20560 5405 20600
rect 5347 20559 5405 20560
rect 576 20432 5952 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 5952 20432
rect 576 20368 5952 20392
rect 74016 20432 99360 20456
rect 74016 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 74016 20368 99360 20392
rect 835 20264 893 20265
rect 835 20224 844 20264
rect 884 20224 893 20264
rect 835 20223 893 20224
rect 4299 20180 4341 20189
rect 4299 20140 4300 20180
rect 4340 20140 4341 20180
rect 4299 20131 4341 20140
rect 1227 20096 1269 20105
rect 1227 20056 1228 20096
rect 1268 20056 1269 20096
rect 1227 20047 1269 20056
rect 1603 20096 1661 20097
rect 1603 20056 1612 20096
rect 1652 20056 1661 20096
rect 1603 20055 1661 20056
rect 2467 20096 2525 20097
rect 2467 20056 2476 20096
rect 2516 20056 2525 20096
rect 2467 20055 2525 20056
rect 3907 20096 3965 20097
rect 3907 20056 3916 20096
rect 3956 20056 3965 20096
rect 3907 20055 3965 20056
rect 4203 20096 4245 20105
rect 4203 20056 4204 20096
rect 4244 20056 4245 20096
rect 4203 20047 4245 20056
rect 98371 20096 98429 20097
rect 98371 20056 98380 20096
rect 98420 20056 98429 20096
rect 98371 20055 98429 20056
rect 4579 19928 4637 19929
rect 4579 19888 4588 19928
rect 4628 19888 4637 19928
rect 4579 19887 4637 19888
rect 96843 19928 96885 19937
rect 96843 19888 96844 19928
rect 96884 19888 96885 19928
rect 96843 19879 96885 19888
rect 3619 19844 3677 19845
rect 3619 19804 3628 19844
rect 3668 19804 3677 19844
rect 3619 19803 3677 19804
rect 576 19676 5952 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 5952 19676
rect 576 19612 5952 19636
rect 74016 19676 99360 19700
rect 74016 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 74016 19612 99360 19636
rect 2275 19508 2333 19509
rect 2275 19468 2284 19508
rect 2324 19468 2333 19508
rect 2275 19467 2333 19468
rect 5067 19508 5109 19517
rect 5067 19468 5068 19508
rect 5108 19468 5109 19508
rect 5067 19459 5109 19468
rect 4675 19424 4733 19425
rect 4675 19384 4684 19424
rect 4724 19384 4733 19424
rect 4675 19383 4733 19384
rect 2467 19340 2525 19341
rect 2467 19300 2476 19340
rect 2516 19300 2525 19340
rect 2467 19299 2525 19300
rect 3523 19340 3581 19341
rect 3523 19300 3532 19340
rect 3572 19300 3581 19340
rect 3523 19299 3581 19300
rect 4867 19340 4925 19341
rect 4867 19300 4876 19340
rect 4916 19300 4925 19340
rect 4867 19299 4925 19300
rect 1603 19256 1661 19257
rect 1603 19216 1612 19256
rect 1652 19216 1661 19256
rect 1603 19215 1661 19216
rect 1899 19256 1941 19265
rect 1899 19216 1900 19256
rect 1940 19216 1941 19256
rect 1899 19207 1941 19216
rect 1995 19256 2037 19265
rect 1995 19216 1996 19256
rect 2036 19216 2037 19256
rect 1995 19207 2037 19216
rect 4003 19256 4061 19257
rect 4003 19216 4012 19256
rect 4052 19216 4061 19256
rect 4003 19215 4061 19216
rect 4299 19256 4341 19265
rect 4299 19216 4300 19256
rect 4340 19216 4341 19256
rect 4299 19207 4341 19216
rect 4395 19256 4437 19265
rect 4395 19216 4396 19256
rect 4436 19216 4437 19256
rect 4395 19207 4437 19216
rect 835 19088 893 19089
rect 835 19048 844 19088
rect 884 19048 893 19088
rect 835 19047 893 19048
rect 2667 19088 2709 19097
rect 2667 19048 2668 19088
rect 2708 19048 2709 19088
rect 2667 19039 2709 19048
rect 3723 19088 3765 19097
rect 3723 19048 3724 19088
rect 3764 19048 3765 19088
rect 3723 19039 3765 19048
rect 576 18920 5952 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 5952 18920
rect 576 18856 5952 18880
rect 74016 18920 80736 18944
rect 74016 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80736 18920
rect 74016 18856 80736 18880
rect 835 18752 893 18753
rect 835 18712 844 18752
rect 884 18712 893 18752
rect 835 18711 893 18712
rect 3435 18668 3477 18677
rect 3435 18628 3436 18668
rect 3476 18628 3477 18668
rect 3435 18619 3477 18628
rect 3811 18584 3869 18585
rect 3811 18544 3820 18584
rect 3860 18544 3869 18584
rect 3811 18543 3869 18544
rect 4675 18584 4733 18585
rect 4675 18544 4684 18584
rect 4724 18544 4733 18584
rect 4675 18543 4733 18544
rect 1891 18500 1949 18501
rect 1891 18460 1900 18500
rect 1940 18460 1949 18500
rect 1891 18459 1949 18460
rect 2275 18500 2333 18501
rect 2275 18460 2284 18500
rect 2324 18460 2333 18500
rect 2275 18459 2333 18460
rect 5835 18500 5877 18509
rect 5835 18460 5836 18500
rect 5876 18460 5877 18500
rect 5835 18451 5877 18460
rect 2091 18416 2133 18425
rect 2091 18376 2092 18416
rect 2132 18376 2133 18416
rect 2091 18367 2133 18376
rect 2475 18332 2517 18341
rect 2475 18292 2476 18332
rect 2516 18292 2517 18332
rect 2475 18283 2517 18292
rect 576 18164 5952 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 5952 18164
rect 576 18100 5952 18124
rect 74016 18164 80736 18188
rect 74016 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 80736 18164
rect 74016 18100 80736 18124
rect 4491 17996 4533 18005
rect 4491 17956 4492 17996
rect 4532 17956 4533 17996
rect 4491 17947 4533 17956
rect 1507 17912 1565 17913
rect 1507 17872 1516 17912
rect 1556 17872 1565 17912
rect 1507 17871 1565 17872
rect 4099 17912 4157 17913
rect 4099 17872 4108 17912
rect 4148 17872 4157 17912
rect 4099 17871 4157 17872
rect 4291 17828 4349 17829
rect 4291 17788 4300 17828
rect 4340 17788 4349 17828
rect 4291 17787 4349 17788
rect 835 17744 893 17745
rect 835 17704 844 17744
rect 884 17704 893 17744
rect 835 17703 893 17704
rect 1131 17744 1173 17753
rect 1131 17704 1132 17744
rect 1172 17704 1173 17744
rect 1131 17695 1173 17704
rect 1227 17744 1269 17753
rect 1227 17704 1228 17744
rect 1268 17704 1269 17744
rect 1227 17695 1269 17704
rect 1707 17744 1749 17753
rect 1707 17704 1708 17744
rect 1748 17704 1749 17744
rect 1707 17695 1749 17704
rect 2083 17744 2141 17745
rect 2083 17704 2092 17744
rect 2132 17704 2141 17744
rect 2083 17703 2141 17704
rect 2947 17744 3005 17745
rect 2947 17704 2956 17744
rect 2996 17704 3005 17744
rect 2947 17703 3005 17704
rect 576 17408 5952 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 5952 17408
rect 576 17344 5952 17368
rect 74016 17408 80736 17432
rect 74016 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80736 17408
rect 74016 17344 80736 17368
rect 835 17240 893 17241
rect 835 17200 844 17240
rect 884 17200 893 17240
rect 835 17199 893 17200
rect 1219 17240 1277 17241
rect 1219 17200 1228 17240
rect 1268 17200 1277 17240
rect 1219 17199 1277 17200
rect 80611 17240 80669 17241
rect 80611 17200 80620 17240
rect 80660 17200 80669 17240
rect 80611 17199 80669 17200
rect 77739 17156 77781 17165
rect 77739 17116 77740 17156
rect 77780 17116 77781 17156
rect 77739 17107 77781 17116
rect 3435 17072 3477 17081
rect 3435 17032 3436 17072
rect 3476 17032 3477 17072
rect 3435 17023 3477 17032
rect 3811 17072 3869 17073
rect 3811 17032 3820 17072
rect 3860 17032 3869 17072
rect 3811 17031 3869 17032
rect 4675 17072 4733 17073
rect 4675 17032 4684 17072
rect 4724 17032 4733 17072
rect 4675 17031 4733 17032
rect 77347 17072 77405 17073
rect 77347 17032 77356 17072
rect 77396 17032 77405 17072
rect 77347 17031 77405 17032
rect 77643 17072 77685 17081
rect 77643 17032 77644 17072
rect 77684 17032 77685 17072
rect 77643 17023 77685 17032
rect 78219 17072 78261 17081
rect 78219 17032 78220 17072
rect 78260 17032 78261 17072
rect 78219 17023 78261 17032
rect 78595 17072 78653 17073
rect 78595 17032 78604 17072
rect 78644 17032 78653 17072
rect 78595 17031 78653 17032
rect 79459 17072 79517 17073
rect 79459 17032 79468 17072
rect 79508 17032 79517 17072
rect 79459 17031 79517 17032
rect 78019 16904 78077 16905
rect 78019 16864 78028 16904
rect 78068 16864 78077 16904
rect 78019 16863 78077 16864
rect 5827 16820 5885 16821
rect 5827 16780 5836 16820
rect 5876 16780 5885 16820
rect 5827 16779 5885 16780
rect 80611 16820 80669 16821
rect 80611 16780 80620 16820
rect 80660 16780 80669 16820
rect 80611 16779 80669 16780
rect 576 16652 5952 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 5952 16652
rect 576 16588 5952 16612
rect 74016 16652 80736 16676
rect 74016 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 80736 16652
rect 74016 16588 80736 16612
rect 4003 16484 4061 16485
rect 4003 16444 4012 16484
rect 4052 16444 4061 16484
rect 4003 16443 4061 16444
rect 4963 16484 5021 16485
rect 4963 16444 4972 16484
rect 5012 16444 5021 16484
rect 4963 16443 5021 16444
rect 1987 16232 2045 16233
rect 1987 16192 1996 16232
rect 2036 16192 2045 16232
rect 1987 16191 2045 16192
rect 2851 16232 2909 16233
rect 2851 16192 2860 16232
rect 2900 16192 2909 16232
rect 2851 16191 2909 16192
rect 4291 16232 4349 16233
rect 4291 16192 4300 16232
rect 4340 16192 4349 16232
rect 4291 16191 4349 16192
rect 4587 16232 4629 16241
rect 4587 16192 4588 16232
rect 4628 16192 4629 16232
rect 4587 16183 4629 16192
rect 4683 16232 4725 16241
rect 4683 16192 4684 16232
rect 4724 16192 4725 16232
rect 4683 16183 4725 16192
rect 1611 16148 1653 16157
rect 1611 16108 1612 16148
rect 1652 16108 1653 16148
rect 1611 16099 1653 16108
rect 835 16064 893 16065
rect 835 16024 844 16064
rect 884 16024 893 16064
rect 835 16023 893 16024
rect 4003 16064 4061 16065
rect 4003 16024 4012 16064
rect 4052 16024 4061 16064
rect 4003 16023 4061 16024
rect 576 15896 5952 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 5952 15896
rect 576 15832 5952 15856
rect 74016 15896 80736 15920
rect 74016 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80736 15896
rect 74016 15832 80736 15856
rect 5827 15728 5885 15729
rect 5827 15688 5836 15728
rect 5876 15688 5885 15728
rect 5827 15687 5885 15688
rect 1507 15560 1565 15561
rect 1507 15520 1516 15560
rect 1556 15520 1565 15560
rect 1507 15519 1565 15520
rect 1803 15560 1845 15569
rect 1803 15520 1804 15560
rect 1844 15520 1845 15560
rect 1803 15511 1845 15520
rect 1899 15560 1941 15569
rect 1899 15520 1900 15560
rect 1940 15520 1941 15560
rect 1899 15511 1941 15520
rect 3435 15560 3477 15569
rect 3435 15520 3436 15560
rect 3476 15520 3477 15560
rect 3435 15511 3477 15520
rect 3811 15560 3869 15561
rect 3811 15520 3820 15560
rect 3860 15520 3869 15560
rect 3811 15519 3869 15520
rect 4675 15560 4733 15561
rect 4675 15520 4684 15560
rect 4724 15520 4733 15560
rect 4675 15519 4733 15520
rect 643 15476 701 15477
rect 643 15436 652 15476
rect 692 15436 701 15476
rect 643 15435 701 15436
rect 2179 15392 2237 15393
rect 2179 15352 2188 15392
rect 2228 15352 2237 15392
rect 2179 15351 2237 15352
rect 843 15308 885 15317
rect 843 15268 844 15308
rect 884 15268 885 15308
rect 843 15259 885 15268
rect 576 15140 5952 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 5952 15140
rect 576 15076 5952 15100
rect 74016 15140 80736 15164
rect 74016 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 80736 15140
rect 74016 15076 80736 15100
rect 4963 14972 5021 14973
rect 4963 14932 4972 14972
rect 5012 14932 5021 14972
rect 4963 14931 5021 14932
rect 4003 14888 4061 14889
rect 4003 14848 4012 14888
rect 4052 14848 4061 14888
rect 4003 14847 4061 14848
rect 643 14804 701 14805
rect 643 14764 652 14804
rect 692 14764 701 14804
rect 643 14763 701 14764
rect 1987 14720 2045 14721
rect 1987 14680 1996 14720
rect 2036 14680 2045 14720
rect 1987 14679 2045 14680
rect 2851 14720 2909 14721
rect 2851 14680 2860 14720
rect 2900 14680 2909 14720
rect 2851 14679 2909 14680
rect 4291 14720 4349 14721
rect 4291 14680 4300 14720
rect 4340 14680 4349 14720
rect 4291 14679 4349 14680
rect 4587 14720 4629 14729
rect 4587 14680 4588 14720
rect 4628 14680 4629 14720
rect 4587 14671 4629 14680
rect 4683 14720 4725 14729
rect 4683 14680 4684 14720
rect 4724 14680 4725 14720
rect 4683 14671 4725 14680
rect 1611 14636 1653 14645
rect 1611 14596 1612 14636
rect 1652 14596 1653 14636
rect 1611 14587 1653 14596
rect 843 14552 885 14561
rect 843 14512 844 14552
rect 884 14512 885 14552
rect 843 14503 885 14512
rect 576 14384 5952 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 5952 14384
rect 576 14320 5952 14344
rect 74016 14384 80736 14408
rect 74016 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80736 14384
rect 74016 14320 80736 14344
rect 1507 14048 1565 14049
rect 1507 14008 1516 14048
rect 1556 14008 1565 14048
rect 1507 14007 1565 14008
rect 1803 14048 1845 14057
rect 1803 14008 1804 14048
rect 1844 14008 1845 14048
rect 1803 13999 1845 14008
rect 1899 14048 1941 14057
rect 1899 14008 1900 14048
rect 1940 14008 1941 14048
rect 1899 13999 1941 14008
rect 3619 14048 3677 14049
rect 3619 14008 3628 14048
rect 3668 14008 3677 14048
rect 3619 14007 3677 14008
rect 3915 14048 3957 14057
rect 3915 14008 3916 14048
rect 3956 14008 3957 14048
rect 3915 13999 3957 14008
rect 4011 14048 4053 14057
rect 4011 14008 4012 14048
rect 4052 14008 4053 14048
rect 4011 13999 4053 14008
rect 2179 13880 2237 13881
rect 2179 13840 2188 13880
rect 2228 13840 2237 13880
rect 2179 13839 2237 13840
rect 4291 13796 4349 13797
rect 4291 13756 4300 13796
rect 4340 13756 4349 13796
rect 4291 13755 4349 13756
rect 576 13628 5952 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 5952 13628
rect 576 13564 5952 13588
rect 74016 13628 80736 13652
rect 74016 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 80736 13628
rect 74016 13564 80736 13588
rect 5827 13460 5885 13461
rect 5827 13420 5836 13460
rect 5876 13420 5885 13460
rect 5827 13419 5885 13420
rect 1219 13208 1277 13209
rect 1219 13168 1228 13208
rect 1268 13168 1277 13208
rect 1219 13167 1277 13168
rect 2083 13208 2141 13209
rect 2083 13168 2092 13208
rect 2132 13168 2141 13208
rect 2083 13167 2141 13168
rect 3435 13208 3477 13217
rect 3435 13168 3436 13208
rect 3476 13168 3477 13208
rect 3435 13159 3477 13168
rect 3811 13208 3869 13209
rect 3811 13168 3820 13208
rect 3860 13168 3869 13208
rect 3811 13167 3869 13168
rect 4675 13208 4733 13209
rect 4675 13168 4684 13208
rect 4724 13168 4733 13208
rect 4675 13167 4733 13168
rect 843 13124 885 13133
rect 843 13084 844 13124
rect 884 13084 885 13124
rect 843 13075 885 13084
rect 3235 13040 3293 13041
rect 3235 13000 3244 13040
rect 3284 13000 3293 13040
rect 3235 12999 3293 13000
rect 5827 13040 5885 13041
rect 5827 13000 5836 13040
rect 5876 13000 5885 13040
rect 5827 12999 5885 13000
rect 576 12872 5952 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 5952 12872
rect 576 12808 5952 12832
rect 74016 12872 80736 12896
rect 74016 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80736 12872
rect 74016 12808 80736 12832
rect 2187 12746 2229 12755
rect 843 12704 885 12713
rect 843 12664 844 12704
rect 884 12664 885 12704
rect 2187 12706 2188 12746
rect 2228 12706 2229 12746
rect 2187 12697 2229 12706
rect 843 12655 885 12664
rect 1507 12536 1565 12537
rect 1507 12496 1516 12536
rect 1556 12496 1565 12536
rect 1507 12495 1565 12496
rect 1803 12536 1845 12545
rect 1803 12496 1804 12536
rect 1844 12496 1845 12536
rect 1803 12487 1845 12496
rect 1899 12536 1941 12545
rect 1899 12496 1900 12536
rect 1940 12496 1941 12536
rect 1899 12487 1941 12496
rect 3435 12536 3477 12545
rect 3435 12496 3436 12536
rect 3476 12496 3477 12536
rect 3435 12487 3477 12496
rect 3811 12536 3869 12537
rect 3811 12496 3820 12536
rect 3860 12496 3869 12536
rect 3811 12495 3869 12496
rect 4675 12536 4733 12537
rect 4675 12496 4684 12536
rect 4724 12496 4733 12536
rect 4675 12495 4733 12496
rect 643 12452 701 12453
rect 643 12412 652 12452
rect 692 12412 701 12452
rect 643 12411 701 12412
rect 1027 12452 1085 12453
rect 1027 12412 1036 12452
rect 1076 12412 1085 12452
rect 1027 12411 1085 12412
rect 1227 12368 1269 12377
rect 1227 12328 1228 12368
rect 1268 12328 1269 12368
rect 1227 12319 1269 12328
rect 5827 12284 5885 12285
rect 5827 12244 5836 12284
rect 5876 12244 5885 12284
rect 5827 12243 5885 12244
rect 576 12116 5952 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 5952 12116
rect 576 12052 5952 12076
rect 74016 12116 80736 12140
rect 74016 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 80736 12116
rect 74016 12052 80736 12076
rect 4579 11948 4637 11949
rect 4579 11908 4588 11948
rect 4628 11908 4637 11948
rect 4579 11907 4637 11908
rect 643 11780 701 11781
rect 643 11740 652 11780
rect 692 11740 701 11780
rect 643 11739 701 11740
rect 3907 11696 3965 11697
rect 3907 11656 3916 11696
rect 3956 11656 3965 11696
rect 3907 11655 3965 11656
rect 4203 11696 4245 11705
rect 4203 11656 4204 11696
rect 4244 11656 4245 11696
rect 4203 11647 4245 11656
rect 4299 11696 4341 11705
rect 4299 11656 4300 11696
rect 4340 11656 4341 11696
rect 4299 11647 4341 11656
rect 843 11528 885 11537
rect 843 11488 844 11528
rect 884 11488 885 11528
rect 843 11479 885 11488
rect 576 11360 5952 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 5952 11360
rect 576 11296 5952 11320
rect 74016 11360 80736 11384
rect 74016 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80736 11360
rect 74016 11296 80736 11320
rect 2379 11234 2421 11243
rect 2379 11194 2380 11234
rect 2420 11194 2421 11234
rect 2379 11185 2421 11194
rect 4963 11192 5021 11193
rect 4963 11152 4972 11192
rect 5012 11152 5021 11192
rect 4963 11151 5021 11152
rect 2091 11108 2133 11117
rect 2091 11068 2092 11108
rect 2132 11068 2133 11108
rect 2091 11059 2133 11068
rect 2571 11108 2613 11117
rect 2571 11068 2572 11108
rect 2612 11068 2613 11108
rect 2571 11059 2613 11068
rect 1699 11024 1757 11025
rect 1699 10984 1708 11024
rect 1748 10984 1757 11024
rect 1699 10983 1757 10984
rect 1995 11024 2037 11033
rect 1995 10984 1996 11024
rect 2036 10984 2037 11024
rect 1995 10975 2037 10984
rect 2947 11024 3005 11025
rect 2947 10984 2956 11024
rect 2996 10984 3005 11024
rect 2947 10983 3005 10984
rect 3811 11024 3869 11025
rect 3811 10984 3820 11024
rect 3860 10984 3869 11024
rect 3811 10983 3869 10984
rect 643 10940 701 10941
rect 643 10900 652 10940
rect 692 10900 701 10940
rect 643 10899 701 10900
rect 843 10772 885 10781
rect 843 10732 844 10772
rect 884 10732 885 10772
rect 843 10723 885 10732
rect 576 10604 5952 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 5952 10604
rect 576 10540 5952 10564
rect 74016 10604 80736 10628
rect 74016 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 80736 10604
rect 74016 10540 80736 10564
rect 643 10268 701 10269
rect 643 10228 652 10268
rect 692 10228 701 10268
rect 643 10227 701 10228
rect 5835 10268 5877 10277
rect 5835 10228 5836 10268
rect 5876 10228 5877 10268
rect 5835 10219 5877 10228
rect 3811 10184 3869 10185
rect 3811 10144 3820 10184
rect 3860 10144 3869 10184
rect 3811 10143 3869 10144
rect 4675 10184 4733 10185
rect 4675 10144 4684 10184
rect 4724 10144 4733 10184
rect 4675 10143 4733 10144
rect 3435 10100 3477 10109
rect 3435 10060 3436 10100
rect 3476 10060 3477 10100
rect 3435 10051 3477 10060
rect 843 10016 885 10025
rect 843 9976 844 10016
rect 884 9976 885 10016
rect 843 9967 885 9976
rect 576 9848 5952 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 5952 9848
rect 576 9784 5952 9808
rect 74016 9848 80736 9872
rect 74016 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80736 9848
rect 74016 9784 80736 9808
rect 4003 9512 4061 9513
rect 4003 9472 4012 9512
rect 4052 9472 4061 9512
rect 4003 9471 4061 9472
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4299 9463 4341 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 643 9428 701 9429
rect 643 9388 652 9428
rect 692 9388 701 9428
rect 643 9387 701 9388
rect 4675 9344 4733 9345
rect 4675 9304 4684 9344
rect 4724 9304 4733 9344
rect 4675 9303 4733 9304
rect 843 9260 885 9269
rect 843 9220 844 9260
rect 884 9220 885 9260
rect 843 9211 885 9220
rect 576 9092 5952 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 5952 9092
rect 576 9028 5952 9052
rect 74016 9092 80736 9116
rect 74016 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 80736 9092
rect 74016 9028 80736 9052
rect 835 8504 893 8505
rect 835 8464 844 8504
rect 884 8464 893 8504
rect 835 8463 893 8464
rect 576 8336 5952 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 5952 8336
rect 576 8272 5952 8296
rect 74016 8336 80736 8360
rect 74016 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80736 8336
rect 74016 8272 80736 8296
rect 835 8168 893 8169
rect 835 8128 844 8168
rect 884 8128 893 8168
rect 835 8127 893 8128
rect 5827 8168 5885 8169
rect 5827 8128 5836 8168
rect 5876 8128 5885 8168
rect 5827 8127 5885 8128
rect 3435 8000 3477 8009
rect 3435 7960 3436 8000
rect 3476 7960 3477 8000
rect 3435 7951 3477 7960
rect 3811 8000 3869 8001
rect 3811 7960 3820 8000
rect 3860 7960 3869 8000
rect 3811 7959 3869 7960
rect 4675 8000 4733 8001
rect 4675 7960 4684 8000
rect 4724 7960 4733 8000
rect 4675 7959 4733 7960
rect 576 7580 5952 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 5952 7580
rect 576 7516 5952 7540
rect 74016 7580 80736 7604
rect 74016 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 80736 7580
rect 74016 7516 80736 7540
rect 5059 7412 5117 7413
rect 5059 7372 5068 7412
rect 5108 7372 5117 7412
rect 5059 7371 5117 7372
rect 4387 7160 4445 7161
rect 4387 7120 4396 7160
rect 4436 7120 4445 7160
rect 4387 7119 4445 7120
rect 4683 7160 4725 7169
rect 4683 7120 4684 7160
rect 4724 7120 4725 7160
rect 4683 7111 4725 7120
rect 4779 7160 4821 7169
rect 4779 7120 4780 7160
rect 4820 7120 4821 7160
rect 4779 7111 4821 7120
rect 835 6992 893 6993
rect 835 6952 844 6992
rect 884 6952 893 6992
rect 835 6951 893 6952
rect 576 6824 5952 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 5952 6824
rect 576 6760 5952 6784
rect 74016 6824 80736 6848
rect 74016 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80736 6824
rect 74016 6760 80736 6784
rect 80227 6488 80285 6489
rect 80227 6448 80236 6488
rect 80276 6448 80285 6488
rect 80227 6447 80285 6448
rect 78883 6404 78941 6405
rect 78883 6364 78892 6404
rect 78932 6364 78941 6404
rect 78883 6363 78941 6364
rect 576 6068 5952 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 5952 6068
rect 576 6004 5952 6028
rect 74016 6068 80736 6092
rect 74016 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 80736 6068
rect 74016 6004 80736 6028
rect 835 5480 893 5481
rect 835 5440 844 5480
rect 884 5440 893 5480
rect 835 5439 893 5440
rect 576 5312 80736 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80736 5312
rect 576 5248 80736 5272
rect 835 5144 893 5145
rect 835 5104 844 5144
rect 884 5104 893 5144
rect 835 5103 893 5104
rect 18403 5144 18461 5145
rect 18403 5104 18412 5144
rect 18452 5104 18461 5144
rect 18403 5103 18461 5104
rect 31947 5144 31989 5153
rect 31947 5104 31948 5144
rect 31988 5104 31989 5144
rect 31947 5095 31989 5104
rect 32131 5144 32189 5145
rect 32131 5104 32140 5144
rect 32180 5104 32189 5144
rect 32131 5103 32189 5104
rect 32715 5144 32757 5153
rect 32715 5104 32716 5144
rect 32756 5104 32757 5144
rect 32715 5095 32757 5104
rect 21771 5060 21813 5069
rect 21771 5020 21772 5060
rect 21812 5020 21813 5060
rect 21771 5011 21813 5020
rect 26091 5060 26133 5069
rect 26091 5020 26092 5060
rect 26132 5020 26133 5060
rect 26091 5011 26133 5020
rect 39243 5060 39285 5069
rect 39243 5020 39244 5060
rect 39284 5020 39285 5060
rect 39243 5011 39285 5020
rect 16011 4976 16053 4985
rect 16011 4936 16012 4976
rect 16052 4936 16053 4976
rect 16011 4927 16053 4936
rect 16387 4976 16445 4977
rect 16387 4936 16396 4976
rect 16436 4936 16445 4976
rect 21379 4976 21437 4977
rect 16387 4935 16445 4936
rect 17251 4965 17309 4966
rect 17251 4925 17260 4965
rect 17300 4925 17309 4965
rect 21379 4936 21388 4976
rect 21428 4936 21437 4976
rect 21379 4935 21437 4936
rect 21675 4976 21717 4985
rect 21675 4936 21676 4976
rect 21716 4936 21717 4976
rect 21675 4927 21717 4936
rect 24067 4976 24125 4977
rect 24067 4936 24076 4976
rect 24116 4936 24125 4976
rect 24067 4935 24125 4936
rect 24363 4976 24405 4985
rect 24363 4936 24364 4976
rect 24404 4936 24405 4976
rect 24363 4927 24405 4936
rect 24459 4976 24501 4985
rect 24459 4936 24460 4976
rect 24500 4936 24501 4976
rect 24459 4927 24501 4936
rect 25699 4976 25757 4977
rect 25699 4936 25708 4976
rect 25748 4936 25757 4976
rect 25699 4935 25757 4936
rect 25995 4976 26037 4985
rect 25995 4936 25996 4976
rect 26036 4936 26037 4976
rect 25995 4927 26037 4936
rect 30307 4976 30365 4977
rect 30307 4936 30316 4976
rect 30356 4936 30365 4976
rect 30307 4935 30365 4936
rect 30603 4976 30645 4985
rect 30603 4936 30604 4976
rect 30644 4936 30645 4976
rect 30603 4927 30645 4936
rect 30699 4976 30741 4985
rect 30699 4936 30700 4976
rect 30740 4936 30741 4976
rect 30699 4927 30741 4936
rect 32227 4976 32285 4977
rect 32227 4936 32236 4976
rect 32276 4936 32285 4976
rect 32227 4935 32285 4936
rect 36939 4976 36981 4985
rect 36939 4936 36940 4976
rect 36980 4936 36981 4976
rect 36939 4927 36981 4936
rect 37123 4976 37181 4977
rect 37123 4936 37132 4976
rect 37172 4936 37181 4976
rect 37123 4935 37181 4936
rect 38571 4976 38613 4985
rect 38571 4936 38572 4976
rect 38612 4936 38613 4976
rect 38571 4927 38613 4936
rect 38947 4976 39005 4977
rect 38947 4936 38956 4976
rect 38996 4936 39005 4976
rect 38947 4935 39005 4936
rect 39147 4976 39189 4985
rect 39147 4936 39148 4976
rect 39188 4936 39189 4976
rect 39147 4927 39189 4936
rect 39331 4976 39389 4977
rect 39331 4936 39340 4976
rect 39380 4936 39389 4976
rect 39331 4935 39389 4936
rect 45187 4976 45245 4977
rect 45187 4936 45196 4976
rect 45236 4936 45245 4976
rect 45187 4935 45245 4936
rect 51715 4976 51773 4977
rect 51715 4936 51724 4976
rect 51764 4936 51773 4976
rect 51715 4935 51773 4936
rect 52011 4976 52053 4985
rect 52011 4936 52012 4976
rect 52052 4936 52053 4976
rect 52011 4927 52053 4936
rect 52107 4976 52149 4985
rect 52107 4936 52108 4976
rect 52148 4936 52149 4976
rect 52107 4927 52149 4936
rect 17251 4924 17309 4925
rect 25219 4892 25277 4893
rect 25219 4852 25228 4892
rect 25268 4852 25277 4892
rect 25219 4851 25277 4852
rect 26563 4892 26621 4893
rect 26563 4852 26572 4892
rect 26612 4852 26621 4892
rect 26563 4851 26621 4852
rect 26947 4892 27005 4893
rect 26947 4852 26956 4892
rect 26996 4852 27005 4892
rect 26947 4851 27005 4852
rect 38667 4892 38709 4901
rect 38667 4852 38668 4892
rect 38708 4852 38709 4892
rect 38667 4843 38709 4852
rect 38859 4892 38901 4901
rect 38859 4852 38860 4892
rect 38900 4852 38901 4892
rect 38859 4843 38901 4852
rect 43843 4892 43901 4893
rect 43843 4852 43852 4892
rect 43892 4852 43901 4892
rect 43843 4851 43901 4852
rect 46819 4892 46877 4893
rect 46819 4852 46828 4892
rect 46868 4852 46877 4892
rect 46819 4851 46877 4852
rect 25419 4808 25461 4817
rect 25419 4768 25420 4808
rect 25460 4768 25461 4808
rect 25419 4759 25461 4768
rect 32419 4808 32477 4809
rect 32419 4768 32428 4808
rect 32468 4768 32477 4808
rect 32419 4767 32477 4768
rect 38763 4808 38805 4817
rect 38763 4768 38764 4808
rect 38804 4768 38805 4808
rect 38763 4759 38805 4768
rect 22051 4724 22109 4725
rect 22051 4684 22060 4724
rect 22100 4684 22109 4724
rect 22051 4683 22109 4684
rect 24739 4724 24797 4725
rect 24739 4684 24748 4724
rect 24788 4684 24797 4724
rect 24739 4683 24797 4684
rect 26371 4724 26429 4725
rect 26371 4684 26380 4724
rect 26420 4684 26429 4724
rect 26371 4683 26429 4684
rect 26763 4724 26805 4733
rect 26763 4684 26764 4724
rect 26804 4684 26805 4724
rect 26763 4675 26805 4684
rect 27147 4724 27189 4733
rect 27147 4684 27148 4724
rect 27188 4684 27189 4724
rect 27147 4675 27189 4684
rect 30979 4724 31037 4725
rect 30979 4684 30988 4724
rect 31028 4684 31037 4724
rect 30979 4683 31037 4684
rect 37035 4724 37077 4733
rect 37035 4684 37036 4724
rect 37076 4684 37077 4724
rect 37035 4675 37077 4684
rect 47019 4724 47061 4733
rect 47019 4684 47020 4724
rect 47060 4684 47061 4724
rect 47019 4675 47061 4684
rect 52387 4724 52445 4725
rect 52387 4684 52396 4724
rect 52436 4684 52445 4724
rect 52387 4683 52445 4684
rect 576 4556 80736 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 80736 4556
rect 576 4492 80736 4516
rect 17251 4388 17309 4389
rect 17251 4348 17260 4388
rect 17300 4348 17309 4388
rect 17251 4347 17309 4348
rect 22435 4388 22493 4389
rect 22435 4348 22444 4388
rect 22484 4348 22493 4388
rect 22435 4347 22493 4348
rect 19843 4304 19901 4305
rect 19843 4264 19852 4304
rect 19892 4264 19901 4304
rect 19843 4263 19901 4264
rect 27043 4304 27101 4305
rect 27043 4264 27052 4304
rect 27092 4264 27101 4304
rect 27043 4263 27101 4264
rect 30883 4304 30941 4305
rect 30883 4264 30892 4304
rect 30932 4264 30941 4304
rect 30883 4263 30941 4264
rect 36363 4304 36405 4313
rect 36363 4264 36364 4304
rect 36404 4264 36405 4304
rect 36363 4255 36405 4264
rect 38667 4304 38709 4313
rect 38667 4264 38668 4304
rect 38708 4264 38709 4304
rect 38667 4255 38709 4264
rect 41259 4304 41301 4313
rect 41259 4264 41260 4304
rect 41300 4264 41301 4304
rect 41259 4255 41301 4264
rect 46531 4304 46589 4305
rect 46531 4264 46540 4304
rect 46580 4264 46589 4304
rect 46531 4263 46589 4264
rect 47779 4304 47837 4305
rect 47779 4264 47788 4304
rect 47828 4264 47837 4304
rect 47779 4263 47837 4264
rect 54019 4304 54077 4305
rect 54019 4264 54028 4304
rect 54068 4264 54077 4304
rect 54019 4263 54077 4264
rect 50379 4220 50421 4229
rect 50379 4180 50380 4220
rect 50420 4180 50421 4220
rect 47491 4178 47549 4179
rect 16579 4136 16637 4137
rect 16579 4096 16588 4136
rect 16628 4096 16637 4136
rect 16579 4095 16637 4096
rect 16875 4136 16917 4145
rect 16875 4096 16876 4136
rect 16916 4096 16917 4136
rect 16875 4087 16917 4096
rect 16971 4136 17013 4145
rect 16971 4096 16972 4136
rect 17012 4096 17013 4136
rect 16971 4087 17013 4096
rect 17827 4136 17885 4137
rect 17827 4096 17836 4136
rect 17876 4096 17885 4136
rect 17827 4095 17885 4096
rect 18691 4136 18749 4137
rect 18691 4096 18700 4136
rect 18740 4096 18749 4136
rect 18691 4095 18749 4096
rect 20419 4136 20477 4137
rect 20419 4096 20428 4136
rect 20468 4096 20477 4136
rect 20419 4095 20477 4096
rect 21283 4136 21341 4137
rect 21283 4096 21292 4136
rect 21332 4096 21341 4136
rect 21283 4095 21341 4096
rect 23403 4136 23445 4145
rect 23403 4096 23404 4136
rect 23444 4096 23445 4136
rect 23403 4087 23445 4096
rect 23779 4136 23837 4137
rect 23779 4096 23788 4136
rect 23828 4096 23837 4136
rect 23779 4095 23837 4096
rect 24643 4136 24701 4137
rect 24643 4096 24652 4136
rect 24692 4096 24701 4136
rect 24643 4095 24701 4096
rect 26371 4136 26429 4137
rect 26371 4096 26380 4136
rect 26420 4096 26429 4136
rect 26371 4095 26429 4096
rect 26667 4136 26709 4145
rect 26667 4096 26668 4136
rect 26708 4096 26709 4136
rect 26667 4087 26709 4096
rect 26763 4136 26805 4145
rect 26763 4096 26764 4136
rect 26804 4096 26805 4136
rect 26763 4087 26805 4096
rect 27243 4136 27285 4145
rect 27243 4096 27244 4136
rect 27284 4096 27285 4136
rect 27243 4087 27285 4096
rect 27619 4136 27677 4137
rect 27619 4096 27628 4136
rect 27668 4096 27677 4136
rect 27619 4095 27677 4096
rect 28483 4136 28541 4137
rect 28483 4096 28492 4136
rect 28532 4096 28541 4136
rect 28483 4095 28541 4096
rect 30211 4136 30269 4137
rect 30211 4096 30220 4136
rect 30260 4096 30269 4136
rect 30211 4095 30269 4096
rect 30507 4136 30549 4145
rect 30507 4096 30508 4136
rect 30548 4096 30549 4136
rect 30507 4087 30549 4096
rect 31083 4136 31125 4145
rect 31083 4096 31084 4136
rect 31124 4096 31125 4136
rect 31083 4087 31125 4096
rect 31459 4136 31517 4137
rect 31459 4096 31468 4136
rect 31508 4096 31517 4136
rect 31459 4095 31517 4096
rect 32323 4136 32381 4137
rect 32323 4096 32332 4136
rect 32372 4096 32381 4136
rect 32323 4095 32381 4096
rect 34723 4136 34781 4137
rect 34723 4096 34732 4136
rect 34772 4096 34781 4136
rect 34723 4095 34781 4096
rect 35115 4136 35157 4145
rect 35115 4096 35116 4136
rect 35156 4096 35157 4136
rect 35115 4087 35157 4096
rect 35307 4136 35349 4145
rect 35307 4096 35308 4136
rect 35348 4096 35349 4136
rect 35307 4087 35349 4096
rect 36267 4136 36309 4145
rect 36267 4096 36268 4136
rect 36308 4096 36309 4136
rect 36267 4087 36309 4096
rect 36451 4136 36509 4137
rect 36451 4096 36460 4136
rect 36500 4096 36509 4136
rect 36451 4095 36509 4096
rect 40011 4136 40053 4145
rect 40011 4096 40012 4136
rect 40052 4096 40053 4136
rect 40011 4087 40053 4096
rect 40107 4136 40149 4145
rect 40107 4096 40108 4136
rect 40148 4096 40149 4136
rect 40107 4087 40149 4096
rect 40683 4136 40725 4145
rect 40683 4096 40684 4136
rect 40724 4096 40725 4136
rect 40683 4087 40725 4096
rect 40779 4136 40821 4145
rect 40779 4096 40780 4136
rect 40820 4096 40821 4136
rect 40779 4087 40821 4096
rect 40875 4136 40917 4145
rect 40875 4096 40876 4136
rect 40916 4096 40917 4136
rect 40875 4087 40917 4096
rect 40971 4136 41013 4145
rect 40971 4096 40972 4136
rect 41012 4096 41013 4136
rect 40971 4087 41013 4096
rect 42315 4136 42357 4145
rect 42315 4096 42316 4136
rect 42356 4096 42357 4136
rect 42315 4087 42357 4096
rect 42507 4136 42549 4145
rect 42507 4096 42508 4136
rect 42548 4096 42549 4136
rect 42507 4087 42549 4096
rect 42795 4136 42837 4145
rect 42795 4096 42796 4136
rect 42836 4096 42837 4136
rect 42795 4087 42837 4096
rect 42891 4136 42933 4145
rect 42891 4096 42892 4136
rect 42932 4096 42933 4136
rect 42891 4087 42933 4096
rect 43275 4136 43317 4145
rect 43275 4096 43276 4136
rect 43316 4096 43317 4136
rect 43275 4087 43317 4096
rect 43371 4136 43413 4145
rect 44331 4141 44373 4150
rect 43371 4096 43372 4136
rect 43412 4096 43413 4136
rect 43371 4087 43413 4096
rect 43843 4136 43901 4137
rect 43843 4096 43852 4136
rect 43892 4096 43901 4136
rect 43843 4095 43901 4096
rect 44331 4101 44332 4141
rect 44372 4101 44373 4141
rect 44331 4092 44373 4101
rect 45859 4136 45917 4137
rect 45859 4096 45868 4136
rect 45908 4096 45917 4136
rect 45859 4095 45917 4096
rect 46155 4136 46197 4145
rect 46155 4096 46156 4136
rect 46196 4096 46197 4136
rect 46155 4087 46197 4096
rect 47107 4136 47165 4137
rect 47107 4096 47116 4136
rect 47156 4096 47165 4136
rect 47107 4095 47165 4096
rect 47403 4136 47445 4145
rect 47491 4138 47500 4178
rect 47540 4138 47549 4178
rect 50379 4171 50421 4180
rect 47491 4137 47549 4138
rect 47403 4096 47404 4136
rect 47444 4096 47445 4136
rect 47403 4087 47445 4096
rect 47979 4136 48021 4145
rect 47979 4096 47980 4136
rect 48020 4096 48021 4136
rect 47979 4087 48021 4096
rect 48355 4136 48413 4137
rect 48355 4096 48364 4136
rect 48404 4096 48413 4136
rect 48355 4095 48413 4096
rect 49219 4136 49277 4137
rect 49219 4096 49228 4136
rect 49268 4096 49277 4136
rect 49219 4095 49277 4096
rect 50947 4136 51005 4137
rect 50947 4096 50956 4136
rect 50996 4096 51005 4136
rect 50947 4095 51005 4096
rect 51811 4136 51869 4137
rect 51811 4096 51820 4136
rect 51860 4096 51869 4136
rect 51811 4095 51869 4096
rect 53347 4136 53405 4137
rect 53347 4096 53356 4136
rect 53396 4096 53405 4136
rect 53347 4095 53405 4096
rect 53643 4136 53685 4145
rect 53643 4096 53644 4136
rect 53684 4096 53685 4136
rect 53643 4087 53685 4096
rect 54219 4136 54261 4145
rect 54219 4096 54220 4136
rect 54260 4096 54261 4136
rect 54219 4087 54261 4096
rect 54595 4136 54653 4137
rect 54595 4096 54604 4136
rect 54644 4096 54653 4136
rect 54595 4095 54653 4096
rect 55459 4136 55517 4137
rect 55459 4096 55468 4136
rect 55508 4096 55517 4136
rect 55459 4095 55517 4096
rect 17451 4052 17493 4061
rect 17451 4012 17452 4052
rect 17492 4012 17493 4052
rect 17451 4003 17493 4012
rect 20043 4052 20085 4061
rect 20043 4012 20044 4052
rect 20084 4012 20085 4052
rect 20043 4003 20085 4012
rect 30603 4052 30645 4061
rect 30603 4012 30604 4052
rect 30644 4012 30645 4052
rect 30603 4003 30645 4012
rect 46251 4052 46293 4061
rect 46251 4012 46252 4052
rect 46292 4012 46293 4052
rect 46251 4003 46293 4012
rect 50571 4052 50613 4061
rect 50571 4012 50572 4052
rect 50612 4012 50613 4052
rect 50571 4003 50613 4012
rect 53739 4052 53781 4061
rect 53739 4012 53740 4052
rect 53780 4012 53781 4052
rect 53739 4003 53781 4012
rect 835 3968 893 3969
rect 835 3928 844 3968
rect 884 3928 893 3968
rect 835 3927 893 3928
rect 25795 3968 25853 3969
rect 25795 3928 25804 3968
rect 25844 3928 25853 3968
rect 25795 3927 25853 3928
rect 29635 3968 29693 3969
rect 29635 3928 29644 3968
rect 29684 3928 29693 3968
rect 29635 3927 29693 3928
rect 33475 3968 33533 3969
rect 33475 3928 33484 3968
rect 33524 3928 33533 3968
rect 33475 3927 33533 3928
rect 34627 3968 34685 3969
rect 34627 3928 34636 3968
rect 34676 3928 34685 3968
rect 34627 3927 34685 3928
rect 34915 3968 34973 3969
rect 34915 3928 34924 3968
rect 34964 3928 34973 3968
rect 34915 3927 34973 3928
rect 35211 3968 35253 3977
rect 35211 3928 35212 3968
rect 35252 3928 35253 3968
rect 35211 3919 35253 3928
rect 40291 3968 40349 3969
rect 40291 3928 40300 3968
rect 40340 3928 40349 3968
rect 40291 3927 40349 3928
rect 42411 3968 42453 3977
rect 42411 3928 42412 3968
rect 42452 3928 42453 3968
rect 42411 3919 42453 3928
rect 44523 3968 44565 3977
rect 44523 3928 44524 3968
rect 44564 3928 44565 3968
rect 44523 3919 44565 3928
rect 52963 3968 53021 3969
rect 52963 3928 52972 3968
rect 53012 3928 53021 3968
rect 52963 3927 53021 3928
rect 56611 3968 56669 3969
rect 56611 3928 56620 3968
rect 56660 3928 56669 3968
rect 56611 3927 56669 3928
rect 576 3800 80736 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80736 3800
rect 576 3736 80736 3760
rect 835 3632 893 3633
rect 835 3592 844 3632
rect 884 3592 893 3632
rect 835 3591 893 3592
rect 23971 3632 24029 3633
rect 23971 3592 23980 3632
rect 24020 3592 24029 3632
rect 23971 3591 24029 3592
rect 28579 3632 28637 3633
rect 28579 3592 28588 3632
rect 28628 3592 28637 3632
rect 28579 3591 28637 3592
rect 31939 3632 31997 3633
rect 31939 3592 31948 3632
rect 31988 3592 31997 3632
rect 31939 3591 31997 3592
rect 32427 3632 32469 3641
rect 32427 3592 32428 3632
rect 32468 3592 32469 3632
rect 32427 3583 32469 3592
rect 41251 3632 41309 3633
rect 41251 3592 41260 3632
rect 41300 3592 41309 3632
rect 41251 3591 41309 3592
rect 48643 3632 48701 3633
rect 48643 3592 48652 3632
rect 48692 3592 48701 3632
rect 48643 3591 48701 3592
rect 54691 3632 54749 3633
rect 54691 3592 54700 3632
rect 54740 3592 54749 3632
rect 54691 3591 54749 3592
rect 17355 3548 17397 3557
rect 17355 3508 17356 3548
rect 17396 3508 17397 3548
rect 17259 3491 17301 3500
rect 17355 3499 17397 3508
rect 20619 3548 20661 3557
rect 20619 3508 20620 3548
rect 20660 3508 20661 3548
rect 20619 3499 20661 3508
rect 21579 3548 21621 3557
rect 21579 3508 21580 3548
rect 21620 3508 21621 3548
rect 21579 3499 21621 3508
rect 26187 3548 26229 3557
rect 26187 3508 26188 3548
rect 26228 3508 26229 3548
rect 26187 3499 26229 3508
rect 29547 3548 29589 3557
rect 29547 3508 29548 3548
rect 29588 3508 29589 3548
rect 29547 3499 29589 3508
rect 43083 3548 43125 3557
rect 43083 3508 43084 3548
rect 43124 3508 43125 3548
rect 43083 3499 43125 3508
rect 45387 3548 45429 3557
rect 45387 3508 45388 3548
rect 45428 3508 45429 3548
rect 45387 3499 45429 3508
rect 46251 3548 46293 3557
rect 46251 3508 46252 3548
rect 46292 3508 46293 3548
rect 46251 3499 46293 3508
rect 52299 3548 52341 3557
rect 52299 3508 52300 3548
rect 52340 3508 52341 3548
rect 52299 3499 52341 3508
rect 16963 3464 17021 3465
rect 16963 3424 16972 3464
rect 17012 3424 17021 3464
rect 17259 3451 17260 3491
rect 17300 3451 17301 3491
rect 17259 3442 17301 3451
rect 20227 3464 20285 3465
rect 16963 3423 17021 3424
rect 20227 3424 20236 3464
rect 20276 3424 20285 3464
rect 20227 3423 20285 3424
rect 20523 3464 20565 3473
rect 20523 3424 20524 3464
rect 20564 3424 20565 3464
rect 20523 3415 20565 3424
rect 21955 3464 22013 3465
rect 21955 3424 21964 3464
rect 22004 3424 22013 3464
rect 21955 3423 22013 3424
rect 22819 3464 22877 3465
rect 22819 3424 22828 3464
rect 22868 3424 22877 3464
rect 22819 3423 22877 3424
rect 26563 3464 26621 3465
rect 26563 3424 26572 3464
rect 26612 3424 26621 3464
rect 26563 3423 26621 3424
rect 27427 3464 27485 3465
rect 27427 3424 27436 3464
rect 27476 3424 27485 3464
rect 27427 3423 27485 3424
rect 29923 3464 29981 3465
rect 29923 3424 29932 3464
rect 29972 3424 29981 3464
rect 29923 3423 29981 3424
rect 30787 3464 30845 3465
rect 30787 3424 30796 3464
rect 30836 3424 30845 3464
rect 30787 3423 30845 3424
rect 32235 3464 32277 3473
rect 32235 3424 32236 3464
rect 32276 3424 32277 3464
rect 32235 3415 32277 3424
rect 32523 3464 32565 3473
rect 32523 3424 32524 3464
rect 32564 3424 32565 3464
rect 32523 3415 32565 3424
rect 34819 3464 34877 3465
rect 34819 3424 34828 3464
rect 34868 3424 34877 3464
rect 34819 3423 34877 3424
rect 35211 3464 35253 3473
rect 35211 3424 35212 3464
rect 35252 3424 35253 3464
rect 35211 3415 35253 3424
rect 36931 3464 36989 3465
rect 36931 3424 36940 3464
rect 36980 3424 36989 3464
rect 36931 3423 36989 3424
rect 37323 3464 37365 3473
rect 37323 3424 37324 3464
rect 37364 3424 37365 3464
rect 37323 3415 37365 3424
rect 38275 3464 38333 3465
rect 38275 3424 38284 3464
rect 38324 3424 38333 3464
rect 38275 3423 38333 3424
rect 38667 3464 38709 3473
rect 38667 3424 38668 3464
rect 38708 3424 38709 3464
rect 38667 3415 38709 3424
rect 40971 3464 41013 3473
rect 40971 3424 40972 3464
rect 41012 3424 41013 3464
rect 40971 3415 41013 3424
rect 41067 3464 41109 3473
rect 41067 3424 41068 3464
rect 41108 3424 41109 3464
rect 41067 3415 41109 3424
rect 41163 3464 41205 3473
rect 41163 3424 41164 3464
rect 41204 3424 41205 3464
rect 41163 3415 41205 3424
rect 42987 3464 43029 3473
rect 42987 3424 42988 3464
rect 43028 3424 43029 3464
rect 43267 3464 43325 3465
rect 42987 3415 43029 3424
rect 43171 3450 43229 3451
rect 43171 3410 43180 3450
rect 43220 3410 43229 3450
rect 43267 3424 43276 3464
rect 43316 3424 43325 3464
rect 43267 3423 43325 3424
rect 43939 3464 43997 3465
rect 43939 3424 43948 3464
rect 43988 3424 43997 3464
rect 43939 3423 43997 3424
rect 45187 3464 45245 3465
rect 45187 3424 45196 3464
rect 45236 3424 45245 3464
rect 45187 3423 45245 3424
rect 46627 3464 46685 3465
rect 46627 3424 46636 3464
rect 46676 3424 46685 3464
rect 49795 3464 49853 3465
rect 46627 3423 46685 3424
rect 47491 3453 47549 3454
rect 47491 3413 47500 3453
rect 47540 3413 47549 3453
rect 49795 3424 49804 3464
rect 49844 3424 49853 3464
rect 49795 3423 49853 3424
rect 50091 3464 50133 3473
rect 50091 3424 50092 3464
rect 50132 3424 50133 3464
rect 50091 3415 50133 3424
rect 50187 3464 50229 3473
rect 50187 3424 50188 3464
rect 50228 3424 50229 3464
rect 50187 3415 50229 3424
rect 52675 3464 52733 3465
rect 52675 3424 52684 3464
rect 52724 3424 52733 3464
rect 52675 3423 52733 3424
rect 53539 3464 53597 3465
rect 53539 3424 53548 3464
rect 53588 3424 53597 3464
rect 53539 3423 53597 3424
rect 47491 3412 47549 3413
rect 43171 3409 43229 3410
rect 21187 3380 21245 3381
rect 21187 3340 21196 3380
rect 21236 3340 21245 3380
rect 21187 3339 21245 3340
rect 34923 3380 34965 3389
rect 34923 3340 34924 3380
rect 34964 3340 34965 3380
rect 34923 3331 34965 3340
rect 35115 3380 35157 3389
rect 35115 3340 35116 3380
rect 35156 3340 35157 3380
rect 35115 3331 35157 3340
rect 37035 3380 37077 3389
rect 37035 3340 37036 3380
rect 37076 3340 37077 3380
rect 37035 3331 37077 3340
rect 37227 3380 37269 3389
rect 37227 3340 37228 3380
rect 37268 3340 37269 3380
rect 37227 3331 37269 3340
rect 38379 3380 38421 3389
rect 38379 3340 38380 3380
rect 38420 3340 38421 3380
rect 38379 3331 38421 3340
rect 38571 3380 38613 3389
rect 38571 3340 38572 3380
rect 38612 3340 38613 3380
rect 38571 3331 38613 3340
rect 17635 3296 17693 3297
rect 17635 3256 17644 3296
rect 17684 3256 17693 3296
rect 17635 3255 17693 3256
rect 20899 3296 20957 3297
rect 20899 3256 20908 3296
rect 20948 3256 20957 3296
rect 20899 3255 20957 3256
rect 35019 3296 35061 3305
rect 35019 3256 35020 3296
rect 35060 3256 35061 3296
rect 35019 3247 35061 3256
rect 37131 3296 37173 3305
rect 37131 3256 37132 3296
rect 37172 3256 37173 3296
rect 37131 3247 37173 3256
rect 38475 3296 38517 3305
rect 38475 3256 38476 3296
rect 38516 3256 38517 3296
rect 38475 3247 38517 3256
rect 50467 3296 50525 3297
rect 50467 3256 50476 3296
rect 50516 3256 50525 3296
rect 50467 3255 50525 3256
rect 21387 3212 21429 3221
rect 21387 3172 21388 3212
rect 21428 3172 21429 3212
rect 21387 3163 21429 3172
rect 32523 3212 32565 3221
rect 32523 3172 32524 3212
rect 32564 3172 32565 3212
rect 32523 3163 32565 3172
rect 576 3044 80736 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 80736 3044
rect 576 2980 80736 3004
rect 32419 2876 32477 2877
rect 32419 2836 32428 2876
rect 32468 2836 32477 2876
rect 32419 2835 32477 2836
rect 28483 2792 28541 2793
rect 28483 2752 28492 2792
rect 28532 2752 28541 2792
rect 28483 2751 28541 2752
rect 30019 2792 30077 2793
rect 30019 2752 30028 2792
rect 30068 2752 30077 2792
rect 30019 2751 30077 2752
rect 34923 2792 34965 2801
rect 34923 2752 34924 2792
rect 34964 2752 34965 2792
rect 34923 2743 34965 2752
rect 39331 2792 39389 2793
rect 39331 2752 39340 2792
rect 39380 2752 39389 2792
rect 39331 2751 39389 2752
rect 40675 2792 40733 2793
rect 40675 2752 40684 2792
rect 40724 2752 40733 2792
rect 40675 2751 40733 2752
rect 49795 2792 49853 2793
rect 49795 2752 49804 2792
rect 49844 2752 49853 2792
rect 49795 2751 49853 2752
rect 21475 2708 21533 2709
rect 21475 2668 21484 2708
rect 21524 2668 21533 2708
rect 21475 2667 21533 2668
rect 24267 2708 24309 2717
rect 24267 2668 24268 2708
rect 24308 2668 24309 2708
rect 24267 2659 24309 2668
rect 42307 2708 42365 2709
rect 42307 2668 42316 2708
rect 42356 2668 42365 2708
rect 42307 2667 42365 2668
rect 52395 2708 52437 2717
rect 52395 2668 52396 2708
rect 52436 2668 52437 2708
rect 52395 2659 52437 2668
rect 22243 2624 22301 2625
rect 22243 2584 22252 2624
rect 22292 2584 22301 2624
rect 22243 2583 22301 2584
rect 23107 2624 23165 2625
rect 23107 2584 23116 2624
rect 23156 2584 23165 2624
rect 23107 2583 23165 2584
rect 27811 2624 27869 2625
rect 27811 2584 27820 2624
rect 27860 2584 27869 2624
rect 27811 2583 27869 2584
rect 28107 2624 28149 2633
rect 28107 2584 28108 2624
rect 28148 2584 28149 2624
rect 28107 2575 28149 2584
rect 29347 2624 29405 2625
rect 29347 2584 29356 2624
rect 29396 2584 29405 2624
rect 29347 2583 29405 2584
rect 29643 2624 29685 2633
rect 29643 2584 29644 2624
rect 29684 2584 29685 2624
rect 29643 2575 29685 2584
rect 29739 2624 29781 2633
rect 29739 2584 29740 2624
rect 29780 2584 29781 2624
rect 29739 2575 29781 2584
rect 31747 2624 31805 2625
rect 31747 2584 31756 2624
rect 31796 2584 31805 2624
rect 31747 2583 31805 2584
rect 32227 2624 32285 2625
rect 32227 2584 32236 2624
rect 32276 2584 32285 2624
rect 32227 2583 32285 2584
rect 34827 2624 34869 2633
rect 34827 2584 34828 2624
rect 34868 2584 34869 2624
rect 34827 2575 34869 2584
rect 35011 2624 35069 2625
rect 35011 2584 35020 2624
rect 35060 2584 35069 2624
rect 35011 2583 35069 2584
rect 38659 2624 38717 2625
rect 38659 2584 38668 2624
rect 38708 2584 38717 2624
rect 38659 2583 38717 2584
rect 38955 2624 38997 2633
rect 38955 2584 38956 2624
rect 38996 2584 38997 2624
rect 38955 2575 38997 2584
rect 39051 2624 39093 2633
rect 39051 2584 39052 2624
rect 39092 2584 39093 2624
rect 39051 2575 39093 2584
rect 40003 2624 40061 2625
rect 40003 2584 40012 2624
rect 40052 2584 40061 2624
rect 40003 2583 40061 2584
rect 40299 2624 40341 2633
rect 40299 2584 40300 2624
rect 40340 2584 40341 2624
rect 40299 2575 40341 2584
rect 40395 2624 40437 2633
rect 40395 2584 40396 2624
rect 40436 2584 40437 2624
rect 40395 2575 40437 2584
rect 46051 2624 46109 2625
rect 46051 2584 46060 2624
rect 46100 2584 46109 2624
rect 46051 2583 46109 2584
rect 47299 2624 47357 2625
rect 47299 2584 47308 2624
rect 47348 2584 47357 2624
rect 47299 2583 47357 2584
rect 49123 2624 49181 2625
rect 49123 2584 49132 2624
rect 49172 2584 49181 2624
rect 49123 2583 49181 2584
rect 49419 2624 49461 2633
rect 49419 2584 49420 2624
rect 49460 2584 49461 2624
rect 49419 2575 49461 2584
rect 49515 2624 49557 2633
rect 49515 2584 49516 2624
rect 49556 2584 49557 2624
rect 49515 2575 49557 2584
rect 49995 2624 50037 2633
rect 49995 2584 49996 2624
rect 50036 2584 50037 2624
rect 49995 2575 50037 2584
rect 50371 2624 50429 2625
rect 50371 2584 50380 2624
rect 50420 2584 50429 2624
rect 50371 2583 50429 2584
rect 51235 2624 51293 2625
rect 51235 2584 51244 2624
rect 51284 2584 51293 2624
rect 51235 2583 51293 2584
rect 21867 2540 21909 2549
rect 21867 2500 21868 2540
rect 21908 2500 21909 2540
rect 21867 2491 21909 2500
rect 28203 2540 28245 2549
rect 28203 2500 28204 2540
rect 28244 2500 28245 2540
rect 28203 2491 28245 2500
rect 47499 2540 47541 2549
rect 47499 2500 47500 2540
rect 47540 2500 47541 2540
rect 47499 2491 47541 2500
rect 835 2456 893 2457
rect 835 2416 844 2456
rect 884 2416 893 2456
rect 835 2415 893 2416
rect 21675 2456 21717 2465
rect 21675 2416 21676 2456
rect 21716 2416 21717 2456
rect 21675 2407 21717 2416
rect 31651 2456 31709 2457
rect 31651 2416 31660 2456
rect 31700 2416 31709 2456
rect 31651 2415 31709 2416
rect 31939 2456 31997 2457
rect 31939 2416 31948 2456
rect 31988 2416 31997 2456
rect 31939 2415 31997 2416
rect 32131 2456 32189 2457
rect 32131 2416 32140 2456
rect 32180 2416 32189 2456
rect 32131 2415 32189 2416
rect 32715 2456 32757 2465
rect 32715 2416 32716 2456
rect 32756 2416 32757 2456
rect 32715 2407 32757 2416
rect 42507 2456 42549 2465
rect 42507 2416 42508 2456
rect 42548 2416 42549 2456
rect 42507 2407 42549 2416
rect 576 2288 80736 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80736 2288
rect 576 2224 80736 2248
rect 25987 2120 26045 2121
rect 25987 2080 25996 2120
rect 26036 2080 26045 2120
rect 25987 2079 26045 2080
rect 31555 2120 31613 2121
rect 31555 2080 31564 2120
rect 31604 2080 31613 2120
rect 31555 2079 31613 2080
rect 34147 2120 34205 2121
rect 34147 2080 34156 2120
rect 34196 2080 34205 2120
rect 34147 2079 34205 2080
rect 39331 2120 39389 2121
rect 39331 2080 39340 2120
rect 39380 2080 39389 2120
rect 39331 2079 39389 2080
rect 42307 2120 42365 2121
rect 42307 2080 42316 2120
rect 42356 2080 42365 2120
rect 42307 2079 42365 2080
rect 22155 2036 22197 2045
rect 22155 1996 22156 2036
rect 22196 1996 22197 2036
rect 22155 1987 22197 1996
rect 23115 2036 23157 2045
rect 23115 1996 23116 2036
rect 23156 1996 23157 2036
rect 23115 1987 23157 1996
rect 29163 2036 29205 2045
rect 29163 1996 29164 2036
rect 29204 1996 29205 2036
rect 29163 1987 29205 1996
rect 39915 2036 39957 2045
rect 39915 1996 39916 2036
rect 39956 1996 39957 2036
rect 39915 1987 39957 1996
rect 21763 1952 21821 1953
rect 21763 1912 21772 1952
rect 21812 1912 21821 1952
rect 21763 1911 21821 1912
rect 22059 1952 22101 1961
rect 22059 1912 22060 1952
rect 22100 1912 22101 1952
rect 22059 1903 22101 1912
rect 22723 1952 22781 1953
rect 22723 1912 22732 1952
rect 22772 1912 22781 1952
rect 22723 1911 22781 1912
rect 23019 1952 23061 1961
rect 23019 1912 23020 1952
rect 23060 1912 23061 1952
rect 23019 1903 23061 1912
rect 23595 1952 23637 1961
rect 23595 1912 23596 1952
rect 23636 1912 23637 1952
rect 23595 1903 23637 1912
rect 23971 1952 24029 1953
rect 23971 1912 23980 1952
rect 24020 1912 24029 1952
rect 23971 1911 24029 1912
rect 24835 1952 24893 1953
rect 24835 1912 24844 1952
rect 24884 1912 24893 1952
rect 24835 1911 24893 1912
rect 26187 1952 26229 1961
rect 26187 1912 26188 1952
rect 26228 1912 26229 1952
rect 26187 1903 26229 1912
rect 26563 1952 26621 1953
rect 26563 1912 26572 1952
rect 26612 1912 26621 1952
rect 26563 1911 26621 1912
rect 27427 1952 27485 1953
rect 27427 1912 27436 1952
rect 27476 1912 27485 1952
rect 27427 1911 27485 1912
rect 29539 1952 29597 1953
rect 29539 1912 29548 1952
rect 29588 1912 29597 1952
rect 29539 1911 29597 1912
rect 30403 1952 30461 1953
rect 30403 1912 30412 1952
rect 30452 1912 30461 1952
rect 30403 1911 30461 1912
rect 31755 1952 31797 1961
rect 31755 1912 31756 1952
rect 31796 1912 31797 1952
rect 31755 1903 31797 1912
rect 32131 1952 32189 1953
rect 32131 1912 32140 1952
rect 32180 1912 32189 1952
rect 32131 1911 32189 1912
rect 32995 1952 33053 1953
rect 32995 1912 33004 1952
rect 33044 1912 33053 1952
rect 32995 1911 33053 1912
rect 34347 1952 34389 1961
rect 34347 1912 34348 1952
rect 34388 1912 34389 1952
rect 34347 1903 34389 1912
rect 34723 1952 34781 1953
rect 34723 1912 34732 1952
rect 34772 1912 34781 1952
rect 34723 1911 34781 1912
rect 35587 1952 35645 1953
rect 35587 1912 35596 1952
rect 35636 1912 35645 1952
rect 35587 1911 35645 1912
rect 36939 1952 36981 1961
rect 36939 1912 36940 1952
rect 36980 1912 36981 1952
rect 36939 1903 36981 1912
rect 37315 1952 37373 1953
rect 37315 1912 37324 1952
rect 37364 1912 37373 1952
rect 37315 1911 37373 1912
rect 38179 1952 38237 1953
rect 38179 1912 38188 1952
rect 38228 1912 38237 1952
rect 38179 1911 38237 1912
rect 40291 1952 40349 1953
rect 40291 1912 40300 1952
rect 40340 1912 40349 1952
rect 40291 1911 40349 1912
rect 41155 1952 41213 1953
rect 41155 1912 41164 1952
rect 41204 1912 41213 1952
rect 41155 1911 41213 1912
rect 42507 1952 42549 1961
rect 42507 1912 42508 1952
rect 42548 1912 42549 1952
rect 42507 1903 42549 1912
rect 42883 1952 42941 1953
rect 42883 1912 42892 1952
rect 42932 1912 42941 1952
rect 42883 1911 42941 1912
rect 43747 1952 43805 1953
rect 43747 1912 43756 1952
rect 43796 1912 43805 1952
rect 43747 1911 43805 1912
rect 45099 1952 45141 1961
rect 45099 1912 45100 1952
rect 45140 1912 45141 1952
rect 45099 1903 45141 1912
rect 45475 1952 45533 1953
rect 45475 1912 45484 1952
rect 45524 1912 45533 1952
rect 45475 1911 45533 1912
rect 46339 1952 46397 1953
rect 46339 1912 46348 1952
rect 46388 1912 46397 1952
rect 46339 1911 46397 1912
rect 47779 1952 47837 1953
rect 47779 1912 47788 1952
rect 47828 1912 47837 1952
rect 47779 1911 47837 1912
rect 48075 1952 48117 1961
rect 48075 1912 48076 1952
rect 48116 1912 48117 1952
rect 48075 1903 48117 1912
rect 48171 1952 48213 1961
rect 48171 1912 48172 1952
rect 48212 1912 48213 1952
rect 48171 1903 48213 1912
rect 48651 1952 48693 1961
rect 48651 1912 48652 1952
rect 48692 1912 48693 1952
rect 48651 1903 48693 1912
rect 49027 1952 49085 1953
rect 49027 1912 49036 1952
rect 49076 1912 49085 1952
rect 49027 1911 49085 1912
rect 49891 1952 49949 1953
rect 49891 1912 49900 1952
rect 49940 1912 49949 1952
rect 49891 1911 49949 1912
rect 52011 1952 52053 1961
rect 52011 1912 52012 1952
rect 52052 1912 52053 1952
rect 52011 1903 52053 1912
rect 52387 1952 52445 1953
rect 52387 1912 52396 1952
rect 52436 1912 52445 1952
rect 52387 1911 52445 1912
rect 53251 1952 53309 1953
rect 53251 1912 53260 1952
rect 53300 1912 53309 1952
rect 53251 1911 53309 1912
rect 22435 1784 22493 1785
rect 22435 1744 22444 1784
rect 22484 1744 22493 1784
rect 22435 1743 22493 1744
rect 23395 1784 23453 1785
rect 23395 1744 23404 1784
rect 23444 1744 23453 1784
rect 23395 1743 23453 1744
rect 36739 1784 36797 1785
rect 36739 1744 36748 1784
rect 36788 1744 36797 1784
rect 36739 1743 36797 1744
rect 48451 1784 48509 1785
rect 48451 1744 48460 1784
rect 48500 1744 48509 1784
rect 48451 1743 48509 1744
rect 51043 1784 51101 1785
rect 51043 1744 51052 1784
rect 51092 1744 51101 1784
rect 51043 1743 51101 1744
rect 25987 1700 26045 1701
rect 25987 1660 25996 1700
rect 26036 1660 26045 1700
rect 25987 1659 26045 1660
rect 28579 1700 28637 1701
rect 28579 1660 28588 1700
rect 28628 1660 28637 1700
rect 28579 1659 28637 1660
rect 44899 1700 44957 1701
rect 44899 1660 44908 1700
rect 44948 1660 44957 1700
rect 44899 1659 44957 1660
rect 47491 1700 47549 1701
rect 47491 1660 47500 1700
rect 47540 1660 47549 1700
rect 47491 1659 47549 1660
rect 54403 1700 54461 1701
rect 54403 1660 54412 1700
rect 54452 1660 54461 1700
rect 54403 1659 54461 1660
rect 576 1532 80736 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 80736 1532
rect 576 1468 80736 1492
rect 26467 1364 26525 1365
rect 26467 1324 26476 1364
rect 26516 1324 26525 1364
rect 26467 1323 26525 1324
rect 30499 1364 30557 1365
rect 30499 1324 30508 1364
rect 30548 1324 30557 1364
rect 30499 1323 30557 1324
rect 32227 1364 32285 1365
rect 32227 1324 32236 1364
rect 32276 1324 32285 1364
rect 32227 1323 32285 1324
rect 34819 1364 34877 1365
rect 34819 1324 34828 1364
rect 34868 1324 34877 1364
rect 34819 1323 34877 1324
rect 35787 1364 35829 1373
rect 35787 1324 35788 1364
rect 35828 1324 35829 1364
rect 35787 1315 35829 1324
rect 37315 1364 37373 1365
rect 37315 1324 37324 1364
rect 37364 1324 37373 1364
rect 37315 1323 37373 1324
rect 41155 1364 41213 1365
rect 41155 1324 41164 1364
rect 41204 1324 41213 1364
rect 41155 1323 41213 1324
rect 42883 1364 42941 1365
rect 42883 1324 42892 1364
rect 42932 1324 42941 1364
rect 42883 1323 42941 1324
rect 45091 1364 45149 1365
rect 45091 1324 45100 1364
rect 45140 1324 45149 1364
rect 45091 1323 45149 1324
rect 52099 1364 52157 1365
rect 52099 1324 52108 1364
rect 52148 1324 52157 1364
rect 52099 1323 52157 1324
rect 25795 1112 25853 1113
rect 25795 1072 25804 1112
rect 25844 1072 25853 1112
rect 25795 1071 25853 1072
rect 26091 1112 26133 1121
rect 26091 1072 26092 1112
rect 26132 1072 26133 1112
rect 26091 1063 26133 1072
rect 26187 1112 26229 1121
rect 26187 1072 26188 1112
rect 26228 1072 26229 1112
rect 26187 1063 26229 1072
rect 28107 1112 28149 1121
rect 28107 1072 28108 1112
rect 28148 1072 28149 1112
rect 28107 1063 28149 1072
rect 28483 1112 28541 1113
rect 28483 1072 28492 1112
rect 28532 1072 28541 1112
rect 28483 1071 28541 1072
rect 29347 1112 29405 1113
rect 29347 1072 29356 1112
rect 29396 1072 29405 1112
rect 29347 1071 29405 1072
rect 31555 1112 31613 1113
rect 31555 1072 31564 1112
rect 31604 1072 31613 1112
rect 31555 1071 31613 1072
rect 31851 1112 31893 1121
rect 31851 1072 31852 1112
rect 31892 1072 31893 1112
rect 31851 1063 31893 1072
rect 31947 1112 31989 1121
rect 31947 1072 31948 1112
rect 31988 1072 31989 1112
rect 31947 1063 31989 1072
rect 34147 1112 34205 1113
rect 34147 1072 34156 1112
rect 34196 1072 34205 1112
rect 34147 1071 34205 1072
rect 34443 1112 34485 1121
rect 34443 1072 34444 1112
rect 34484 1072 34485 1112
rect 34443 1063 34485 1072
rect 34539 1112 34581 1121
rect 34539 1072 34540 1112
rect 34580 1072 34581 1112
rect 34539 1063 34581 1072
rect 35691 1112 35733 1121
rect 35691 1072 35692 1112
rect 35732 1072 35733 1112
rect 35691 1063 35733 1072
rect 35875 1112 35933 1113
rect 35875 1072 35884 1112
rect 35924 1072 35933 1112
rect 35875 1071 35933 1072
rect 36643 1112 36701 1113
rect 36643 1072 36652 1112
rect 36692 1072 36701 1112
rect 36643 1071 36701 1072
rect 36939 1112 36981 1121
rect 36939 1072 36940 1112
rect 36980 1072 36981 1112
rect 36939 1063 36981 1072
rect 37035 1112 37077 1121
rect 37035 1072 37036 1112
rect 37076 1072 37077 1112
rect 37035 1063 37077 1072
rect 38763 1112 38805 1121
rect 38763 1072 38764 1112
rect 38804 1072 38805 1112
rect 38763 1063 38805 1072
rect 39139 1112 39197 1113
rect 39139 1072 39148 1112
rect 39188 1072 39197 1112
rect 39139 1071 39197 1072
rect 40003 1112 40061 1113
rect 40003 1072 40012 1112
rect 40052 1072 40061 1112
rect 40003 1071 40061 1072
rect 42211 1112 42269 1113
rect 42211 1072 42220 1112
rect 42260 1072 42269 1112
rect 42211 1071 42269 1072
rect 42507 1112 42549 1121
rect 42507 1072 42508 1112
rect 42548 1072 42549 1112
rect 42507 1063 42549 1072
rect 42603 1112 42645 1121
rect 42603 1072 42604 1112
rect 42644 1072 42645 1112
rect 42603 1063 42645 1072
rect 44419 1112 44477 1113
rect 44419 1072 44428 1112
rect 44468 1072 44477 1112
rect 44419 1071 44477 1072
rect 44715 1112 44757 1121
rect 44715 1072 44716 1112
rect 44756 1072 44757 1112
rect 44715 1063 44757 1072
rect 44811 1112 44853 1121
rect 44811 1072 44812 1112
rect 44852 1072 44853 1112
rect 44811 1063 44853 1072
rect 51427 1112 51485 1113
rect 51427 1072 51436 1112
rect 51476 1072 51485 1112
rect 51427 1071 51485 1072
rect 51723 1112 51765 1121
rect 51723 1072 51724 1112
rect 51764 1072 51765 1112
rect 51723 1063 51765 1072
rect 51819 1112 51861 1121
rect 51819 1072 51820 1112
rect 51860 1072 51861 1112
rect 51819 1063 51861 1072
rect 576 776 80736 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80736 776
rect 576 712 80736 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 21004 38368 21044 38408
rect 27148 38368 27188 38408
rect 27052 38284 27092 38324
rect 28972 38284 29012 38324
rect 21100 38200 21140 38240
rect 26860 38200 26900 38240
rect 26956 38200 26996 38240
rect 28492 38200 28532 38240
rect 28876 38200 28916 38240
rect 29260 38200 29300 38240
rect 29452 38200 29492 38240
rect 38476 38200 38516 38240
rect 38764 38200 38804 38240
rect 38860 38200 38900 38240
rect 41068 38200 41108 38240
rect 41356 38200 41396 38240
rect 41452 38200 41492 38240
rect 70348 38200 70388 38240
rect 652 38116 692 38156
rect 21772 38116 21812 38156
rect 23212 38116 23252 38156
rect 23596 38116 23636 38156
rect 23980 38116 24020 38156
rect 844 37948 884 37988
rect 21292 37948 21332 37988
rect 21964 37948 22004 37988
rect 23404 37948 23444 37988
rect 23788 37948 23828 37988
rect 24172 37948 24212 37988
rect 26956 37948 26996 37988
rect 29356 37948 29396 37988
rect 39148 37948 39188 37988
rect 41740 37948 41780 37988
rect 70540 37948 70580 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 26092 37528 26132 37568
rect 41932 37528 41972 37568
rect 19276 37360 19316 37400
rect 19372 37360 19412 37400
rect 20524 37360 20564 37400
rect 21388 37360 21428 37400
rect 23116 37360 23156 37400
rect 23980 37360 24020 37400
rect 25900 37360 25940 37400
rect 26092 37360 26132 37400
rect 26284 37360 26324 37400
rect 26668 37360 26708 37400
rect 27532 37360 27572 37400
rect 29356 37360 29396 37400
rect 29452 37360 29492 37400
rect 30316 37360 30356 37400
rect 31180 37360 31220 37400
rect 38188 37360 38228 37400
rect 39052 37360 39092 37400
rect 41260 37360 41300 37400
rect 41548 37360 41588 37400
rect 42124 37360 42164 37400
rect 42508 37360 42548 37400
rect 43372 37360 43412 37400
rect 20140 37276 20180 37316
rect 22732 37276 22772 37316
rect 29932 37276 29972 37316
rect 37804 37276 37844 37316
rect 41644 37276 41684 37316
rect 19564 37192 19604 37232
rect 22540 37192 22580 37232
rect 25132 37192 25172 37232
rect 28684 37192 28724 37232
rect 29740 37192 29780 37232
rect 32332 37192 32372 37232
rect 40204 37192 40244 37232
rect 44524 37192 44564 37232
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 21772 36914 21812 36954
rect 20620 36856 20660 36896
rect 22636 36856 22676 36896
rect 24364 36856 24404 36896
rect 25228 36856 25268 36896
rect 25996 36856 26036 36896
rect 26956 36856 26996 36896
rect 27244 36856 27284 36896
rect 27628 36856 27668 36896
rect 31468 36856 31508 36896
rect 43468 36856 43508 36896
rect 24652 36772 24692 36812
rect 27916 36772 27956 36812
rect 29068 36772 29108 36812
rect 41068 36772 41108 36812
rect 17836 36688 17876 36728
rect 18220 36688 18260 36728
rect 19084 36688 19124 36728
rect 20428 36688 20468 36728
rect 20716 36688 20756 36728
rect 20908 36688 20948 36728
rect 21580 36688 21620 36728
rect 21676 36688 21716 36728
rect 22252 36688 22292 36728
rect 22348 36688 22388 36728
rect 22924 36688 22964 36728
rect 23020 36688 23060 36728
rect 23212 36688 23252 36728
rect 23308 36688 23348 36728
rect 23500 36688 23540 36728
rect 23692 36688 23732 36728
rect 23884 36688 23924 36728
rect 23980 36688 24020 36728
rect 24460 36688 24500 36728
rect 25228 36688 25268 36728
rect 25324 36688 25364 36728
rect 25900 36688 25940 36728
rect 26092 36688 26132 36728
rect 26188 36688 26228 36728
rect 26476 36688 26516 36728
rect 26572 36688 26612 36728
rect 26668 36688 26708 36728
rect 26764 36688 26804 36728
rect 27148 36688 27188 36728
rect 27340 36688 27380 36728
rect 27436 36688 27476 36728
rect 27724 36688 27764 36728
rect 29452 36688 29492 36728
rect 30316 36688 30356 36728
rect 32428 36688 32468 36728
rect 32812 36688 32852 36728
rect 33676 36688 33716 36728
rect 35116 36688 35156 36728
rect 35404 36688 35444 36728
rect 35500 36688 35540 36728
rect 38476 36688 38516 36728
rect 38860 36688 38900 36728
rect 39724 36688 39764 36728
rect 41452 36688 41492 36728
rect 42316 36688 42356 36728
rect 20236 36604 20276 36644
rect 44908 36604 44948 36644
rect 45292 36604 45332 36644
rect 21292 36520 21332 36560
rect 23500 36520 23540 36560
rect 21004 36436 21044 36476
rect 23692 36436 23732 36476
rect 25516 36436 25556 36476
rect 34828 36436 34868 36476
rect 35788 36436 35828 36476
rect 40876 36436 40916 36476
rect 45100 36436 45140 36476
rect 45484 36436 45524 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 18892 36100 18932 36140
rect 21868 36100 21908 36140
rect 24844 36100 24884 36140
rect 28012 36100 28052 36140
rect 32236 36100 32276 36140
rect 39148 36100 39188 36140
rect 14860 36016 14900 36056
rect 20428 36016 20468 36056
rect 40204 36016 40244 36056
rect 44236 36016 44276 36056
rect 47980 36016 48020 36056
rect 52972 36016 53012 36056
rect 53932 36016 53972 36056
rect 13708 35932 13748 35972
rect 20620 35932 20660 35972
rect 21004 35932 21044 35972
rect 31084 35932 31124 35972
rect 41356 35932 41396 35972
rect 14188 35848 14228 35888
rect 14476 35848 14516 35888
rect 15244 35848 15284 35888
rect 15628 35848 15668 35888
rect 16492 35848 16532 35888
rect 19180 35848 19220 35888
rect 19276 35848 19316 35888
rect 19756 35848 19796 35888
rect 20044 35848 20084 35888
rect 21580 35848 21620 35888
rect 21676 35848 21716 35888
rect 21868 35848 21908 35888
rect 22444 35848 22484 35888
rect 22828 35848 22868 35888
rect 23692 35848 23732 35888
rect 25996 35848 26036 35888
rect 26860 35848 26900 35888
rect 31564 35848 31604 35888
rect 31852 35848 31892 35888
rect 34444 35848 34484 35888
rect 35788 35848 35828 35888
rect 36652 35848 36692 35888
rect 38476 35848 38516 35888
rect 38764 35848 38804 35888
rect 38860 35848 38900 35888
rect 39532 35848 39572 35888
rect 39820 35848 39860 35888
rect 39916 35848 39956 35888
rect 41836 35848 41876 35888
rect 42124 35848 42164 35888
rect 42220 35848 42260 35888
rect 43564 35848 43604 35888
rect 43852 35848 43892 35888
rect 44428 35848 44468 35888
rect 44812 35848 44852 35888
rect 45676 35848 45716 35888
rect 49516 35848 49556 35888
rect 52300 35848 52340 35888
rect 52588 35848 52628 35888
rect 53260 35848 53300 35888
rect 53548 35848 53588 35888
rect 72268 35848 72308 35888
rect 14572 35764 14612 35804
rect 20140 35764 20180 35804
rect 25612 35764 25652 35804
rect 31948 35764 31988 35804
rect 35404 35764 35444 35804
rect 43948 35764 43988 35804
rect 52684 35764 52724 35804
rect 53644 35764 53684 35804
rect 13900 35680 13940 35720
rect 17644 35680 17684 35720
rect 19372 35676 19412 35716
rect 20812 35680 20852 35720
rect 21196 35680 21236 35720
rect 31276 35680 31316 35720
rect 32908 35680 32948 35720
rect 37804 35680 37844 35720
rect 41548 35680 41588 35720
rect 46828 35680 46868 35720
rect 72652 35680 72692 35720
rect 42508 35638 42548 35678
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 17452 35344 17492 35384
rect 21580 35344 21620 35384
rect 27244 35344 27284 35384
rect 27724 35344 27764 35384
rect 32236 35344 32276 35384
rect 43564 35344 43604 35384
rect 18700 35260 18740 35300
rect 28396 35260 28436 35300
rect 29356 35260 29396 35300
rect 44044 35260 44084 35300
rect 53164 35260 53204 35300
rect 13420 35176 13460 35216
rect 13708 35176 13748 35216
rect 13804 35176 13844 35216
rect 14284 35176 14324 35216
rect 14668 35176 14708 35216
rect 15532 35176 15572 35216
rect 17068 35176 17108 35216
rect 18316 35176 18356 35216
rect 18604 35176 18644 35216
rect 19180 35176 19220 35216
rect 19564 35176 19604 35216
rect 20428 35176 20468 35216
rect 24460 35176 24500 35216
rect 25708 35176 25748 35216
rect 26764 35176 26804 35216
rect 27052 35176 27092 35216
rect 28012 35176 28052 35216
rect 28300 35176 28340 35216
rect 28972 35176 29012 35216
rect 29260 35176 29300 35216
rect 29836 35176 29876 35216
rect 30220 35176 30260 35216
rect 31084 35176 31124 35216
rect 33484 35176 33524 35216
rect 34636 35176 34676 35216
rect 35020 35176 35060 35216
rect 35884 35176 35924 35216
rect 37612 35176 37652 35216
rect 38764 35176 38804 35216
rect 39052 35176 39092 35216
rect 39148 35176 39188 35216
rect 40396 35176 40436 35216
rect 40588 35176 40628 35216
rect 40780 35176 40820 35216
rect 41164 35176 41204 35216
rect 42028 35176 42068 35216
rect 43468 35176 43508 35216
rect 43660 35176 43700 35216
rect 43756 35176 43796 35216
rect 44428 35176 44468 35216
rect 45292 35176 45332 35216
rect 46732 35176 46772 35216
rect 47020 35176 47060 35216
rect 47116 35176 47156 35216
rect 47980 35176 48020 35216
rect 48364 35176 48404 35216
rect 49228 35176 49268 35216
rect 50572 35176 50612 35216
rect 50956 35176 50996 35216
rect 51820 35176 51860 35216
rect 53548 35176 53588 35216
rect 54412 35176 54452 35216
rect 12268 35092 12308 35132
rect 27532 35092 27572 35132
rect 47596 35092 47636 35132
rect 14092 35008 14132 35048
rect 18988 35008 19028 35048
rect 29644 35008 29684 35048
rect 12460 34924 12500 34964
rect 16684 34924 16724 34964
rect 17644 34924 17684 34964
rect 24844 34924 24884 34964
rect 26092 34924 26132 34964
rect 28684 34924 28724 34964
rect 32236 34924 32276 34964
rect 33772 34924 33812 34964
rect 37036 34924 37076 34964
rect 37804 34924 37844 34964
rect 39436 34924 39476 34964
rect 40588 34924 40628 34964
rect 43180 34924 43220 34964
rect 46444 34924 46484 34964
rect 47404 34924 47444 34964
rect 47788 34924 47828 34964
rect 50380 34924 50420 34964
rect 52972 34924 53012 34964
rect 55564 34924 55604 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 20332 34588 20372 34628
rect 35500 34588 35540 34628
rect 47212 34588 47252 34628
rect 50764 34588 50804 34628
rect 51916 34588 51956 34628
rect 11596 34504 11636 34544
rect 16300 34504 16340 34544
rect 23404 34504 23444 34544
rect 24460 34504 24500 34544
rect 31948 34504 31988 34544
rect 42892 34504 42932 34544
rect 43372 34504 43412 34544
rect 49804 34504 49844 34544
rect 18892 34420 18932 34460
rect 27052 34420 27092 34460
rect 30412 34420 30452 34460
rect 7372 34336 7412 34376
rect 10924 34336 10964 34376
rect 11212 34336 11252 34376
rect 11788 34336 11828 34376
rect 12172 34336 12212 34376
rect 13036 34336 13076 34376
rect 15244 34336 15284 34376
rect 15628 34336 15668 34376
rect 15916 34336 15956 34376
rect 16012 34336 16052 34376
rect 16492 34336 16532 34376
rect 16876 34336 16916 34376
rect 17740 34336 17780 34376
rect 19852 34336 19892 34376
rect 20812 34336 20852 34376
rect 21004 34336 21044 34376
rect 21388 34336 21428 34376
rect 22252 34336 22292 34376
rect 23788 34336 23828 34376
rect 24076 34336 24116 34376
rect 24652 34336 24692 34376
rect 25036 34336 25076 34376
rect 25900 34336 25940 34376
rect 28012 34336 28052 34376
rect 28396 34336 28436 34376
rect 29260 34336 29300 34376
rect 31276 34336 31316 34376
rect 31564 34336 31604 34376
rect 32140 34336 32180 34376
rect 32524 34336 32564 34376
rect 33388 34336 33428 34376
rect 34828 34336 34868 34376
rect 35116 34336 35156 34376
rect 37324 34336 37364 34376
rect 37708 34336 37748 34376
rect 38572 34336 38612 34376
rect 41068 34336 41108 34376
rect 41260 34336 41300 34376
rect 41356 34336 41396 34376
rect 41644 34336 41684 34376
rect 41836 34336 41876 34376
rect 42220 34336 42260 34376
rect 42700 34336 42740 34376
rect 42892 34336 42932 34376
rect 43756 34336 43796 34376
rect 45196 34336 45236 34376
rect 46540 34336 46580 34376
rect 46828 34336 46868 34376
rect 46924 34336 46964 34376
rect 47404 34336 47444 34376
rect 47788 34336 47828 34376
rect 48652 34336 48692 34376
rect 50092 34336 50132 34376
rect 50380 34336 50420 34376
rect 51532 34336 51572 34376
rect 52780 34336 52820 34376
rect 53644 34336 53684 34376
rect 54124 34336 54164 34376
rect 54508 34336 54548 34376
rect 55372 34336 55412 34376
rect 61516 34336 61556 34376
rect 62476 34336 62516 34376
rect 63340 34336 63380 34376
rect 64684 34336 64724 34376
rect 65932 34336 65972 34376
rect 66892 34336 66932 34376
rect 81196 34336 81236 34376
rect 82060 34336 82100 34376
rect 11308 34252 11348 34292
rect 24172 34252 24212 34292
rect 31660 34252 31700 34292
rect 35212 34252 35252 34292
rect 41164 34252 41204 34292
rect 50476 34252 50516 34292
rect 80812 34252 80852 34292
rect 7756 34168 7796 34208
rect 14188 34168 14228 34208
rect 34540 34168 34580 34208
rect 39724 34168 39764 34208
rect 41740 34168 41780 34208
rect 42316 34168 42356 34208
rect 56524 34168 56564 34208
rect 83212 34168 83252 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 80140 33748 80180 33788
rect 79756 33664 79796 33704
rect 80044 33664 80084 33704
rect 80716 33664 80756 33704
rect 81004 33664 81044 33704
rect 81100 33664 81140 33704
rect 81772 33580 81812 33620
rect 80428 33496 80468 33536
rect 81388 33412 81428 33452
rect 81964 33412 82004 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 5644 33076 5684 33116
rect 5452 32908 5492 32948
rect 80428 32908 80468 32948
rect 80812 32824 80852 32864
rect 81196 32824 81236 32864
rect 82060 32824 82100 32864
rect 5644 32656 5684 32696
rect 80620 32656 80660 32696
rect 83212 32656 83252 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 83212 32320 83252 32360
rect 4972 32152 5012 32192
rect 80812 32152 80852 32192
rect 81196 32152 81236 32192
rect 82060 32152 82100 32192
rect 4396 32068 4436 32108
rect 4588 31900 4628 31940
rect 5164 31900 5204 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 81388 31564 81428 31604
rect 5836 31396 5876 31436
rect 81676 31396 81716 31436
rect 3820 31312 3860 31352
rect 4684 31312 4724 31352
rect 80716 31312 80756 31352
rect 81004 31312 81044 31352
rect 81100 31312 81140 31352
rect 3436 31228 3476 31268
rect 81868 31144 81908 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 83212 30808 83252 30848
rect 4876 30724 4916 30764
rect 4492 30640 4532 30680
rect 4780 30640 4820 30680
rect 80812 30640 80852 30680
rect 81196 30640 81236 30680
rect 82060 30640 82100 30680
rect 79948 30556 79988 30596
rect 5164 30472 5204 30512
rect 80140 30388 80180 30428
rect 83212 30388 83252 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 82444 30052 82484 30092
rect 79852 29968 79892 30008
rect 79180 29800 79220 29840
rect 79468 29800 79508 29840
rect 79564 29800 79604 29840
rect 80044 29800 80084 29840
rect 80428 29800 80468 29840
rect 81292 29800 81332 29840
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 80428 29212 80468 29252
rect 80044 29128 80084 29168
rect 80332 29128 80372 29168
rect 81004 29128 81044 29168
rect 81292 29128 81332 29168
rect 81388 29128 81428 29168
rect 80716 28960 80756 29000
rect 81676 28876 81716 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 82636 28540 82676 28580
rect 80044 28456 80084 28496
rect 74764 28288 74804 28328
rect 76108 28288 76148 28328
rect 79372 28288 79412 28328
rect 79660 28288 79700 28328
rect 79756 28288 79796 28328
rect 80236 28288 80276 28328
rect 80620 28288 80660 28328
rect 81484 28288 81524 28328
rect 82636 28120 82676 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 83212 27784 83252 27824
rect 80812 27700 80852 27740
rect 3436 27616 3476 27656
rect 3820 27616 3860 27656
rect 4684 27616 4724 27656
rect 81196 27616 81236 27656
rect 82060 27616 82100 27656
rect 5836 27364 5876 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 5164 27028 5204 27068
rect 82828 27028 82868 27068
rect 4492 26776 4532 26816
rect 4780 26776 4820 26816
rect 80812 26776 80852 26816
rect 81676 26776 81716 26816
rect 4876 26692 4916 26732
rect 80428 26692 80468 26732
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 80620 26188 80660 26228
rect 80236 26104 80276 26144
rect 80524 26104 80564 26144
rect 81292 26104 81332 26144
rect 81580 26104 81620 26144
rect 81676 26104 81716 26144
rect 80908 25936 80948 25976
rect 81964 25852 82004 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 5836 25516 5876 25556
rect 83212 25516 83252 25556
rect 80620 25432 80660 25472
rect 652 25348 692 25388
rect 3820 25264 3860 25304
rect 4684 25264 4724 25304
rect 79948 25264 79988 25304
rect 80236 25264 80276 25304
rect 80812 25264 80852 25304
rect 81196 25264 81236 25304
rect 82060 25264 82100 25304
rect 3436 25180 3476 25220
rect 80332 25180 80372 25220
rect 844 25096 884 25136
rect 5836 25096 5876 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 5068 24802 5108 24842
rect 4780 24676 4820 24716
rect 80524 24676 80564 24716
rect 4396 24592 4436 24632
rect 4684 24592 4724 24632
rect 74092 24592 74132 24632
rect 80908 24592 80948 24632
rect 81772 24592 81812 24632
rect 652 24508 692 24548
rect 82924 24508 82964 24548
rect 844 24424 884 24464
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 844 24004 884 24044
rect 652 23836 692 23876
rect 74188 23752 74228 23792
rect 74668 23584 74708 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 844 23248 884 23288
rect 3436 23080 3476 23120
rect 3820 23080 3860 23120
rect 4684 23080 4724 23120
rect 74188 23080 74228 23120
rect 652 22996 692 23036
rect 5836 22828 5876 22868
rect 74476 22828 74516 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 4396 22492 4436 22532
rect 3724 22240 3764 22280
rect 4012 22240 4052 22280
rect 4108 22240 4148 22280
rect 844 22072 884 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3436 21568 3476 21608
rect 3820 21568 3860 21608
rect 4684 21568 4724 21608
rect 82732 21568 82772 21608
rect 83116 21568 83156 21608
rect 83980 21568 84020 21608
rect 5836 21484 5876 21524
rect 85132 21316 85172 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 82348 20980 82388 21020
rect 2764 20896 2804 20936
rect 2092 20728 2132 20768
rect 2380 20728 2420 20768
rect 2956 20728 2996 20768
rect 3340 20728 3380 20768
rect 4204 20728 4244 20768
rect 81676 20728 81716 20768
rect 81964 20728 82004 20768
rect 82060 20728 82100 20768
rect 2476 20644 2516 20684
rect 844 20560 884 20600
rect 5356 20560 5396 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 844 20224 884 20264
rect 4300 20140 4340 20180
rect 1228 20056 1268 20096
rect 1612 20056 1652 20096
rect 2476 20056 2516 20096
rect 3916 20056 3956 20096
rect 4204 20056 4244 20096
rect 98380 20056 98420 20096
rect 4588 19888 4628 19928
rect 96844 19888 96884 19928
rect 3628 19804 3668 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 2284 19468 2324 19508
rect 5068 19468 5108 19508
rect 4684 19384 4724 19424
rect 2476 19300 2516 19340
rect 3532 19300 3572 19340
rect 4876 19300 4916 19340
rect 1612 19216 1652 19256
rect 1900 19216 1940 19256
rect 1996 19216 2036 19256
rect 4012 19216 4052 19256
rect 4300 19216 4340 19256
rect 4396 19216 4436 19256
rect 844 19048 884 19088
rect 2668 19048 2708 19088
rect 3724 19048 3764 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 844 18712 884 18752
rect 3436 18628 3476 18668
rect 3820 18544 3860 18584
rect 4684 18544 4724 18584
rect 1900 18460 1940 18500
rect 2284 18460 2324 18500
rect 5836 18460 5876 18500
rect 2092 18376 2132 18416
rect 2476 18292 2516 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 4492 17956 4532 17996
rect 1516 17872 1556 17912
rect 4108 17872 4148 17912
rect 4300 17788 4340 17828
rect 844 17704 884 17744
rect 1132 17704 1172 17744
rect 1228 17704 1268 17744
rect 1708 17704 1748 17744
rect 2092 17704 2132 17744
rect 2956 17704 2996 17744
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 844 17200 884 17240
rect 1228 17200 1268 17240
rect 80620 17200 80660 17240
rect 77740 17116 77780 17156
rect 3436 17032 3476 17072
rect 3820 17032 3860 17072
rect 4684 17032 4724 17072
rect 77356 17032 77396 17072
rect 77644 17032 77684 17072
rect 78220 17032 78260 17072
rect 78604 17032 78644 17072
rect 79468 17032 79508 17072
rect 78028 16864 78068 16904
rect 5836 16780 5876 16820
rect 80620 16780 80660 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 4012 16444 4052 16484
rect 4972 16444 5012 16484
rect 1996 16192 2036 16232
rect 2860 16192 2900 16232
rect 4300 16192 4340 16232
rect 4588 16192 4628 16232
rect 4684 16192 4724 16232
rect 1612 16108 1652 16148
rect 844 16024 884 16064
rect 4012 16024 4052 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 5836 15688 5876 15728
rect 1516 15520 1556 15560
rect 1804 15520 1844 15560
rect 1900 15520 1940 15560
rect 3436 15520 3476 15560
rect 3820 15520 3860 15560
rect 4684 15520 4724 15560
rect 652 15436 692 15476
rect 2188 15352 2228 15392
rect 844 15268 884 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 4972 14932 5012 14972
rect 4012 14848 4052 14888
rect 652 14764 692 14804
rect 1996 14680 2036 14720
rect 2860 14680 2900 14720
rect 4300 14680 4340 14720
rect 4588 14680 4628 14720
rect 4684 14680 4724 14720
rect 1612 14596 1652 14636
rect 844 14512 884 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 1516 14008 1556 14048
rect 1804 14008 1844 14048
rect 1900 14008 1940 14048
rect 3628 14008 3668 14048
rect 3916 14008 3956 14048
rect 4012 14008 4052 14048
rect 2188 13840 2228 13880
rect 4300 13756 4340 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 5836 13420 5876 13460
rect 1228 13168 1268 13208
rect 2092 13168 2132 13208
rect 3436 13168 3476 13208
rect 3820 13168 3860 13208
rect 4684 13168 4724 13208
rect 844 13084 884 13124
rect 3244 13000 3284 13040
rect 5836 13000 5876 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 844 12664 884 12704
rect 2188 12706 2228 12746
rect 1516 12496 1556 12536
rect 1804 12496 1844 12536
rect 1900 12496 1940 12536
rect 3436 12496 3476 12536
rect 3820 12496 3860 12536
rect 4684 12496 4724 12536
rect 652 12412 692 12452
rect 1036 12412 1076 12452
rect 1228 12328 1268 12368
rect 5836 12244 5876 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 4588 11908 4628 11948
rect 652 11740 692 11780
rect 3916 11656 3956 11696
rect 4204 11656 4244 11696
rect 4300 11656 4340 11696
rect 844 11488 884 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 2380 11194 2420 11234
rect 4972 11152 5012 11192
rect 2092 11068 2132 11108
rect 2572 11068 2612 11108
rect 1708 10984 1748 11024
rect 1996 10984 2036 11024
rect 2956 10984 2996 11024
rect 3820 10984 3860 11024
rect 652 10900 692 10940
rect 844 10732 884 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 652 10228 692 10268
rect 5836 10228 5876 10268
rect 3820 10144 3860 10184
rect 4684 10144 4724 10184
rect 3436 10060 3476 10100
rect 844 9976 884 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 4012 9472 4052 9512
rect 4300 9472 4340 9512
rect 4396 9472 4436 9512
rect 652 9388 692 9428
rect 4684 9304 4724 9344
rect 844 9220 884 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 844 8464 884 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 844 8128 884 8168
rect 5836 8128 5876 8168
rect 3436 7960 3476 8000
rect 3820 7960 3860 8000
rect 4684 7960 4724 8000
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 5068 7372 5108 7412
rect 4396 7120 4436 7160
rect 4684 7120 4724 7160
rect 4780 7120 4820 7160
rect 844 6952 884 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 80236 6448 80276 6488
rect 78892 6364 78932 6404
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 844 5440 884 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 844 5104 884 5144
rect 18412 5104 18452 5144
rect 31948 5104 31988 5144
rect 32140 5104 32180 5144
rect 32716 5104 32756 5144
rect 21772 5020 21812 5060
rect 26092 5020 26132 5060
rect 39244 5020 39284 5060
rect 16012 4936 16052 4976
rect 16396 4936 16436 4976
rect 17260 4925 17300 4965
rect 21388 4936 21428 4976
rect 21676 4936 21716 4976
rect 24076 4936 24116 4976
rect 24364 4936 24404 4976
rect 24460 4936 24500 4976
rect 25708 4936 25748 4976
rect 25996 4936 26036 4976
rect 30316 4936 30356 4976
rect 30604 4936 30644 4976
rect 30700 4936 30740 4976
rect 32236 4936 32276 4976
rect 36940 4936 36980 4976
rect 37132 4936 37172 4976
rect 38572 4936 38612 4976
rect 38956 4936 38996 4976
rect 39148 4936 39188 4976
rect 39340 4936 39380 4976
rect 45196 4936 45236 4976
rect 51724 4936 51764 4976
rect 52012 4936 52052 4976
rect 52108 4936 52148 4976
rect 25228 4852 25268 4892
rect 26572 4852 26612 4892
rect 26956 4852 26996 4892
rect 38668 4852 38708 4892
rect 38860 4852 38900 4892
rect 43852 4852 43892 4892
rect 46828 4852 46868 4892
rect 25420 4768 25460 4808
rect 32428 4768 32468 4808
rect 38764 4768 38804 4808
rect 22060 4684 22100 4724
rect 24748 4684 24788 4724
rect 26380 4684 26420 4724
rect 26764 4684 26804 4724
rect 27148 4684 27188 4724
rect 30988 4684 31028 4724
rect 37036 4684 37076 4724
rect 47020 4684 47060 4724
rect 52396 4684 52436 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 17260 4348 17300 4388
rect 22444 4348 22484 4388
rect 19852 4264 19892 4304
rect 27052 4264 27092 4304
rect 30892 4264 30932 4304
rect 36364 4264 36404 4304
rect 38668 4264 38708 4304
rect 41260 4264 41300 4304
rect 46540 4264 46580 4304
rect 47788 4264 47828 4304
rect 54028 4264 54068 4304
rect 50380 4180 50420 4220
rect 16588 4096 16628 4136
rect 16876 4096 16916 4136
rect 16972 4096 17012 4136
rect 17836 4096 17876 4136
rect 18700 4096 18740 4136
rect 20428 4096 20468 4136
rect 21292 4096 21332 4136
rect 23404 4096 23444 4136
rect 23788 4096 23828 4136
rect 24652 4096 24692 4136
rect 26380 4096 26420 4136
rect 26668 4096 26708 4136
rect 26764 4096 26804 4136
rect 27244 4096 27284 4136
rect 27628 4096 27668 4136
rect 28492 4096 28532 4136
rect 30220 4096 30260 4136
rect 30508 4096 30548 4136
rect 31084 4096 31124 4136
rect 31468 4096 31508 4136
rect 32332 4096 32372 4136
rect 34732 4096 34772 4136
rect 35116 4096 35156 4136
rect 35308 4096 35348 4136
rect 36268 4096 36308 4136
rect 36460 4096 36500 4136
rect 40012 4096 40052 4136
rect 40108 4096 40148 4136
rect 40684 4096 40724 4136
rect 40780 4096 40820 4136
rect 40876 4096 40916 4136
rect 40972 4096 41012 4136
rect 42316 4096 42356 4136
rect 42508 4096 42548 4136
rect 42796 4096 42836 4136
rect 42892 4096 42932 4136
rect 43276 4096 43316 4136
rect 43372 4096 43412 4136
rect 43852 4096 43892 4136
rect 44332 4101 44372 4141
rect 45868 4096 45908 4136
rect 46156 4096 46196 4136
rect 47116 4096 47156 4136
rect 47500 4138 47540 4178
rect 47404 4096 47444 4136
rect 47980 4096 48020 4136
rect 48364 4096 48404 4136
rect 49228 4096 49268 4136
rect 50956 4096 50996 4136
rect 51820 4096 51860 4136
rect 53356 4096 53396 4136
rect 53644 4096 53684 4136
rect 54220 4096 54260 4136
rect 54604 4096 54644 4136
rect 55468 4096 55508 4136
rect 17452 4012 17492 4052
rect 20044 4012 20084 4052
rect 30604 4012 30644 4052
rect 46252 4012 46292 4052
rect 50572 4012 50612 4052
rect 53740 4012 53780 4052
rect 844 3928 884 3968
rect 25804 3928 25844 3968
rect 29644 3928 29684 3968
rect 33484 3928 33524 3968
rect 34636 3928 34676 3968
rect 34924 3928 34964 3968
rect 35212 3928 35252 3968
rect 40300 3928 40340 3968
rect 42412 3928 42452 3968
rect 44524 3928 44564 3968
rect 52972 3928 53012 3968
rect 56620 3928 56660 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 844 3592 884 3632
rect 23980 3592 24020 3632
rect 28588 3592 28628 3632
rect 31948 3592 31988 3632
rect 32428 3592 32468 3632
rect 41260 3592 41300 3632
rect 48652 3592 48692 3632
rect 54700 3592 54740 3632
rect 17356 3508 17396 3548
rect 20620 3508 20660 3548
rect 21580 3508 21620 3548
rect 26188 3508 26228 3548
rect 29548 3508 29588 3548
rect 43084 3508 43124 3548
rect 45388 3508 45428 3548
rect 46252 3508 46292 3548
rect 52300 3508 52340 3548
rect 16972 3424 17012 3464
rect 17260 3451 17300 3491
rect 20236 3424 20276 3464
rect 20524 3424 20564 3464
rect 21964 3424 22004 3464
rect 22828 3424 22868 3464
rect 26572 3424 26612 3464
rect 27436 3424 27476 3464
rect 29932 3424 29972 3464
rect 30796 3424 30836 3464
rect 32236 3424 32276 3464
rect 32524 3424 32564 3464
rect 34828 3424 34868 3464
rect 35212 3424 35252 3464
rect 36940 3424 36980 3464
rect 37324 3424 37364 3464
rect 38284 3424 38324 3464
rect 38668 3424 38708 3464
rect 40972 3424 41012 3464
rect 41068 3424 41108 3464
rect 41164 3424 41204 3464
rect 42988 3424 43028 3464
rect 43180 3410 43220 3450
rect 43276 3424 43316 3464
rect 43948 3424 43988 3464
rect 45196 3424 45236 3464
rect 46636 3424 46676 3464
rect 47500 3413 47540 3453
rect 49804 3424 49844 3464
rect 50092 3424 50132 3464
rect 50188 3424 50228 3464
rect 52684 3424 52724 3464
rect 53548 3424 53588 3464
rect 21196 3340 21236 3380
rect 34924 3340 34964 3380
rect 35116 3340 35156 3380
rect 37036 3340 37076 3380
rect 37228 3340 37268 3380
rect 38380 3340 38420 3380
rect 38572 3340 38612 3380
rect 17644 3256 17684 3296
rect 20908 3256 20948 3296
rect 35020 3256 35060 3296
rect 37132 3256 37172 3296
rect 38476 3256 38516 3296
rect 50476 3256 50516 3296
rect 21388 3172 21428 3212
rect 32524 3172 32564 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 32428 2836 32468 2876
rect 28492 2752 28532 2792
rect 30028 2752 30068 2792
rect 34924 2752 34964 2792
rect 39340 2752 39380 2792
rect 40684 2752 40724 2792
rect 49804 2752 49844 2792
rect 21484 2668 21524 2708
rect 24268 2668 24308 2708
rect 42316 2668 42356 2708
rect 52396 2668 52436 2708
rect 22252 2584 22292 2624
rect 23116 2584 23156 2624
rect 27820 2584 27860 2624
rect 28108 2584 28148 2624
rect 29356 2584 29396 2624
rect 29644 2584 29684 2624
rect 29740 2584 29780 2624
rect 31756 2584 31796 2624
rect 32236 2584 32276 2624
rect 34828 2584 34868 2624
rect 35020 2584 35060 2624
rect 38668 2584 38708 2624
rect 38956 2584 38996 2624
rect 39052 2584 39092 2624
rect 40012 2584 40052 2624
rect 40300 2584 40340 2624
rect 40396 2584 40436 2624
rect 46060 2584 46100 2624
rect 47308 2584 47348 2624
rect 49132 2584 49172 2624
rect 49420 2584 49460 2624
rect 49516 2584 49556 2624
rect 49996 2584 50036 2624
rect 50380 2584 50420 2624
rect 51244 2584 51284 2624
rect 21868 2500 21908 2540
rect 28204 2500 28244 2540
rect 47500 2500 47540 2540
rect 844 2416 884 2456
rect 21676 2416 21716 2456
rect 31660 2416 31700 2456
rect 31948 2416 31988 2456
rect 32140 2416 32180 2456
rect 32716 2416 32756 2456
rect 42508 2416 42548 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 25996 2080 26036 2120
rect 31564 2080 31604 2120
rect 34156 2080 34196 2120
rect 39340 2080 39380 2120
rect 42316 2080 42356 2120
rect 22156 1996 22196 2036
rect 23116 1996 23156 2036
rect 29164 1996 29204 2036
rect 39916 1996 39956 2036
rect 21772 1912 21812 1952
rect 22060 1912 22100 1952
rect 22732 1912 22772 1952
rect 23020 1912 23060 1952
rect 23596 1912 23636 1952
rect 23980 1912 24020 1952
rect 24844 1912 24884 1952
rect 26188 1912 26228 1952
rect 26572 1912 26612 1952
rect 27436 1912 27476 1952
rect 29548 1912 29588 1952
rect 30412 1912 30452 1952
rect 31756 1912 31796 1952
rect 32140 1912 32180 1952
rect 33004 1912 33044 1952
rect 34348 1912 34388 1952
rect 34732 1912 34772 1952
rect 35596 1912 35636 1952
rect 36940 1912 36980 1952
rect 37324 1912 37364 1952
rect 38188 1912 38228 1952
rect 40300 1912 40340 1952
rect 41164 1912 41204 1952
rect 42508 1912 42548 1952
rect 42892 1912 42932 1952
rect 43756 1912 43796 1952
rect 45100 1912 45140 1952
rect 45484 1912 45524 1952
rect 46348 1912 46388 1952
rect 47788 1912 47828 1952
rect 48076 1912 48116 1952
rect 48172 1912 48212 1952
rect 48652 1912 48692 1952
rect 49036 1912 49076 1952
rect 49900 1912 49940 1952
rect 52012 1912 52052 1952
rect 52396 1912 52436 1952
rect 53260 1912 53300 1952
rect 22444 1744 22484 1784
rect 23404 1744 23444 1784
rect 36748 1744 36788 1784
rect 48460 1744 48500 1784
rect 51052 1744 51092 1784
rect 25996 1660 26036 1700
rect 28588 1660 28628 1700
rect 44908 1660 44948 1700
rect 47500 1660 47540 1700
rect 54412 1660 54452 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 26476 1324 26516 1364
rect 30508 1324 30548 1364
rect 32236 1324 32276 1364
rect 34828 1324 34868 1364
rect 35788 1324 35828 1364
rect 37324 1324 37364 1364
rect 41164 1324 41204 1364
rect 42892 1324 42932 1364
rect 45100 1324 45140 1364
rect 52108 1324 52148 1364
rect 25804 1072 25844 1112
rect 26092 1072 26132 1112
rect 26188 1072 26228 1112
rect 28108 1072 28148 1112
rect 28492 1072 28532 1112
rect 29356 1072 29396 1112
rect 31564 1072 31604 1112
rect 31852 1072 31892 1112
rect 31948 1072 31988 1112
rect 34156 1072 34196 1112
rect 34444 1072 34484 1112
rect 34540 1072 34580 1112
rect 35692 1072 35732 1112
rect 35884 1072 35924 1112
rect 36652 1072 36692 1112
rect 36940 1072 36980 1112
rect 37036 1072 37076 1112
rect 38764 1072 38804 1112
rect 39148 1072 39188 1112
rect 40012 1072 40052 1112
rect 42220 1072 42260 1112
rect 42508 1072 42548 1112
rect 42604 1072 42644 1112
rect 44428 1072 44468 1112
rect 44716 1072 44756 1112
rect 44812 1072 44852 1112
rect 51436 1072 51476 1112
rect 51724 1072 51764 1112
rect 51820 1072 51860 1112
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 21003 38408 21045 38417
rect 21003 38368 21004 38408
rect 21044 38368 21045 38408
rect 21003 38359 21045 38368
rect 22251 38408 22293 38417
rect 27148 38408 27188 38417
rect 22251 38368 22252 38408
rect 22292 38368 22293 38408
rect 22251 38359 22293 38368
rect 26764 38368 26996 38408
rect 21004 38274 21044 38359
rect 21100 38240 21140 38249
rect 652 38156 692 38165
rect 652 37577 692 38116
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 5451 37988 5493 37997
rect 5451 37948 5452 37988
rect 5492 37948 5493 37988
rect 5451 37939 5493 37948
rect 844 37854 884 37939
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 651 37568 693 37577
rect 651 37528 652 37568
rect 692 37528 693 37568
rect 651 37519 693 37528
rect 747 37400 789 37409
rect 747 37360 748 37400
rect 788 37360 789 37400
rect 747 37351 789 37360
rect 652 25388 692 25397
rect 652 24977 692 25348
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 652 24548 692 24557
rect 652 24137 692 24508
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 652 23876 692 23885
rect 652 23297 692 23836
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 748 23288 788 37351
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 5452 36233 5492 37939
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 19276 37400 19316 37409
rect 19180 37360 19276 37400
rect 7083 36728 7125 36737
rect 7083 36688 7084 36728
rect 7124 36688 7125 36728
rect 7083 36679 7125 36688
rect 17835 36728 17877 36737
rect 18220 36728 18260 36737
rect 17835 36688 17836 36728
rect 17876 36688 17877 36728
rect 17835 36679 17877 36688
rect 18124 36688 18220 36728
rect 5451 36224 5493 36233
rect 5451 36184 5452 36224
rect 5492 36184 5493 36224
rect 5451 36175 5493 36184
rect 2571 35888 2613 35897
rect 2571 35848 2572 35888
rect 2612 35848 2613 35888
rect 2571 35839 2613 35848
rect 1131 33788 1173 33797
rect 1131 33748 1132 33788
rect 1172 33748 1173 33788
rect 1131 33739 1173 33748
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 844 25002 884 25087
rect 844 24464 884 24473
rect 884 24424 1076 24464
rect 844 24415 884 24424
rect 843 24044 885 24053
rect 843 24004 844 24044
rect 884 24004 885 24044
rect 843 23995 885 24004
rect 844 23910 884 23995
rect 844 23288 884 23297
rect 748 23248 844 23288
rect 651 23239 693 23248
rect 844 23239 884 23248
rect 652 23036 692 23045
rect 652 22457 692 22996
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 844 22112 884 22121
rect 844 21617 884 22072
rect 843 21608 885 21617
rect 843 21568 844 21608
rect 884 21568 885 21608
rect 843 21559 885 21568
rect 843 20768 885 20777
rect 843 20728 844 20768
rect 884 20728 885 20768
rect 843 20719 885 20728
rect 844 20600 884 20719
rect 844 20551 884 20560
rect 844 20264 884 20273
rect 844 19937 884 20224
rect 843 19928 885 19937
rect 843 19888 844 19928
rect 884 19888 885 19928
rect 843 19879 885 19888
rect 843 19088 885 19097
rect 843 19048 844 19088
rect 884 19048 885 19088
rect 843 19039 885 19048
rect 844 18954 884 19039
rect 844 18752 884 18761
rect 844 18257 884 18712
rect 843 18248 885 18257
rect 843 18208 844 18248
rect 884 18208 885 18248
rect 843 18199 885 18208
rect 843 18080 885 18089
rect 843 18040 844 18080
rect 884 18040 885 18080
rect 843 18031 885 18040
rect 844 17744 884 18031
rect 844 17695 884 17704
rect 843 17408 885 17417
rect 843 17368 844 17408
rect 884 17368 885 17408
rect 843 17359 885 17368
rect 844 17240 884 17359
rect 1036 17300 1076 24424
rect 1132 24053 1172 33739
rect 1323 25136 1365 25145
rect 1323 25096 1324 25136
rect 1364 25096 1365 25136
rect 1323 25087 1365 25096
rect 1131 24044 1173 24053
rect 1131 24004 1132 24044
rect 1172 24004 1173 24044
rect 1131 23995 1173 24004
rect 1227 20096 1269 20105
rect 1227 20056 1228 20096
rect 1268 20056 1269 20096
rect 1227 20047 1269 20056
rect 1228 19962 1268 20047
rect 1227 17912 1269 17921
rect 1227 17872 1228 17912
rect 1268 17872 1269 17912
rect 1227 17863 1269 17872
rect 844 17191 884 17200
rect 940 17260 1076 17300
rect 1132 17744 1172 17753
rect 844 16064 884 16073
rect 844 15737 884 16024
rect 843 15728 885 15737
rect 843 15688 844 15728
rect 884 15688 885 15728
rect 843 15679 885 15688
rect 651 15476 693 15485
rect 651 15436 652 15476
rect 692 15436 693 15476
rect 651 15427 693 15436
rect 652 15342 692 15427
rect 844 15308 884 15317
rect 844 14897 884 15268
rect 843 14888 885 14897
rect 843 14848 844 14888
rect 884 14848 885 14888
rect 843 14839 885 14848
rect 652 14804 692 14813
rect 556 14764 652 14804
rect 556 5489 596 14764
rect 652 14755 692 14764
rect 844 14552 884 14561
rect 844 14057 884 14512
rect 843 14048 885 14057
rect 843 14008 844 14048
rect 884 14008 885 14048
rect 843 13999 885 14008
rect 747 13208 789 13217
rect 747 13168 748 13208
rect 788 13168 789 13208
rect 747 13159 789 13168
rect 748 12704 788 13159
rect 844 13124 884 13133
rect 844 12881 884 13084
rect 843 12872 885 12881
rect 843 12832 844 12872
rect 884 12832 885 12872
rect 843 12823 885 12832
rect 844 12704 884 12713
rect 748 12664 844 12704
rect 844 12655 884 12664
rect 651 12452 693 12461
rect 651 12412 652 12452
rect 692 12412 693 12452
rect 651 12403 693 12412
rect 652 12318 692 12403
rect 940 12242 980 17260
rect 1132 16073 1172 17704
rect 1228 17744 1268 17863
rect 1228 17695 1268 17704
rect 1228 17240 1268 17249
rect 1228 16577 1268 17200
rect 1227 16568 1269 16577
rect 1227 16528 1228 16568
rect 1268 16528 1269 16568
rect 1227 16519 1269 16528
rect 1131 16064 1173 16073
rect 1131 16024 1132 16064
rect 1172 16024 1173 16064
rect 1131 16015 1173 16024
rect 1227 14384 1269 14393
rect 1227 14344 1228 14384
rect 1268 14344 1269 14384
rect 1227 14335 1269 14344
rect 1228 13385 1268 14335
rect 1227 13376 1269 13385
rect 1227 13336 1228 13376
rect 1268 13336 1269 13376
rect 1227 13327 1269 13336
rect 1228 13208 1268 13327
rect 1228 13159 1268 13168
rect 1036 12452 1076 12461
rect 1076 12412 1172 12452
rect 1036 12403 1076 12412
rect 940 12202 1076 12242
rect 651 11780 693 11789
rect 651 11740 652 11780
rect 692 11740 693 11780
rect 651 11731 693 11740
rect 652 11646 692 11731
rect 843 11528 885 11537
rect 843 11488 844 11528
rect 884 11488 885 11528
rect 843 11479 885 11488
rect 844 11394 884 11479
rect 651 10940 693 10949
rect 651 10900 652 10940
rect 692 10900 693 10940
rect 651 10891 693 10900
rect 652 10806 692 10891
rect 843 10772 885 10781
rect 843 10732 844 10772
rect 884 10732 885 10772
rect 843 10723 885 10732
rect 844 10638 884 10723
rect 651 10268 693 10277
rect 651 10228 652 10268
rect 692 10228 693 10268
rect 651 10219 693 10228
rect 939 10268 981 10277
rect 939 10228 940 10268
rect 980 10228 981 10268
rect 939 10219 981 10228
rect 652 10134 692 10219
rect 844 10016 884 10025
rect 844 9857 884 9976
rect 843 9848 885 9857
rect 843 9808 844 9848
rect 884 9808 885 9848
rect 843 9799 885 9808
rect 652 9428 692 9437
rect 555 5480 597 5489
rect 555 5440 556 5480
rect 596 5440 597 5480
rect 555 5431 597 5440
rect 652 4901 692 9388
rect 844 9260 884 9269
rect 844 9017 884 9220
rect 843 9008 885 9017
rect 843 8968 844 9008
rect 884 8968 885 9008
rect 843 8959 885 8968
rect 844 8504 884 8513
rect 748 8464 844 8504
rect 748 8177 788 8464
rect 844 8455 884 8464
rect 747 8168 789 8177
rect 747 8128 748 8168
rect 788 8128 789 8168
rect 747 8119 789 8128
rect 844 8168 884 8177
rect 844 7337 884 8128
rect 843 7328 885 7337
rect 843 7288 844 7328
rect 884 7288 885 7328
rect 843 7279 885 7288
rect 844 6992 884 7001
rect 844 6497 884 6952
rect 843 6488 885 6497
rect 843 6448 844 6488
rect 884 6448 885 6488
rect 843 6439 885 6448
rect 843 5648 885 5657
rect 843 5608 844 5648
rect 884 5608 885 5648
rect 843 5599 885 5608
rect 844 5480 884 5599
rect 844 5431 884 5440
rect 844 5144 884 5153
rect 651 4892 693 4901
rect 651 4852 652 4892
rect 692 4852 693 4892
rect 651 4843 693 4852
rect 844 4817 884 5104
rect 843 4808 885 4817
rect 843 4768 844 4808
rect 884 4768 885 4808
rect 843 4759 885 4768
rect 843 3968 885 3977
rect 843 3928 844 3968
rect 884 3928 885 3968
rect 843 3919 885 3928
rect 844 3834 884 3919
rect 844 3632 884 3641
rect 844 3137 884 3592
rect 843 3128 885 3137
rect 843 3088 844 3128
rect 884 3088 885 3128
rect 843 3079 885 3088
rect 940 2465 980 10219
rect 1036 3557 1076 12202
rect 1132 11621 1172 12412
rect 1227 12368 1269 12377
rect 1227 12328 1228 12368
rect 1268 12328 1269 12368
rect 1227 12319 1269 12328
rect 1228 12234 1268 12319
rect 1227 11780 1269 11789
rect 1227 11740 1228 11780
rect 1268 11740 1269 11780
rect 1227 11731 1269 11740
rect 1131 11612 1173 11621
rect 1131 11572 1132 11612
rect 1172 11572 1173 11612
rect 1131 11563 1173 11572
rect 1131 10940 1173 10949
rect 1131 10900 1132 10940
rect 1172 10900 1173 10940
rect 1131 10891 1173 10900
rect 1035 3548 1077 3557
rect 1035 3508 1036 3548
rect 1076 3508 1077 3548
rect 1035 3499 1077 3508
rect 1132 2885 1172 10891
rect 1228 4229 1268 11731
rect 1227 4220 1269 4229
rect 1227 4180 1228 4220
rect 1268 4180 1269 4220
rect 1227 4171 1269 4180
rect 1324 3725 1364 25087
rect 2091 20852 2133 20861
rect 2091 20812 2092 20852
rect 2132 20812 2133 20852
rect 2091 20803 2133 20812
rect 1611 20768 1653 20777
rect 1611 20728 1612 20768
rect 1652 20728 1653 20768
rect 1611 20719 1653 20728
rect 2092 20768 2132 20803
rect 1612 20096 1652 20719
rect 2092 20717 2132 20728
rect 2380 20768 2420 20777
rect 1612 20047 1652 20056
rect 2283 20096 2325 20105
rect 2283 20056 2284 20096
rect 2324 20056 2325 20096
rect 2283 20047 2325 20056
rect 1995 19592 2037 19601
rect 1995 19552 1996 19592
rect 2036 19552 2037 19592
rect 1995 19543 2037 19552
rect 1612 19256 1652 19265
rect 1900 19256 1940 19265
rect 1612 18677 1652 19216
rect 1804 19216 1900 19256
rect 1611 18668 1653 18677
rect 1611 18628 1612 18668
rect 1652 18628 1653 18668
rect 1611 18619 1653 18628
rect 1612 18089 1652 18619
rect 1611 18080 1653 18089
rect 1611 18040 1612 18080
rect 1652 18040 1653 18080
rect 1611 18031 1653 18040
rect 1804 17921 1844 19216
rect 1900 19207 1940 19216
rect 1996 19256 2036 19543
rect 2284 19508 2324 20047
rect 2284 19459 2324 19468
rect 2380 19265 2420 20728
rect 2475 20684 2517 20693
rect 2475 20644 2476 20684
rect 2516 20644 2517 20684
rect 2475 20635 2517 20644
rect 2476 20550 2516 20635
rect 2475 20096 2517 20105
rect 2475 20056 2476 20096
rect 2516 20056 2517 20096
rect 2475 20047 2517 20056
rect 2476 19962 2516 20047
rect 2475 19340 2517 19349
rect 2475 19300 2476 19340
rect 2516 19300 2517 19340
rect 2475 19291 2517 19300
rect 1996 19207 2036 19216
rect 2379 19256 2421 19265
rect 2379 19216 2380 19256
rect 2420 19216 2421 19256
rect 2379 19207 2421 19216
rect 2476 19206 2516 19291
rect 1900 18628 2516 18668
rect 1900 18500 1940 18628
rect 1900 18451 1940 18460
rect 2283 18500 2325 18509
rect 2283 18460 2284 18500
rect 2324 18460 2420 18500
rect 2283 18451 2325 18460
rect 2091 18416 2133 18425
rect 2091 18376 2092 18416
rect 2132 18376 2133 18416
rect 2091 18367 2133 18376
rect 1516 17912 1556 17921
rect 1803 17912 1845 17921
rect 1556 17872 1748 17912
rect 1516 17863 1556 17872
rect 1708 17744 1748 17872
rect 1803 17872 1804 17912
rect 1844 17872 1845 17912
rect 1803 17863 1845 17872
rect 1708 17695 1748 17704
rect 2092 17744 2132 18367
rect 2284 18366 2324 18451
rect 2283 18248 2325 18257
rect 2283 18208 2284 18248
rect 2324 18208 2325 18248
rect 2283 18199 2325 18208
rect 1996 16232 2036 16241
rect 2092 16232 2132 17704
rect 2036 16192 2132 16232
rect 1612 16148 1652 16157
rect 1516 15560 1556 15569
rect 1516 14729 1556 15520
rect 1612 15401 1652 16108
rect 1899 16064 1941 16073
rect 1899 16024 1900 16064
rect 1940 16024 1941 16064
rect 1899 16015 1941 16024
rect 1804 15560 1844 15569
rect 1611 15392 1653 15401
rect 1611 15352 1612 15392
rect 1652 15352 1653 15392
rect 1611 15343 1653 15352
rect 1804 14897 1844 15520
rect 1900 15560 1940 16015
rect 1900 15511 1940 15520
rect 1803 14888 1845 14897
rect 1803 14848 1804 14888
rect 1844 14848 1845 14888
rect 1803 14839 1845 14848
rect 1515 14720 1557 14729
rect 1515 14680 1516 14720
rect 1556 14680 1557 14720
rect 1515 14671 1557 14680
rect 1516 14048 1556 14671
rect 1516 12536 1556 14008
rect 1612 14636 1652 14645
rect 1612 13889 1652 14596
rect 1804 14300 1844 14839
rect 1996 14720 2036 16192
rect 2187 15392 2229 15401
rect 2187 15352 2188 15392
rect 2228 15352 2229 15392
rect 2187 15343 2229 15352
rect 2188 15258 2228 15343
rect 1996 14393 2036 14680
rect 1995 14384 2037 14393
rect 1995 14344 1996 14384
rect 2036 14344 2037 14384
rect 1995 14335 2037 14344
rect 1804 14260 1940 14300
rect 1804 14048 1844 14057
rect 1611 13880 1653 13889
rect 1611 13840 1612 13880
rect 1652 13840 1653 13880
rect 1611 13831 1653 13840
rect 1804 12956 1844 14008
rect 1900 14048 1940 14260
rect 1900 13999 1940 14008
rect 2187 13880 2229 13889
rect 2187 13840 2188 13880
rect 2228 13840 2229 13880
rect 2187 13831 2229 13840
rect 2188 13746 2228 13831
rect 2091 13208 2133 13217
rect 2091 13168 2092 13208
rect 2132 13168 2133 13208
rect 2091 13159 2133 13168
rect 2092 13074 2132 13159
rect 1804 12916 1940 12956
rect 1804 12536 1844 12545
rect 1556 12496 1748 12536
rect 1516 12487 1556 12496
rect 1708 11024 1748 12496
rect 1804 11705 1844 12496
rect 1900 12536 1940 12916
rect 2187 12872 2229 12881
rect 2187 12832 2188 12872
rect 2228 12832 2229 12872
rect 2187 12823 2229 12832
rect 2188 12746 2228 12823
rect 2188 12697 2228 12706
rect 1900 12293 1940 12496
rect 2284 12452 2324 18199
rect 2092 12412 2324 12452
rect 1899 12284 1941 12293
rect 1899 12244 1900 12284
rect 1940 12244 1941 12284
rect 1899 12235 1941 12244
rect 2092 12116 2132 12412
rect 2380 12242 2420 18460
rect 2476 18332 2516 18628
rect 2476 17165 2516 18292
rect 2572 17300 2612 35839
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 4971 34376 5013 34385
rect 4971 34336 4972 34376
rect 5012 34336 5013 34376
rect 4971 34327 5013 34336
rect 4779 34208 4821 34217
rect 4779 34168 4780 34208
rect 4820 34168 4821 34208
rect 4779 34159 4821 34168
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4395 32108 4437 32117
rect 4395 32068 4396 32108
rect 4436 32068 4437 32108
rect 4395 32059 4437 32068
rect 3819 31940 3861 31949
rect 3819 31900 3820 31940
rect 3860 31900 3861 31940
rect 3819 31891 3861 31900
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 2667 31688 2709 31697
rect 2667 31648 2668 31688
rect 2708 31648 2709 31688
rect 2667 31639 2709 31648
rect 2668 19349 2708 31639
rect 3820 31352 3860 31891
rect 4396 31781 4436 32059
rect 4587 31940 4629 31949
rect 4587 31900 4588 31940
rect 4628 31900 4629 31940
rect 4587 31891 4629 31900
rect 4588 31806 4628 31891
rect 4395 31772 4437 31781
rect 4395 31732 4396 31772
rect 4436 31732 4437 31772
rect 4395 31723 4437 31732
rect 3436 31268 3476 31277
rect 3436 30521 3476 31228
rect 3435 30512 3477 30521
rect 3435 30472 3436 30512
rect 3476 30472 3477 30512
rect 3435 30463 3477 30472
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3435 27656 3477 27665
rect 3435 27616 3436 27656
rect 3476 27616 3477 27656
rect 3435 27607 3477 27616
rect 3820 27656 3860 31312
rect 4684 31352 4724 31361
rect 4780 31352 4820 34159
rect 4972 32192 5012 34327
rect 5259 34040 5301 34049
rect 5259 34000 5260 34040
rect 5300 34000 5301 34040
rect 5259 33991 5301 34000
rect 4972 32143 5012 32152
rect 5164 31940 5204 31949
rect 5068 31900 5164 31940
rect 4724 31312 4820 31352
rect 4875 31352 4917 31361
rect 4875 31312 4876 31352
rect 4916 31312 4917 31352
rect 4684 31303 4724 31312
rect 4875 31303 4917 31312
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 4491 30764 4533 30773
rect 4491 30724 4492 30764
rect 4532 30724 4533 30764
rect 4491 30715 4533 30724
rect 4876 30764 4916 31303
rect 4876 30715 4916 30724
rect 4492 30680 4532 30715
rect 4492 29672 4532 30640
rect 4779 30680 4821 30689
rect 4779 30640 4780 30680
rect 4820 30640 4821 30680
rect 4779 30631 4821 30640
rect 4780 30546 4820 30631
rect 4875 30596 4917 30605
rect 4875 30556 4876 30596
rect 4916 30556 4917 30596
rect 4875 30547 4917 30556
rect 4204 29632 4532 29672
rect 4204 29336 4244 29632
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 4204 29296 4340 29336
rect 4300 28160 4340 29296
rect 4779 28328 4821 28337
rect 4779 28288 4780 28328
rect 4820 28288 4821 28328
rect 4779 28279 4821 28288
rect 4204 28120 4340 28160
rect 4204 27824 4244 28120
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 4204 27784 4532 27824
rect 3436 27522 3476 27607
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3820 25304 3860 27616
rect 4492 26816 4532 27784
rect 4300 26776 4492 26816
rect 4300 26648 4340 26776
rect 4492 26767 4532 26776
rect 4684 27656 4724 27665
rect 4780 27656 4820 28279
rect 4724 27616 4820 27656
rect 4204 26608 4340 26648
rect 4684 26648 4724 27616
rect 4876 27572 4916 30547
rect 5068 28337 5108 31900
rect 5164 31891 5204 31900
rect 5260 30773 5300 33991
rect 5452 32948 5492 36175
rect 7084 36065 7124 36679
rect 17836 36594 17876 36679
rect 7083 36056 7125 36065
rect 7083 36016 7084 36056
rect 7124 36016 7125 36056
rect 7083 36007 7125 36016
rect 14860 36056 14900 36065
rect 6411 35888 6453 35897
rect 6411 35848 6412 35888
rect 6452 35848 6453 35888
rect 6411 35839 6453 35848
rect 5547 33872 5589 33881
rect 5547 33832 5548 33872
rect 5588 33832 5589 33872
rect 5547 33823 5589 33832
rect 5452 32899 5492 32908
rect 5259 30764 5301 30773
rect 5259 30724 5260 30764
rect 5300 30724 5301 30764
rect 5259 30715 5301 30724
rect 5355 30680 5397 30689
rect 5355 30640 5356 30680
rect 5396 30640 5397 30680
rect 5355 30631 5397 30640
rect 5163 30512 5205 30521
rect 5163 30472 5164 30512
rect 5204 30472 5205 30512
rect 5163 30463 5205 30472
rect 5164 30378 5204 30463
rect 5067 28328 5109 28337
rect 5067 28288 5068 28328
rect 5108 28288 5109 28328
rect 5067 28279 5109 28288
rect 4971 28076 5013 28085
rect 4971 28036 4972 28076
rect 5012 28036 5013 28076
rect 4971 28027 5013 28036
rect 4780 27532 4916 27572
rect 4780 26816 4820 27532
rect 4780 26767 4820 26776
rect 4875 26732 4917 26741
rect 4875 26692 4876 26732
rect 4916 26692 4917 26732
rect 4875 26683 4917 26692
rect 4684 26608 4820 26648
rect 4204 26312 4244 26608
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 4204 26272 4340 26312
rect 3435 25220 3477 25229
rect 3435 25180 3436 25220
rect 3476 25180 3477 25220
rect 3435 25171 3477 25180
rect 3436 25086 3476 25171
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 3436 23129 3476 23214
rect 3435 23120 3477 23129
rect 3435 23080 3436 23120
rect 3476 23080 3477 23120
rect 3435 23071 3477 23080
rect 3820 23120 3860 25264
rect 4300 25136 4340 26272
rect 4684 25304 4724 25313
rect 4780 25304 4820 26608
rect 4876 26598 4916 26683
rect 4724 25264 4916 25304
rect 4684 25255 4724 25264
rect 4204 25096 4340 25136
rect 4204 24800 4244 25096
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 4204 24760 4436 24800
rect 4300 23624 4340 24760
rect 4396 24632 4436 24760
rect 4779 24716 4821 24725
rect 4779 24676 4780 24716
rect 4820 24676 4821 24716
rect 4779 24667 4821 24676
rect 4396 24583 4436 24592
rect 4684 24632 4724 24641
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 3723 22364 3765 22373
rect 3723 22324 3724 22364
rect 3764 22324 3765 22364
rect 3723 22315 3765 22324
rect 3724 22280 3764 22315
rect 3724 22229 3764 22240
rect 3436 21608 3476 21617
rect 3820 21608 3860 23080
rect 4204 23584 4340 23624
rect 4684 23624 4724 24592
rect 4780 24582 4820 24667
rect 4684 23584 4820 23624
rect 4204 22373 4244 23584
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 4780 23288 4820 23584
rect 4588 23248 4820 23288
rect 4395 23120 4437 23129
rect 4395 23080 4396 23120
rect 4436 23080 4437 23120
rect 4395 23071 4437 23080
rect 4396 22532 4436 23071
rect 4396 22483 4436 22492
rect 3915 22364 3957 22373
rect 3915 22324 3916 22364
rect 3956 22324 3957 22364
rect 3915 22315 3957 22324
rect 4203 22364 4245 22373
rect 4203 22324 4204 22364
rect 4244 22324 4245 22364
rect 4203 22315 4245 22324
rect 3476 21568 3572 21608
rect 3436 21559 3476 21568
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 2764 20936 2804 20945
rect 2804 20896 2996 20936
rect 2764 20887 2804 20896
rect 2956 20768 2996 20896
rect 2956 20719 2996 20728
rect 3339 20768 3381 20777
rect 3339 20728 3340 20768
rect 3380 20728 3381 20768
rect 3339 20719 3381 20728
rect 3340 20634 3380 20719
rect 3532 19937 3572 21568
rect 3820 20777 3860 21568
rect 3916 20861 3956 22315
rect 4588 22289 4628 23248
rect 4684 23120 4724 23129
rect 4724 23080 4820 23120
rect 4684 23071 4724 23080
rect 4780 23060 4820 23080
rect 4876 23060 4916 25264
rect 4780 23020 4916 23060
rect 4012 22280 4052 22289
rect 3915 20852 3957 20861
rect 3915 20812 3916 20852
rect 3956 20812 3957 20852
rect 3915 20803 3957 20812
rect 3819 20768 3861 20777
rect 3819 20728 3820 20768
rect 3860 20728 3861 20768
rect 3819 20719 3861 20728
rect 3916 20096 3956 20803
rect 4012 20693 4052 22240
rect 4107 22280 4149 22289
rect 4107 22240 4108 22280
rect 4148 22240 4149 22280
rect 4107 22231 4149 22240
rect 4587 22280 4629 22289
rect 4587 22240 4588 22280
rect 4628 22240 4629 22280
rect 4587 22231 4629 22240
rect 4108 22146 4148 22231
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 4684 21608 4724 21617
rect 4780 21608 4820 23020
rect 4204 21568 4684 21608
rect 4724 21568 4820 21608
rect 4204 20768 4244 21568
rect 4684 21559 4724 21568
rect 4779 20852 4821 20861
rect 4779 20812 4780 20852
rect 4820 20812 4821 20852
rect 4779 20803 4821 20812
rect 4108 20728 4204 20768
rect 4011 20684 4053 20693
rect 4011 20644 4012 20684
rect 4052 20644 4053 20684
rect 4011 20635 4053 20644
rect 4108 20105 4148 20728
rect 4204 20719 4244 20728
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4299 20180 4341 20189
rect 4299 20140 4300 20180
rect 4340 20140 4341 20180
rect 4299 20131 4341 20140
rect 3916 20047 3956 20056
rect 4107 20096 4149 20105
rect 4107 20056 4108 20096
rect 4148 20056 4149 20096
rect 4107 20047 4149 20056
rect 4204 20096 4244 20105
rect 3531 19928 3573 19937
rect 3531 19888 3532 19928
rect 3572 19888 3573 19928
rect 3531 19879 3573 19888
rect 3628 19844 3668 19853
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3628 19601 3668 19804
rect 4204 19601 4244 20056
rect 4300 20046 4340 20131
rect 4587 19928 4629 19937
rect 4587 19888 4588 19928
rect 4628 19888 4629 19928
rect 4587 19879 4629 19888
rect 4588 19794 4628 19879
rect 3627 19592 3669 19601
rect 3627 19552 3628 19592
rect 3668 19552 3669 19592
rect 3627 19543 3669 19552
rect 4203 19592 4245 19601
rect 4203 19552 4204 19592
rect 4244 19552 4245 19592
rect 4203 19543 4245 19552
rect 3531 19508 3573 19517
rect 3531 19468 3532 19508
rect 3572 19468 3573 19508
rect 3531 19459 3573 19468
rect 3435 19424 3477 19433
rect 3435 19384 3436 19424
rect 3476 19384 3477 19424
rect 3435 19375 3477 19384
rect 2667 19340 2709 19349
rect 2667 19300 2668 19340
rect 2708 19300 2804 19340
rect 2667 19291 2709 19300
rect 2668 19088 2708 19097
rect 2668 18509 2708 19048
rect 2667 18500 2709 18509
rect 2667 18460 2668 18500
rect 2708 18460 2709 18500
rect 2667 18451 2709 18460
rect 2764 18257 2804 19300
rect 3436 18668 3476 19375
rect 3436 18619 3476 18628
rect 3532 19340 3572 19459
rect 4683 19424 4725 19433
rect 2763 18248 2805 18257
rect 2763 18208 2764 18248
rect 2804 18208 2805 18248
rect 2763 18199 2805 18208
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 2956 17744 2996 17753
rect 2956 17300 2996 17704
rect 2572 17260 2708 17300
rect 2475 17156 2517 17165
rect 2475 17116 2476 17156
rect 2516 17116 2517 17156
rect 2475 17107 2517 17116
rect 2284 12202 2420 12242
rect 2092 12076 2228 12116
rect 1803 11696 1845 11705
rect 1803 11656 1804 11696
rect 1844 11656 1845 11696
rect 1803 11647 1845 11656
rect 2091 11696 2133 11705
rect 2091 11656 2092 11696
rect 2132 11656 2133 11696
rect 2091 11647 2133 11656
rect 1899 11612 1941 11621
rect 1899 11572 1900 11612
rect 1940 11572 1941 11612
rect 1899 11563 1941 11572
rect 1708 10975 1748 10984
rect 1900 9857 1940 11563
rect 2092 11108 2132 11647
rect 2092 11059 2132 11068
rect 1995 11024 2037 11033
rect 1995 10984 1996 11024
rect 2036 10984 2037 11024
rect 1995 10975 2037 10984
rect 1996 10890 2036 10975
rect 2188 10697 2228 12076
rect 2187 10688 2229 10697
rect 2187 10648 2188 10688
rect 2228 10648 2229 10688
rect 2187 10639 2229 10648
rect 1899 9848 1941 9857
rect 1899 9808 1900 9848
rect 1940 9808 1941 9848
rect 1899 9799 1941 9808
rect 2284 6665 2324 12202
rect 2380 11234 2420 11243
rect 2380 11108 2420 11194
rect 2572 11108 2612 11117
rect 2380 11068 2572 11108
rect 2572 11059 2612 11068
rect 2475 10688 2517 10697
rect 2475 10648 2476 10688
rect 2516 10648 2517 10688
rect 2475 10639 2517 10648
rect 2379 9848 2421 9857
rect 2379 9808 2380 9848
rect 2420 9808 2421 9848
rect 2379 9799 2421 9808
rect 2283 6656 2325 6665
rect 2283 6616 2284 6656
rect 2324 6616 2325 6656
rect 2283 6607 2325 6616
rect 1323 3716 1365 3725
rect 1323 3676 1324 3716
rect 1364 3676 1365 3716
rect 1323 3667 1365 3676
rect 1131 2876 1173 2885
rect 1131 2836 1132 2876
rect 1172 2836 1173 2876
rect 1131 2827 1173 2836
rect 2380 2801 2420 9799
rect 2476 5405 2516 10639
rect 2668 7220 2708 17260
rect 2860 17260 2996 17300
rect 3532 17300 3572 19300
rect 3916 19384 4148 19424
rect 3724 19088 3764 19097
rect 3724 18677 3764 19048
rect 3723 18668 3765 18677
rect 3723 18628 3724 18668
rect 3764 18628 3765 18668
rect 3723 18619 3765 18628
rect 3820 18584 3860 18593
rect 3820 18425 3860 18544
rect 3819 18416 3861 18425
rect 3819 18376 3820 18416
rect 3860 18376 3861 18416
rect 3819 18367 3861 18376
rect 3532 17260 3764 17300
rect 2860 16232 2900 17260
rect 3435 17072 3477 17081
rect 3435 17032 3436 17072
rect 3476 17032 3477 17072
rect 3435 17023 3477 17032
rect 3436 16938 3476 17023
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 2860 15989 2900 16192
rect 2859 15980 2901 15989
rect 2859 15940 2860 15980
rect 2900 15940 2901 15980
rect 2859 15931 2901 15940
rect 2860 14720 2900 15931
rect 3435 15560 3477 15569
rect 3435 15520 3436 15560
rect 3476 15520 3477 15560
rect 3435 15511 3477 15520
rect 3436 15426 3476 15511
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 2860 14671 2900 14680
rect 3627 14720 3669 14729
rect 3627 14680 3628 14720
rect 3668 14680 3669 14720
rect 3627 14671 3669 14680
rect 3531 14384 3573 14393
rect 3531 14344 3532 14384
rect 3572 14344 3573 14384
rect 3531 14335 3573 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 2955 13376 2997 13385
rect 2955 13336 2956 13376
rect 2996 13336 2997 13376
rect 2955 13327 2997 13336
rect 2763 12452 2805 12461
rect 2763 12412 2764 12452
rect 2804 12412 2805 12452
rect 2763 12403 2805 12412
rect 2572 7180 2708 7220
rect 2572 6917 2612 7180
rect 2571 6908 2613 6917
rect 2571 6868 2572 6908
rect 2612 6868 2613 6908
rect 2571 6859 2613 6868
rect 2764 6497 2804 12403
rect 2956 11024 2996 13327
rect 3435 13292 3477 13301
rect 3435 13252 3436 13292
rect 3476 13252 3477 13292
rect 3435 13243 3477 13252
rect 3436 13208 3476 13243
rect 3436 13157 3476 13168
rect 3244 13040 3284 13049
rect 3244 12293 3284 13000
rect 3435 12536 3477 12545
rect 3435 12496 3436 12536
rect 3476 12496 3477 12536
rect 3435 12487 3477 12496
rect 3436 12402 3476 12487
rect 3243 12284 3285 12293
rect 3243 12244 3244 12284
rect 3284 12244 3285 12284
rect 3243 12235 3285 12244
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 2956 10975 2996 10984
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3435 10100 3477 10109
rect 3435 10060 3436 10100
rect 3476 10060 3477 10100
rect 3435 10051 3477 10060
rect 3436 9966 3476 10051
rect 3532 10025 3572 14335
rect 3628 14048 3668 14671
rect 3628 11621 3668 14008
rect 3627 11612 3669 11621
rect 3627 11572 3628 11612
rect 3668 11572 3669 11612
rect 3627 11563 3669 11572
rect 3627 11024 3669 11033
rect 3627 10984 3628 11024
rect 3668 10984 3669 11024
rect 3627 10975 3669 10984
rect 3628 10277 3668 10975
rect 3627 10268 3669 10277
rect 3627 10228 3628 10268
rect 3668 10228 3669 10268
rect 3627 10219 3669 10228
rect 3531 10016 3573 10025
rect 3531 9976 3532 10016
rect 3572 9976 3573 10016
rect 3531 9967 3573 9976
rect 3628 9521 3668 10219
rect 3724 9605 3764 17260
rect 3820 17165 3860 17196
rect 3819 17156 3861 17165
rect 3819 17116 3820 17156
rect 3860 17116 3861 17156
rect 3819 17107 3861 17116
rect 3820 17072 3860 17107
rect 3820 15560 3860 17032
rect 3820 14216 3860 15520
rect 3916 14393 3956 19384
rect 4012 19256 4052 19265
rect 4108 19256 4148 19384
rect 4683 19384 4684 19424
rect 4724 19384 4725 19424
rect 4683 19375 4725 19384
rect 4684 19290 4724 19375
rect 4300 19256 4340 19265
rect 4108 19216 4300 19256
rect 4012 18005 4052 19216
rect 4300 19207 4340 19216
rect 4395 19256 4437 19265
rect 4395 19216 4396 19256
rect 4436 19216 4437 19256
rect 4395 19207 4437 19216
rect 4396 19122 4436 19207
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4299 18668 4341 18677
rect 4299 18628 4300 18668
rect 4340 18628 4341 18668
rect 4299 18619 4341 18628
rect 4011 17996 4053 18005
rect 4011 17956 4012 17996
rect 4052 17956 4053 17996
rect 4011 17947 4053 17956
rect 4012 17300 4052 17947
rect 4107 17912 4149 17921
rect 4107 17872 4108 17912
rect 4148 17872 4149 17912
rect 4107 17863 4149 17872
rect 4108 17778 4148 17863
rect 4300 17828 4340 18619
rect 4684 18584 4724 18593
rect 4780 18584 4820 20803
rect 4875 19340 4917 19349
rect 4875 19300 4876 19340
rect 4916 19300 4917 19340
rect 4875 19291 4917 19300
rect 4876 19206 4916 19291
rect 4724 18544 4820 18584
rect 4684 18535 4724 18544
rect 4491 17996 4533 18005
rect 4491 17956 4492 17996
rect 4532 17956 4533 17996
rect 4491 17947 4533 17956
rect 4492 17862 4532 17947
rect 4204 17788 4300 17828
rect 4204 17300 4244 17788
rect 4300 17779 4340 17788
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4012 17260 4148 17300
rect 4204 17260 4340 17300
rect 4011 16904 4053 16913
rect 4011 16864 4012 16904
rect 4052 16864 4053 16904
rect 4011 16855 4053 16864
rect 4012 16484 4052 16855
rect 4012 16435 4052 16444
rect 4011 16064 4053 16073
rect 4011 16024 4012 16064
rect 4052 16024 4053 16064
rect 4011 16015 4053 16024
rect 4012 15930 4052 16015
rect 4011 14888 4053 14897
rect 4011 14848 4012 14888
rect 4052 14848 4053 14888
rect 4011 14839 4053 14848
rect 4012 14754 4052 14839
rect 4108 14729 4148 17260
rect 4300 16232 4340 17260
rect 4684 17072 4724 17081
rect 4780 17072 4820 18544
rect 4972 17300 5012 28027
rect 5163 27656 5205 27665
rect 5163 27616 5164 27656
rect 5204 27616 5205 27656
rect 5163 27607 5205 27616
rect 5164 27068 5204 27607
rect 5259 27404 5301 27413
rect 5259 27364 5260 27404
rect 5300 27364 5301 27404
rect 5259 27355 5301 27364
rect 5164 27019 5204 27028
rect 5163 26732 5205 26741
rect 5260 26732 5300 27355
rect 5163 26692 5164 26732
rect 5204 26692 5300 26732
rect 5163 26683 5205 26692
rect 5067 25220 5109 25229
rect 5067 25180 5068 25220
rect 5108 25180 5109 25220
rect 5067 25171 5109 25180
rect 5068 24842 5108 25171
rect 5068 24793 5108 24802
rect 5067 19508 5109 19517
rect 5067 19468 5068 19508
rect 5108 19468 5109 19508
rect 5067 19459 5109 19468
rect 5068 19374 5108 19459
rect 4724 17032 4820 17072
rect 4684 17023 4724 17032
rect 4683 16736 4725 16745
rect 4683 16696 4684 16736
rect 4724 16696 4725 16736
rect 4683 16687 4725 16696
rect 4300 16183 4340 16192
rect 4587 16232 4629 16241
rect 4587 16192 4588 16232
rect 4628 16192 4629 16232
rect 4587 16183 4629 16192
rect 4684 16232 4724 16687
rect 4684 16183 4724 16192
rect 4588 16098 4628 16183
rect 4780 15989 4820 17032
rect 4876 17260 5012 17300
rect 4779 15980 4821 15989
rect 4779 15940 4780 15980
rect 4820 15940 4821 15980
rect 4779 15931 4821 15940
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4684 15560 4724 15569
rect 4780 15560 4820 15931
rect 4724 15520 4820 15560
rect 4684 15511 4724 15520
rect 4684 14729 4724 14814
rect 4107 14720 4149 14729
rect 4300 14720 4340 14729
rect 4107 14680 4108 14720
rect 4148 14680 4300 14720
rect 4107 14671 4149 14680
rect 4300 14671 4340 14680
rect 4588 14720 4628 14729
rect 4108 14586 4148 14671
rect 4588 14552 4628 14680
rect 4683 14720 4725 14729
rect 4683 14680 4684 14720
rect 4724 14680 4725 14720
rect 4683 14671 4725 14680
rect 4588 14512 4820 14552
rect 3915 14384 3957 14393
rect 3915 14344 3916 14384
rect 3956 14344 3957 14384
rect 3915 14335 3957 14344
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3820 14176 4148 14216
rect 3916 14048 3956 14057
rect 3819 13376 3861 13385
rect 3819 13336 3820 13376
rect 3860 13336 3861 13376
rect 3819 13327 3861 13336
rect 3820 13208 3860 13327
rect 3820 12536 3860 13168
rect 3820 12487 3860 12496
rect 3916 11873 3956 14008
rect 4011 14048 4053 14057
rect 4011 14008 4012 14048
rect 4052 14008 4053 14048
rect 4011 13999 4053 14008
rect 4012 13914 4052 13999
rect 4011 11948 4053 11957
rect 4011 11908 4012 11948
rect 4052 11908 4053 11948
rect 4011 11899 4053 11908
rect 3915 11864 3957 11873
rect 3915 11824 3916 11864
rect 3956 11824 3957 11864
rect 3915 11815 3957 11824
rect 3916 11696 3956 11707
rect 3916 11621 3956 11656
rect 3915 11612 3957 11621
rect 3915 11572 3916 11612
rect 3956 11572 3957 11612
rect 3915 11563 3957 11572
rect 3819 11024 3861 11033
rect 3819 10984 3820 11024
rect 3860 10984 3861 11024
rect 3819 10975 3861 10984
rect 3820 10890 3860 10975
rect 3819 10772 3861 10781
rect 3819 10732 3820 10772
rect 3860 10732 3861 10772
rect 3819 10723 3861 10732
rect 3820 10184 3860 10723
rect 4012 10604 4052 11899
rect 4108 10781 4148 14176
rect 4780 14057 4820 14512
rect 4779 14048 4821 14057
rect 4779 14008 4780 14048
rect 4820 14008 4821 14048
rect 4779 13999 4821 14008
rect 4300 13796 4340 13805
rect 4300 13301 4340 13756
rect 4299 13292 4341 13301
rect 4299 13252 4300 13292
rect 4340 13252 4341 13292
rect 4299 13243 4341 13252
rect 4683 13208 4725 13217
rect 4876 13208 4916 17260
rect 4971 17072 5013 17081
rect 4971 17032 4972 17072
rect 5012 17032 5013 17072
rect 4971 17023 5013 17032
rect 4972 16484 5012 17023
rect 4972 16435 5012 16444
rect 5067 16232 5109 16241
rect 5067 16192 5068 16232
rect 5108 16192 5109 16232
rect 5067 16183 5109 16192
rect 4971 15560 5013 15569
rect 4971 15520 4972 15560
rect 5012 15520 5013 15560
rect 4971 15511 5013 15520
rect 4972 14972 5012 15511
rect 4972 14923 5012 14932
rect 5068 14729 5108 16183
rect 5067 14720 5109 14729
rect 5067 14680 5068 14720
rect 5108 14680 5109 14720
rect 5067 14671 5109 14680
rect 4683 13168 4684 13208
rect 4724 13168 4916 13208
rect 4683 13159 4725 13168
rect 4684 13074 4724 13159
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4203 12788 4245 12797
rect 4203 12748 4204 12788
rect 4244 12748 4245 12788
rect 4203 12739 4245 12748
rect 4204 11696 4244 12739
rect 4587 12536 4629 12545
rect 4587 12496 4588 12536
rect 4628 12496 4629 12536
rect 4587 12487 4629 12496
rect 4684 12536 4724 12545
rect 4780 12536 4820 13168
rect 4724 12496 4820 12536
rect 4684 12487 4724 12496
rect 4588 11948 4628 12487
rect 4588 11899 4628 11908
rect 4299 11864 4341 11873
rect 4299 11824 4300 11864
rect 4340 11824 4341 11864
rect 4299 11815 4341 11824
rect 4204 11647 4244 11656
rect 4300 11696 4340 11815
rect 4300 11647 4340 11656
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4780 11033 4820 12496
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 4971 12487 5013 12496
rect 4972 11705 5012 12487
rect 5164 11957 5204 26683
rect 5356 21533 5396 30631
rect 5548 28085 5588 33823
rect 5643 33116 5685 33125
rect 5643 33076 5644 33116
rect 5684 33076 5685 33116
rect 5643 33067 5685 33076
rect 5644 32982 5684 33067
rect 5644 32696 5684 32705
rect 5644 32117 5684 32656
rect 5643 32108 5685 32117
rect 5643 32068 5644 32108
rect 5684 32068 5685 32108
rect 5643 32059 5685 32068
rect 5739 31688 5781 31697
rect 5739 31648 5740 31688
rect 5780 31648 5781 31688
rect 5739 31639 5781 31648
rect 5740 30605 5780 31639
rect 5931 31520 5973 31529
rect 5931 31480 5932 31520
rect 5972 31480 5973 31520
rect 5931 31471 5973 31480
rect 5836 31436 5876 31447
rect 5836 31361 5876 31396
rect 5835 31352 5877 31361
rect 5835 31312 5836 31352
rect 5876 31312 5877 31352
rect 5835 31303 5877 31312
rect 5739 30596 5781 30605
rect 5739 30556 5740 30596
rect 5780 30556 5781 30596
rect 5739 30547 5781 30556
rect 5547 28076 5589 28085
rect 5547 28036 5548 28076
rect 5588 28036 5589 28076
rect 5547 28027 5589 28036
rect 5835 27404 5877 27413
rect 5835 27364 5836 27404
rect 5876 27364 5877 27404
rect 5835 27355 5877 27364
rect 5836 27270 5876 27355
rect 5836 25556 5876 25565
rect 5932 25556 5972 31471
rect 6027 25976 6069 25985
rect 6027 25936 6028 25976
rect 6068 25936 6069 25976
rect 6027 25927 6069 25936
rect 5876 25516 5972 25556
rect 5836 25507 5876 25516
rect 5836 25136 5876 25145
rect 5836 24725 5876 25096
rect 5835 24716 5877 24725
rect 5835 24676 5836 24716
rect 5876 24676 5877 24716
rect 5835 24667 5877 24676
rect 5836 22868 5876 22877
rect 5876 22828 5972 22868
rect 5836 22819 5876 22828
rect 5932 22289 5972 22828
rect 5931 22280 5973 22289
rect 5931 22240 5932 22280
rect 5972 22240 5973 22280
rect 5931 22231 5973 22240
rect 5835 21944 5877 21953
rect 5835 21904 5836 21944
rect 5876 21904 5877 21944
rect 5835 21895 5877 21904
rect 5836 21533 5876 21895
rect 5355 21524 5397 21533
rect 5260 21484 5356 21524
rect 5396 21484 5397 21524
rect 5260 20189 5300 21484
rect 5355 21475 5397 21484
rect 5835 21524 5877 21533
rect 5835 21484 5836 21524
rect 5876 21484 5877 21524
rect 5835 21475 5877 21484
rect 5836 21390 5876 21475
rect 5932 20945 5972 22231
rect 5931 20936 5973 20945
rect 5931 20896 5932 20936
rect 5972 20896 5973 20936
rect 5931 20887 5973 20896
rect 5356 20693 5396 20724
rect 5355 20684 5397 20693
rect 5355 20644 5356 20684
rect 5396 20644 5397 20684
rect 5355 20635 5397 20644
rect 5356 20600 5396 20635
rect 5259 20180 5301 20189
rect 5259 20140 5260 20180
rect 5300 20140 5301 20180
rect 5259 20131 5301 20140
rect 5356 18929 5396 20560
rect 6028 19265 6068 25927
rect 6412 19349 6452 35839
rect 6411 19340 6453 19349
rect 6411 19300 6412 19340
rect 6452 19300 6453 19340
rect 6411 19291 6453 19300
rect 6027 19256 6069 19265
rect 6027 19216 6028 19256
rect 6068 19216 6069 19256
rect 6027 19207 6069 19216
rect 5355 18920 5397 18929
rect 5355 18880 5356 18920
rect 5396 18880 5397 18920
rect 5355 18871 5397 18880
rect 5836 18500 5876 18509
rect 6028 18500 6068 19207
rect 5876 18460 6068 18500
rect 5836 18451 5876 18460
rect 5836 16820 5876 16831
rect 5836 16745 5876 16780
rect 5835 16736 5877 16745
rect 5835 16696 5836 16736
rect 5876 16696 5877 16736
rect 5835 16687 5877 16696
rect 5835 16568 5877 16577
rect 5835 16528 5836 16568
rect 5876 16528 5877 16568
rect 5835 16519 5877 16528
rect 5836 16241 5876 16519
rect 5835 16232 5877 16241
rect 5835 16192 5836 16232
rect 5876 16192 5877 16232
rect 5835 16183 5877 16192
rect 5836 15728 5876 16183
rect 5836 15679 5876 15688
rect 5835 14048 5877 14057
rect 5835 14008 5836 14048
rect 5876 14008 5877 14048
rect 5835 13999 5877 14008
rect 5836 13460 5876 13999
rect 5836 13411 5876 13420
rect 5836 13040 5876 13049
rect 5739 12788 5781 12797
rect 5739 12748 5740 12788
rect 5780 12748 5781 12788
rect 5739 12739 5781 12748
rect 5163 11948 5205 11957
rect 5163 11908 5164 11948
rect 5204 11908 5205 11948
rect 5163 11899 5205 11908
rect 4971 11696 5013 11705
rect 4971 11656 4972 11696
rect 5012 11656 5013 11696
rect 4971 11647 5013 11656
rect 4972 11192 5012 11647
rect 4972 11143 5012 11152
rect 4779 11024 4821 11033
rect 4779 10984 4780 11024
rect 4820 10984 4821 11024
rect 4779 10975 4821 10984
rect 4107 10772 4149 10781
rect 4107 10732 4108 10772
rect 4148 10732 4149 10772
rect 4107 10723 4149 10732
rect 4012 10564 4148 10604
rect 3723 9596 3765 9605
rect 3723 9556 3724 9596
rect 3764 9556 3765 9596
rect 3723 9547 3765 9556
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3435 8000 3477 8009
rect 3435 7960 3436 8000
rect 3476 7960 3477 8000
rect 3435 7951 3477 7960
rect 3820 8000 3860 10144
rect 4011 9596 4053 9605
rect 4011 9556 4012 9596
rect 4052 9556 4053 9596
rect 4011 9547 4053 9556
rect 3820 7951 3860 7960
rect 4012 9512 4052 9547
rect 4108 9512 4148 10564
rect 4684 10184 4724 10193
rect 4780 10184 4820 10975
rect 4724 10144 4820 10184
rect 4684 10135 4724 10144
rect 4203 10100 4245 10109
rect 4203 10060 4204 10100
rect 4244 10060 4245 10100
rect 4203 10051 4245 10060
rect 4204 9680 4244 10051
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4204 9640 4724 9680
rect 4300 9512 4340 9521
rect 4108 9472 4300 9512
rect 3436 7866 3476 7951
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4012 7085 4052 9472
rect 4300 9463 4340 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4396 9378 4436 9463
rect 4684 9344 4724 9640
rect 4684 9295 4724 9304
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4684 8000 4724 8009
rect 4780 8000 4820 10144
rect 5740 8168 5780 12739
rect 5836 12713 5876 13000
rect 5835 12704 5877 12713
rect 5835 12664 5836 12704
rect 5876 12664 5877 12704
rect 5835 12655 5877 12664
rect 5836 12377 5876 12408
rect 5835 12368 5877 12377
rect 5835 12328 5836 12368
rect 5876 12328 5877 12368
rect 5835 12319 5877 12328
rect 5836 12284 5876 12319
rect 5836 11873 5876 12244
rect 5835 11864 5877 11873
rect 5835 11824 5836 11864
rect 5876 11824 5877 11864
rect 5835 11815 5877 11824
rect 5835 10268 5877 10277
rect 5835 10228 5836 10268
rect 5876 10228 5972 10268
rect 5835 10219 5877 10228
rect 5836 10134 5876 10219
rect 5836 8168 5876 8177
rect 5740 8128 5836 8168
rect 4724 7960 4820 8000
rect 5067 8000 5109 8009
rect 5067 7960 5068 8000
rect 5108 7960 5109 8000
rect 4684 7951 4724 7960
rect 5067 7951 5109 7960
rect 4779 7748 4821 7757
rect 4779 7708 4780 7748
rect 4820 7708 4821 7748
rect 4779 7699 4821 7708
rect 4396 7160 4436 7171
rect 4396 7085 4436 7120
rect 4683 7160 4725 7169
rect 4683 7120 4684 7160
rect 4724 7120 4725 7160
rect 4683 7111 4725 7120
rect 4780 7160 4820 7699
rect 5068 7412 5108 7951
rect 5740 7757 5780 8128
rect 5836 8119 5876 8128
rect 5739 7748 5781 7757
rect 5739 7708 5740 7748
rect 5780 7708 5781 7748
rect 5739 7699 5781 7708
rect 5068 7363 5108 7372
rect 4011 7076 4053 7085
rect 4011 7036 4012 7076
rect 4052 7036 4053 7076
rect 4011 7027 4053 7036
rect 4395 7076 4437 7085
rect 4395 7036 4396 7076
rect 4436 7036 4437 7076
rect 4395 7027 4437 7036
rect 4684 7026 4724 7111
rect 4780 7110 4820 7120
rect 5932 6833 5972 10228
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 5931 6824 5973 6833
rect 5931 6784 5932 6824
rect 5972 6784 5973 6824
rect 5931 6775 5973 6784
rect 6412 6581 6452 19291
rect 6411 6572 6453 6581
rect 6411 6532 6412 6572
rect 6452 6532 6453 6572
rect 6411 6523 6453 6532
rect 2763 6488 2805 6497
rect 2763 6448 2764 6488
rect 2804 6448 2805 6488
rect 2763 6439 2805 6448
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 2475 5396 2517 5405
rect 2475 5356 2476 5396
rect 2516 5356 2517 5396
rect 2475 5347 2517 5356
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 7084 5153 7124 36007
rect 13708 35972 13748 35983
rect 13708 35897 13748 35932
rect 13707 35888 13749 35897
rect 13707 35848 13708 35888
rect 13748 35848 13749 35888
rect 13707 35839 13749 35848
rect 14188 35888 14228 35897
rect 13900 35720 13940 35729
rect 13900 35384 13940 35680
rect 13612 35344 13940 35384
rect 13420 35216 13460 35225
rect 13612 35216 13652 35344
rect 14188 35225 14228 35848
rect 14476 35888 14516 35897
rect 14860 35888 14900 36016
rect 15244 35888 15284 35897
rect 14860 35848 15244 35888
rect 13460 35176 13652 35216
rect 13708 35216 13748 35225
rect 12267 35132 12309 35141
rect 12267 35092 12268 35132
rect 12308 35092 12309 35132
rect 12267 35083 12309 35092
rect 12459 35132 12501 35141
rect 12459 35092 12460 35132
rect 12500 35092 12501 35132
rect 12459 35083 12501 35092
rect 12268 34998 12308 35083
rect 12460 34964 12500 35083
rect 7371 34544 7413 34553
rect 7371 34504 7372 34544
rect 7412 34504 7413 34544
rect 7371 34495 7413 34504
rect 11596 34544 11636 34553
rect 11636 34504 11828 34544
rect 11596 34495 11636 34504
rect 7372 34385 7412 34495
rect 7371 34376 7413 34385
rect 7371 34336 7372 34376
rect 7412 34336 7413 34376
rect 7371 34327 7413 34336
rect 10924 34376 10964 34385
rect 7372 34242 7412 34327
rect 7756 34208 7796 34217
rect 7756 20861 7796 34168
rect 10924 34049 10964 34336
rect 11212 34376 11252 34385
rect 10923 34040 10965 34049
rect 10923 34000 10924 34040
rect 10964 34000 10965 34040
rect 10923 33991 10965 34000
rect 8235 33956 8277 33965
rect 8235 33916 8236 33956
rect 8276 33916 8277 33956
rect 8235 33907 8277 33916
rect 7851 31604 7893 31613
rect 7851 31564 7852 31604
rect 7892 31564 7893 31604
rect 7851 31555 7893 31564
rect 7755 20852 7797 20861
rect 7755 20812 7756 20852
rect 7796 20812 7797 20852
rect 7755 20803 7797 20812
rect 7755 16736 7797 16745
rect 7755 16696 7756 16736
rect 7796 16696 7797 16736
rect 7755 16687 7797 16696
rect 7756 16409 7796 16687
rect 7755 16400 7797 16409
rect 7755 16360 7756 16400
rect 7796 16360 7797 16400
rect 7755 16351 7797 16360
rect 7852 5825 7892 31555
rect 7947 16400 7989 16409
rect 7947 16360 7948 16400
rect 7988 16360 7989 16400
rect 7947 16351 7989 16360
rect 7948 7001 7988 16351
rect 7947 6992 7989 7001
rect 7947 6952 7948 6992
rect 7988 6952 7989 6992
rect 7947 6943 7989 6952
rect 7851 5816 7893 5825
rect 7851 5776 7852 5816
rect 7892 5776 7893 5816
rect 7851 5767 7893 5776
rect 7083 5144 7125 5153
rect 7083 5104 7084 5144
rect 7124 5104 7125 5144
rect 7083 5095 7125 5104
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 8236 4061 8276 33907
rect 8331 32528 8373 32537
rect 8331 32488 8332 32528
rect 8372 32488 8373 32528
rect 8331 32479 8373 32488
rect 8235 4052 8277 4061
rect 8235 4012 8236 4052
rect 8276 4012 8277 4052
rect 8235 4003 8277 4012
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 2379 2792 2421 2801
rect 2379 2752 2380 2792
rect 2420 2752 2421 2792
rect 2379 2743 2421 2752
rect 844 2456 884 2465
rect 844 2297 884 2416
rect 939 2456 981 2465
rect 939 2416 940 2456
rect 980 2416 981 2456
rect 939 2407 981 2416
rect 843 2288 885 2297
rect 843 2248 844 2288
rect 884 2248 885 2288
rect 843 2239 885 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 8332 1961 8372 32479
rect 11212 31529 11252 34336
rect 11788 34376 11828 34504
rect 11788 34327 11828 34336
rect 12172 34376 12212 34385
rect 12460 34376 12500 34924
rect 12212 34336 12500 34376
rect 13036 34376 13076 34385
rect 12172 34327 12212 34336
rect 11307 34292 11349 34301
rect 11307 34252 11308 34292
rect 11348 34252 11349 34292
rect 11307 34243 11349 34252
rect 11308 34158 11348 34243
rect 13036 34217 13076 34336
rect 13035 34208 13077 34217
rect 13035 34168 13036 34208
rect 13076 34168 13077 34208
rect 13035 34159 13077 34168
rect 13420 34049 13460 35176
rect 13708 34301 13748 35176
rect 13804 35216 13844 35225
rect 13804 34973 13844 35176
rect 14187 35216 14229 35225
rect 14187 35176 14188 35216
rect 14228 35176 14229 35216
rect 14187 35167 14229 35176
rect 14284 35216 14324 35225
rect 14092 35048 14132 35057
rect 14284 35048 14324 35176
rect 14132 35008 14324 35048
rect 14092 34999 14132 35008
rect 14476 34973 14516 35848
rect 15244 35839 15284 35848
rect 15531 35888 15573 35897
rect 15531 35848 15532 35888
rect 15572 35848 15573 35888
rect 15531 35839 15573 35848
rect 15628 35888 15668 35897
rect 14571 35804 14613 35813
rect 14571 35764 14572 35804
rect 14612 35764 14613 35804
rect 14571 35755 14613 35764
rect 14572 35670 14612 35755
rect 14667 35636 14709 35645
rect 14667 35596 14668 35636
rect 14708 35596 14709 35636
rect 14667 35587 14709 35596
rect 14668 35216 14708 35587
rect 14668 35141 14708 35176
rect 15532 35216 15572 35839
rect 15628 35645 15668 35848
rect 16491 35888 16533 35897
rect 16491 35848 16492 35888
rect 16532 35848 16533 35888
rect 16491 35839 16533 35848
rect 17451 35888 17493 35897
rect 17451 35848 17452 35888
rect 17492 35848 17493 35888
rect 17451 35839 17493 35848
rect 16492 35754 16532 35839
rect 17355 35804 17397 35813
rect 17355 35764 17356 35804
rect 17396 35764 17397 35804
rect 17355 35755 17397 35764
rect 15627 35636 15669 35645
rect 15627 35596 15628 35636
rect 15668 35596 15669 35636
rect 15627 35587 15669 35596
rect 16875 35636 16917 35645
rect 16875 35596 16876 35636
rect 16916 35596 16917 35636
rect 16875 35587 16917 35596
rect 14667 35132 14709 35141
rect 14667 35092 14668 35132
rect 14708 35092 14709 35132
rect 14667 35083 14709 35092
rect 13803 34964 13845 34973
rect 13803 34924 13804 34964
rect 13844 34924 13845 34964
rect 13803 34915 13845 34924
rect 14475 34964 14517 34973
rect 14475 34924 14476 34964
rect 14516 34924 14517 34964
rect 14475 34915 14517 34924
rect 15244 34376 15284 34385
rect 13707 34292 13749 34301
rect 13707 34252 13708 34292
rect 13748 34252 13749 34292
rect 13707 34243 13749 34252
rect 14187 34292 14229 34301
rect 14187 34252 14188 34292
rect 14228 34252 14229 34292
rect 14187 34243 14229 34252
rect 14188 34208 14228 34243
rect 15244 34217 15284 34336
rect 15532 34217 15572 35176
rect 15627 35216 15669 35225
rect 15627 35176 15628 35216
rect 15668 35176 15669 35216
rect 15627 35167 15669 35176
rect 15628 34376 15668 35167
rect 16683 34964 16725 34973
rect 16683 34924 16684 34964
rect 16724 34924 16725 34964
rect 16683 34915 16725 34924
rect 16684 34830 16724 34915
rect 16300 34544 16340 34553
rect 16340 34504 16532 34544
rect 16300 34495 16340 34504
rect 15628 34327 15668 34336
rect 15916 34376 15956 34385
rect 14188 34157 14228 34168
rect 15243 34208 15285 34217
rect 15243 34168 15244 34208
rect 15284 34168 15285 34208
rect 15243 34159 15285 34168
rect 15531 34208 15573 34217
rect 15531 34168 15532 34208
rect 15572 34168 15573 34208
rect 15531 34159 15573 34168
rect 13419 34040 13461 34049
rect 13419 34000 13420 34040
rect 13460 34000 13461 34040
rect 13419 33991 13461 34000
rect 15916 31529 15956 34336
rect 16011 34376 16053 34385
rect 16011 34336 16012 34376
rect 16052 34336 16053 34376
rect 16011 34327 16053 34336
rect 16492 34376 16532 34504
rect 16492 34327 16532 34336
rect 16876 34376 16916 35587
rect 17068 35216 17108 35225
rect 17068 34553 17108 35176
rect 17067 34544 17109 34553
rect 17067 34504 17068 34544
rect 17108 34504 17109 34544
rect 17067 34495 17109 34504
rect 16876 34327 16916 34336
rect 16012 34242 16052 34327
rect 17356 31697 17396 35755
rect 17452 35384 17492 35839
rect 17643 35720 17685 35729
rect 17643 35680 17644 35720
rect 17684 35680 17685 35720
rect 17643 35671 17685 35680
rect 17644 35586 17684 35671
rect 18124 35561 18164 36688
rect 18220 36679 18260 36688
rect 18891 36728 18933 36737
rect 18891 36688 18892 36728
rect 18932 36688 18933 36728
rect 18891 36679 18933 36688
rect 19083 36728 19125 36737
rect 19083 36688 19084 36728
rect 19124 36688 19125 36728
rect 19083 36679 19125 36688
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 18892 36140 18932 36679
rect 19084 36594 19124 36679
rect 19180 36653 19220 37360
rect 19276 37351 19316 37360
rect 19372 37400 19412 37411
rect 20524 37400 20564 37409
rect 19372 37325 19412 37360
rect 20332 37360 20524 37400
rect 19371 37316 19413 37325
rect 19371 37276 19372 37316
rect 19412 37276 19413 37316
rect 19371 37267 19413 37276
rect 20139 37316 20181 37325
rect 20139 37276 20140 37316
rect 20180 37276 20181 37316
rect 20139 37267 20181 37276
rect 19372 36821 19412 37267
rect 19564 37232 19604 37241
rect 19604 37192 19988 37232
rect 19564 37183 19604 37192
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 19371 36812 19413 36821
rect 19276 36772 19372 36812
rect 19412 36772 19413 36812
rect 19179 36644 19221 36653
rect 19179 36604 19180 36644
rect 19220 36604 19221 36644
rect 19179 36595 19221 36604
rect 18892 36091 18932 36100
rect 18315 35888 18357 35897
rect 18315 35848 18316 35888
rect 18356 35848 18357 35888
rect 18315 35839 18357 35848
rect 19180 35888 19220 36595
rect 19180 35839 19220 35848
rect 19276 35888 19316 36772
rect 19371 36763 19413 36772
rect 19372 36678 19412 36763
rect 19371 36476 19413 36485
rect 19371 36436 19372 36476
rect 19412 36436 19413 36476
rect 19371 36427 19413 36436
rect 19276 35839 19316 35848
rect 18123 35552 18165 35561
rect 18123 35512 18124 35552
rect 18164 35512 18165 35552
rect 18123 35503 18165 35512
rect 17452 35335 17492 35344
rect 18316 35225 18356 35839
rect 19372 35716 19412 36427
rect 19755 35888 19797 35897
rect 19755 35848 19756 35888
rect 19796 35848 19797 35888
rect 19755 35839 19797 35848
rect 19756 35754 19796 35839
rect 19948 35813 19988 37192
rect 20140 37182 20180 37267
rect 20235 36644 20277 36653
rect 20235 36604 20236 36644
rect 20276 36604 20277 36644
rect 20235 36595 20277 36604
rect 20236 36510 20276 36595
rect 20044 35888 20084 35897
rect 19947 35804 19989 35813
rect 19947 35764 19948 35804
rect 19988 35764 19989 35804
rect 19947 35755 19989 35764
rect 19372 35667 19412 35676
rect 19371 35552 19413 35561
rect 19371 35512 19372 35552
rect 19412 35512 19413 35552
rect 19371 35503 19413 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 18699 35384 18741 35393
rect 18699 35344 18700 35384
rect 18740 35344 18741 35384
rect 18699 35335 18741 35344
rect 18700 35300 18740 35335
rect 18315 35216 18357 35225
rect 18315 35176 18316 35216
rect 18356 35176 18357 35216
rect 18315 35167 18357 35176
rect 18604 35216 18644 35225
rect 18316 35082 18356 35167
rect 18604 35057 18644 35176
rect 18603 35048 18645 35057
rect 18603 35008 18604 35048
rect 18644 35008 18645 35048
rect 18603 34999 18645 35008
rect 17644 34964 17684 34973
rect 17644 34376 17684 34924
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 17740 34376 17780 34385
rect 17644 34336 17740 34376
rect 17740 34327 17780 34336
rect 18700 31697 18740 35260
rect 19180 35216 19220 35225
rect 19372 35216 19412 35503
rect 19564 35216 19604 35225
rect 19372 35176 19564 35216
rect 18988 35048 19028 35057
rect 19180 35048 19220 35176
rect 19028 35008 19220 35048
rect 18988 34999 19028 35008
rect 19564 34889 19604 35176
rect 19851 35216 19893 35225
rect 19851 35176 19852 35216
rect 19892 35176 19893 35216
rect 19851 35167 19893 35176
rect 19563 34880 19605 34889
rect 19563 34840 19564 34880
rect 19604 34840 19605 34880
rect 19563 34831 19605 34840
rect 19852 34553 19892 35167
rect 19851 34544 19893 34553
rect 19851 34504 19852 34544
rect 19892 34504 19893 34544
rect 19851 34495 19893 34504
rect 18892 34460 18932 34471
rect 18892 34385 18932 34420
rect 18891 34376 18933 34385
rect 18891 34336 18892 34376
rect 18932 34336 18933 34376
rect 18891 34327 18933 34336
rect 19371 34376 19413 34385
rect 19371 34336 19372 34376
rect 19412 34336 19413 34376
rect 19371 34327 19413 34336
rect 19852 34376 19892 34495
rect 20044 34385 20084 35848
rect 20140 35804 20180 35813
rect 20140 35057 20180 35764
rect 20332 35300 20372 37360
rect 20524 37351 20564 37360
rect 20619 37232 20661 37241
rect 20619 37192 20620 37232
rect 20660 37192 20661 37232
rect 20619 37183 20661 37192
rect 20620 36896 20660 37183
rect 20907 37148 20949 37157
rect 20907 37108 20908 37148
rect 20948 37108 20949 37148
rect 20907 37099 20949 37108
rect 20620 36847 20660 36856
rect 20427 36812 20469 36821
rect 20427 36772 20428 36812
rect 20468 36772 20469 36812
rect 20427 36763 20469 36772
rect 20428 36728 20468 36763
rect 20428 36677 20468 36688
rect 20716 36728 20756 36739
rect 20716 36653 20756 36688
rect 20908 36728 20948 37099
rect 20908 36679 20948 36688
rect 20715 36644 20757 36653
rect 20715 36604 20716 36644
rect 20756 36604 20757 36644
rect 20715 36595 20757 36604
rect 21100 36560 21140 38200
rect 21772 38156 21812 38165
rect 21292 37988 21332 37997
rect 21292 37325 21332 37948
rect 21387 37400 21429 37409
rect 21387 37360 21388 37400
rect 21428 37360 21429 37400
rect 21387 37351 21429 37360
rect 21291 37316 21333 37325
rect 21291 37276 21292 37316
rect 21332 37276 21333 37316
rect 21291 37267 21333 37276
rect 21388 36737 21428 37351
rect 21772 37325 21812 38116
rect 21964 37988 22004 37997
rect 21771 37316 21813 37325
rect 21771 37276 21772 37316
rect 21812 37276 21813 37316
rect 21771 37267 21813 37276
rect 21483 37148 21525 37157
rect 21483 37108 21484 37148
rect 21524 37108 21525 37148
rect 21483 37099 21525 37108
rect 21771 37148 21813 37157
rect 21771 37108 21772 37148
rect 21812 37108 21813 37148
rect 21771 37099 21813 37108
rect 21387 36728 21429 36737
rect 21387 36688 21388 36728
rect 21428 36688 21429 36728
rect 21387 36679 21429 36688
rect 21292 36560 21332 36569
rect 21100 36520 21292 36560
rect 21292 36511 21332 36520
rect 21003 36476 21045 36485
rect 21003 36436 21004 36476
rect 21044 36436 21045 36476
rect 21003 36427 21045 36436
rect 21004 36342 21044 36427
rect 20428 36056 20468 36065
rect 20428 35384 20468 36016
rect 20620 35972 20660 35981
rect 20620 35813 20660 35932
rect 21004 35972 21044 35981
rect 20619 35804 20661 35813
rect 20619 35764 20620 35804
rect 20660 35764 20661 35804
rect 20619 35755 20661 35764
rect 21004 35729 21044 35932
rect 21195 35888 21237 35897
rect 21195 35848 21196 35888
rect 21236 35848 21237 35888
rect 21195 35839 21237 35848
rect 20811 35720 20853 35729
rect 20811 35680 20812 35720
rect 20852 35680 20853 35720
rect 20811 35671 20853 35680
rect 21003 35720 21045 35729
rect 21003 35680 21004 35720
rect 21044 35680 21045 35720
rect 21003 35671 21045 35680
rect 21196 35720 21236 35839
rect 21291 35804 21333 35813
rect 21291 35764 21292 35804
rect 21332 35764 21333 35804
rect 21291 35755 21333 35764
rect 21196 35671 21236 35680
rect 20812 35586 20852 35671
rect 20428 35344 21044 35384
rect 20236 35260 20372 35300
rect 20139 35048 20181 35057
rect 20139 35008 20140 35048
rect 20180 35008 20181 35048
rect 20139 34999 20181 35008
rect 20140 34637 20180 34999
rect 20139 34628 20181 34637
rect 20139 34588 20140 34628
rect 20180 34588 20181 34628
rect 20139 34579 20181 34588
rect 19852 34327 19892 34336
rect 20043 34376 20085 34385
rect 20043 34336 20044 34376
rect 20084 34336 20085 34376
rect 20043 34327 20085 34336
rect 18795 34208 18837 34217
rect 18795 34168 18796 34208
rect 18836 34168 18837 34208
rect 18795 34159 18837 34168
rect 18796 31772 18836 34159
rect 19372 31772 19412 34327
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 20236 31949 20276 35260
rect 20428 35216 20468 35225
rect 20332 35176 20428 35216
rect 20332 34628 20372 35176
rect 20428 35167 20468 35176
rect 20332 34579 20372 34588
rect 20811 34544 20853 34553
rect 20811 34504 20812 34544
rect 20852 34504 20853 34544
rect 20811 34495 20853 34504
rect 20812 34376 20852 34495
rect 20812 34327 20852 34336
rect 21004 34376 21044 35344
rect 21292 35057 21332 35755
rect 21291 35048 21333 35057
rect 21291 35008 21292 35048
rect 21332 35008 21333 35048
rect 21291 34999 21333 35008
rect 21291 34880 21333 34889
rect 21291 34840 21292 34880
rect 21332 34840 21333 34880
rect 21291 34831 21333 34840
rect 21292 34376 21332 34831
rect 21388 34553 21428 36679
rect 21484 35888 21524 37099
rect 21579 37064 21621 37073
rect 21579 37024 21580 37064
rect 21620 37024 21621 37064
rect 21579 37015 21621 37024
rect 21580 36737 21620 37015
rect 21772 36954 21812 37099
rect 21772 36905 21812 36914
rect 21579 36728 21621 36737
rect 21579 36688 21580 36728
rect 21620 36688 21621 36728
rect 21579 36679 21621 36688
rect 21676 36728 21716 36737
rect 21580 36594 21620 36679
rect 21676 36317 21716 36688
rect 21771 36728 21813 36737
rect 21771 36688 21772 36728
rect 21812 36688 21813 36728
rect 21771 36679 21813 36688
rect 21675 36308 21717 36317
rect 21675 36268 21676 36308
rect 21716 36268 21717 36308
rect 21675 36259 21717 36268
rect 21580 35888 21620 35897
rect 21484 35848 21580 35888
rect 21580 35839 21620 35848
rect 21676 35888 21716 36259
rect 21772 35888 21812 36679
rect 21964 36317 22004 37948
rect 22252 36728 22292 38359
rect 23212 38156 23252 38165
rect 23596 38156 23636 38165
rect 23980 38156 24020 38165
rect 23252 38116 23540 38156
rect 23212 38107 23252 38116
rect 23404 37988 23444 37997
rect 23500 37988 23540 38116
rect 23636 38116 23924 38156
rect 23596 38107 23636 38116
rect 23788 37988 23828 37997
rect 23500 37948 23788 37988
rect 23884 37988 23924 38116
rect 24020 38116 24308 38156
rect 23980 38107 24020 38116
rect 24172 37988 24212 37997
rect 23884 37948 24172 37988
rect 23116 37400 23156 37409
rect 23404 37400 23444 37948
rect 23156 37360 23444 37400
rect 22732 37316 22772 37325
rect 22540 37232 22580 37241
rect 22540 37073 22580 37192
rect 22539 37064 22581 37073
rect 22539 37024 22540 37064
rect 22580 37024 22581 37064
rect 22539 37015 22581 37024
rect 22636 36896 22676 36905
rect 22732 36896 22772 37276
rect 22676 36856 22772 36896
rect 22923 36896 22965 36905
rect 22923 36856 22924 36896
rect 22964 36856 22965 36896
rect 22636 36847 22676 36856
rect 22923 36847 22965 36856
rect 21963 36308 22005 36317
rect 21963 36268 21964 36308
rect 22004 36268 22005 36308
rect 21963 36259 22005 36268
rect 21868 36140 21908 36149
rect 22252 36140 22292 36688
rect 22347 36728 22389 36737
rect 22347 36688 22348 36728
rect 22388 36688 22389 36728
rect 22347 36679 22389 36688
rect 22924 36728 22964 36847
rect 22924 36679 22964 36688
rect 23019 36728 23061 36737
rect 23019 36688 23020 36728
rect 23060 36688 23061 36728
rect 23019 36679 23061 36688
rect 22348 36594 22388 36679
rect 23020 36594 23060 36679
rect 22443 36476 22485 36485
rect 22443 36436 22444 36476
rect 22484 36436 22485 36476
rect 22443 36427 22485 36436
rect 21908 36100 22292 36140
rect 21868 36091 21908 36100
rect 21868 35888 21908 35897
rect 21772 35848 21868 35888
rect 21676 35839 21716 35848
rect 21868 35839 21908 35848
rect 22444 35888 22484 36427
rect 23116 35897 23156 37360
rect 23499 37064 23541 37073
rect 23499 37024 23500 37064
rect 23540 37024 23541 37064
rect 23499 37015 23541 37024
rect 23307 36980 23349 36989
rect 23307 36940 23308 36980
rect 23348 36940 23349 36980
rect 23307 36931 23349 36940
rect 23308 36821 23348 36931
rect 23307 36812 23349 36821
rect 23307 36772 23308 36812
rect 23348 36772 23349 36812
rect 23307 36763 23349 36772
rect 23212 36728 23252 36737
rect 23212 36317 23252 36688
rect 23308 36728 23348 36763
rect 23308 36677 23348 36688
rect 23500 36728 23540 37015
rect 23500 36679 23540 36688
rect 23499 36560 23541 36569
rect 23499 36520 23500 36560
rect 23540 36520 23541 36560
rect 23499 36511 23541 36520
rect 23500 36426 23540 36511
rect 23211 36308 23253 36317
rect 23211 36268 23212 36308
rect 23252 36268 23253 36308
rect 23211 36259 23253 36268
rect 22444 35839 22484 35848
rect 22827 35888 22869 35897
rect 22827 35848 22828 35888
rect 22868 35848 22869 35888
rect 22827 35839 22869 35848
rect 23115 35888 23157 35897
rect 23115 35848 23116 35888
rect 23156 35848 23157 35888
rect 23115 35839 23157 35848
rect 22828 35754 22868 35839
rect 23596 35561 23636 37948
rect 23788 37939 23828 37948
rect 23787 37400 23829 37409
rect 23787 37360 23788 37400
rect 23828 37360 23829 37400
rect 23787 37351 23829 37360
rect 23979 37400 24021 37409
rect 23979 37360 23980 37400
rect 24020 37360 24021 37400
rect 23979 37351 24021 37360
rect 23692 36728 23732 36739
rect 23692 36653 23732 36688
rect 23691 36644 23733 36653
rect 23691 36604 23692 36644
rect 23732 36604 23733 36644
rect 23691 36595 23733 36604
rect 23691 36476 23733 36485
rect 23691 36436 23692 36476
rect 23732 36436 23733 36476
rect 23691 36427 23733 36436
rect 23692 36342 23732 36427
rect 23692 35888 23732 35897
rect 23788 35888 23828 37351
rect 23980 37266 24020 37351
rect 23883 36728 23925 36737
rect 23883 36688 23884 36728
rect 23924 36688 23925 36728
rect 23883 36679 23925 36688
rect 23980 36728 24020 36737
rect 23884 36594 23924 36679
rect 23980 36569 24020 36688
rect 23979 36560 24021 36569
rect 23979 36520 23980 36560
rect 24020 36520 24021 36560
rect 23979 36511 24021 36520
rect 23883 36308 23925 36317
rect 23883 36268 23884 36308
rect 23924 36268 23925 36308
rect 23883 36259 23925 36268
rect 23732 35848 23828 35888
rect 23692 35839 23732 35848
rect 23595 35552 23637 35561
rect 23595 35512 23596 35552
rect 23636 35512 23637 35552
rect 23595 35503 23637 35512
rect 21579 35384 21621 35393
rect 21579 35344 21580 35384
rect 21620 35344 21621 35384
rect 21579 35335 21621 35344
rect 21580 35250 21620 35335
rect 23403 34628 23445 34637
rect 23403 34588 23404 34628
rect 23444 34588 23445 34628
rect 23403 34579 23445 34588
rect 21387 34544 21429 34553
rect 21387 34504 21388 34544
rect 21428 34504 21429 34544
rect 21387 34495 21429 34504
rect 22251 34544 22293 34553
rect 22251 34504 22252 34544
rect 22292 34504 22293 34544
rect 22251 34495 22293 34504
rect 23404 34544 23444 34579
rect 21388 34376 21428 34385
rect 21292 34336 21388 34376
rect 21004 34327 21044 34336
rect 21388 34327 21428 34336
rect 22252 34376 22292 34495
rect 22252 34327 22292 34336
rect 20235 31940 20277 31949
rect 20235 31900 20236 31940
rect 20276 31900 20277 31940
rect 20235 31891 20277 31900
rect 23404 31772 23444 34504
rect 23788 34376 23828 34385
rect 23884 34376 23924 36259
rect 24172 35645 24212 37948
rect 24268 35813 24308 38116
rect 26092 37568 26132 37577
rect 26132 37528 26324 37568
rect 26092 37519 26132 37528
rect 25899 37484 25941 37493
rect 25899 37444 25900 37484
rect 25940 37444 25941 37484
rect 25899 37435 25941 37444
rect 25900 37400 25940 37435
rect 25900 37349 25940 37360
rect 26092 37400 26132 37409
rect 25132 37232 25172 37241
rect 25172 37192 25268 37232
rect 25132 37183 25172 37192
rect 24363 37064 24405 37073
rect 24363 37024 24364 37064
rect 24404 37024 24405 37064
rect 24363 37015 24405 37024
rect 24364 36896 24404 37015
rect 25228 36989 25268 37192
rect 25227 36980 25269 36989
rect 25227 36940 25228 36980
rect 25268 36940 25269 36980
rect 25227 36931 25269 36940
rect 24364 36847 24404 36856
rect 24459 36896 24501 36905
rect 24459 36856 24460 36896
rect 24500 36856 24501 36896
rect 24459 36847 24501 36856
rect 24843 36896 24885 36905
rect 24843 36856 24844 36896
rect 24884 36856 24885 36896
rect 24843 36847 24885 36856
rect 25228 36896 25268 36931
rect 24460 36728 24500 36847
rect 24651 36812 24693 36821
rect 24651 36772 24652 36812
rect 24692 36772 24693 36812
rect 24651 36763 24693 36772
rect 24460 36679 24500 36688
rect 24652 36678 24692 36763
rect 24844 36140 24884 36847
rect 25228 36845 25268 36856
rect 25323 36896 25365 36905
rect 25323 36856 25324 36896
rect 25364 36856 25365 36896
rect 25323 36847 25365 36856
rect 25996 36896 26036 36905
rect 26092 36896 26132 37360
rect 26284 37400 26324 37528
rect 26284 37351 26324 37360
rect 26668 37400 26708 37411
rect 26668 37325 26708 37360
rect 26379 37316 26421 37325
rect 26379 37276 26380 37316
rect 26420 37276 26421 37316
rect 26379 37267 26421 37276
rect 26667 37316 26709 37325
rect 26667 37276 26668 37316
rect 26708 37276 26709 37316
rect 26667 37267 26709 37276
rect 26036 36856 26132 36896
rect 25996 36847 26036 36856
rect 25227 36728 25269 36737
rect 25227 36688 25228 36728
rect 25268 36688 25269 36728
rect 25227 36679 25269 36688
rect 25324 36728 25364 36847
rect 25324 36679 25364 36688
rect 25900 36728 25940 36737
rect 25228 36317 25268 36679
rect 25515 36644 25557 36653
rect 25515 36604 25516 36644
rect 25556 36604 25557 36644
rect 25515 36595 25557 36604
rect 25516 36476 25556 36595
rect 25900 36569 25940 36688
rect 26091 36728 26133 36737
rect 26091 36688 26092 36728
rect 26132 36688 26133 36728
rect 26091 36679 26133 36688
rect 26188 36728 26228 36737
rect 26092 36594 26132 36679
rect 25899 36560 25941 36569
rect 25899 36520 25900 36560
rect 25940 36520 25941 36560
rect 25899 36511 25941 36520
rect 25516 36401 25556 36436
rect 26188 36401 26228 36688
rect 25515 36392 25557 36401
rect 25515 36352 25516 36392
rect 25556 36352 25557 36392
rect 25515 36343 25557 36352
rect 26187 36392 26229 36401
rect 26187 36352 26188 36392
rect 26228 36352 26229 36392
rect 26187 36343 26229 36352
rect 26380 36317 26420 37267
rect 26764 37064 26804 38368
rect 26859 38240 26901 38249
rect 26859 38200 26860 38240
rect 26900 38200 26901 38240
rect 26859 38191 26901 38200
rect 26956 38240 26996 38368
rect 26956 38191 26996 38200
rect 27052 38324 27092 38333
rect 26860 38106 26900 38191
rect 26956 37988 26996 37997
rect 26859 37484 26901 37493
rect 26859 37444 26860 37484
rect 26900 37444 26901 37484
rect 26859 37435 26901 37444
rect 26668 37024 26804 37064
rect 26475 36980 26517 36989
rect 26475 36940 26476 36980
rect 26516 36940 26517 36980
rect 26475 36931 26517 36940
rect 26476 36728 26516 36931
rect 26668 36905 26708 37024
rect 26667 36896 26709 36905
rect 26667 36856 26668 36896
rect 26708 36856 26709 36896
rect 26860 36896 26900 37435
rect 26956 37157 26996 37948
rect 27052 37409 27092 38284
rect 27051 37400 27093 37409
rect 27051 37360 27052 37400
rect 27092 37360 27093 37400
rect 27051 37351 27093 37360
rect 27148 37232 27188 38368
rect 28875 38408 28917 38417
rect 28875 38368 28876 38408
rect 28916 38368 28917 38408
rect 28875 38359 28917 38368
rect 29259 38408 29301 38417
rect 29259 38368 29260 38408
rect 29300 38368 29301 38408
rect 29259 38359 29301 38368
rect 27339 38240 27381 38249
rect 27339 38200 27340 38240
rect 27380 38200 27381 38240
rect 27339 38191 27381 38200
rect 28491 38240 28533 38249
rect 28491 38200 28492 38240
rect 28532 38200 28533 38240
rect 28491 38191 28533 38200
rect 28876 38240 28916 38359
rect 27052 37192 27188 37232
rect 26955 37148 26997 37157
rect 26955 37108 26956 37148
rect 26996 37108 26997 37148
rect 26955 37099 26997 37108
rect 26956 36896 26996 36905
rect 26860 36856 26956 36896
rect 26667 36847 26709 36856
rect 26956 36847 26996 36856
rect 26476 36679 26516 36688
rect 26572 36728 26612 36737
rect 26572 36653 26612 36688
rect 26668 36728 26708 36847
rect 26763 36812 26805 36821
rect 26763 36772 26764 36812
rect 26804 36772 26805 36812
rect 26763 36763 26805 36772
rect 26668 36679 26708 36688
rect 26764 36728 26804 36763
rect 26764 36677 26804 36688
rect 26859 36728 26901 36737
rect 26859 36688 26860 36728
rect 26900 36688 26901 36728
rect 26859 36679 26901 36688
rect 26571 36644 26613 36653
rect 26571 36604 26572 36644
rect 26612 36604 26613 36644
rect 26571 36595 26613 36604
rect 25227 36308 25269 36317
rect 25227 36268 25228 36308
rect 25268 36268 25269 36308
rect 25227 36259 25269 36268
rect 25995 36308 26037 36317
rect 25995 36268 25996 36308
rect 26036 36268 26037 36308
rect 25995 36259 26037 36268
rect 26379 36308 26421 36317
rect 26379 36268 26380 36308
rect 26420 36268 26421 36308
rect 26379 36259 26421 36268
rect 24844 36091 24884 36100
rect 25900 35897 25940 35916
rect 25899 35888 25941 35897
rect 25996 35888 26036 36259
rect 25899 35848 25900 35888
rect 25940 35848 25996 35888
rect 25899 35839 25941 35848
rect 24267 35804 24309 35813
rect 24267 35764 24268 35804
rect 24308 35764 24309 35804
rect 24267 35755 24309 35764
rect 25612 35804 25652 35813
rect 24171 35636 24213 35645
rect 24171 35596 24172 35636
rect 24212 35596 24213 35636
rect 24171 35587 24213 35596
rect 25612 35393 25652 35764
rect 25611 35384 25653 35393
rect 25611 35344 25612 35384
rect 25652 35344 25653 35384
rect 25611 35335 25653 35344
rect 24459 35216 24501 35225
rect 24459 35176 24460 35216
rect 24500 35176 24501 35216
rect 24459 35167 24501 35176
rect 25707 35216 25749 35225
rect 25707 35176 25708 35216
rect 25748 35176 25749 35216
rect 25707 35167 25749 35176
rect 24460 35082 24500 35167
rect 25708 35082 25748 35167
rect 23979 34964 24021 34973
rect 23979 34924 23980 34964
rect 24020 34924 24021 34964
rect 23979 34915 24021 34924
rect 24844 34964 24884 34973
rect 23828 34336 23924 34376
rect 23788 34327 23828 34336
rect 23980 31772 24020 34915
rect 24460 34544 24500 34553
rect 24500 34504 24692 34544
rect 24460 34495 24500 34504
rect 24075 34376 24117 34385
rect 24075 34336 24076 34376
rect 24116 34336 24117 34376
rect 24075 34327 24117 34336
rect 24652 34376 24692 34504
rect 24652 34327 24692 34336
rect 24076 34242 24116 34327
rect 24172 34292 24212 34301
rect 24172 33797 24212 34252
rect 24844 33965 24884 34924
rect 25899 34544 25941 34553
rect 25899 34504 25900 34544
rect 25940 34504 25941 34544
rect 25899 34495 25941 34504
rect 25035 34460 25077 34469
rect 25035 34420 25036 34460
rect 25076 34420 25077 34460
rect 25035 34411 25077 34420
rect 25036 34376 25076 34411
rect 25036 34325 25076 34336
rect 25900 34376 25940 34495
rect 25996 34469 26036 35848
rect 26092 34964 26132 34973
rect 25995 34460 26037 34469
rect 25995 34420 25996 34460
rect 26036 34420 26037 34460
rect 25995 34411 26037 34420
rect 25900 34327 25940 34336
rect 24843 33956 24885 33965
rect 24843 33916 24844 33956
rect 24884 33916 24885 33956
rect 24843 33907 24885 33916
rect 24171 33788 24213 33797
rect 24171 33748 24172 33788
rect 24212 33748 24213 33788
rect 24171 33739 24213 33748
rect 26092 32537 26132 34924
rect 26572 34721 26612 36595
rect 26860 36224 26900 36679
rect 27052 36569 27092 37192
rect 27147 36980 27189 36989
rect 27147 36940 27148 36980
rect 27188 36940 27189 36980
rect 27147 36931 27189 36940
rect 27148 36728 27188 36931
rect 27244 36896 27284 36905
rect 27340 36896 27380 38191
rect 27435 38156 27477 38165
rect 27435 38116 27436 38156
rect 27476 38116 27477 38156
rect 27435 38107 27477 38116
rect 27284 36856 27380 36896
rect 27244 36847 27284 36856
rect 27148 36679 27188 36688
rect 27339 36728 27381 36737
rect 27339 36688 27340 36728
rect 27380 36688 27381 36728
rect 27339 36679 27381 36688
rect 27436 36728 27476 38107
rect 28492 38106 28532 38191
rect 28876 37493 28916 38200
rect 28972 38324 29012 38333
rect 28875 37484 28917 37493
rect 28875 37444 28876 37484
rect 28916 37444 28917 37484
rect 28875 37435 28917 37444
rect 27532 37400 27572 37409
rect 27532 36737 27572 37360
rect 28779 37316 28821 37325
rect 28779 37276 28780 37316
rect 28820 37276 28821 37316
rect 28779 37267 28821 37276
rect 28684 37232 28724 37241
rect 27628 36896 27668 36905
rect 27436 36679 27476 36688
rect 27531 36728 27573 36737
rect 27531 36688 27532 36728
rect 27572 36688 27573 36728
rect 27531 36679 27573 36688
rect 27340 36594 27380 36679
rect 27628 36653 27668 36856
rect 27915 36812 27957 36821
rect 27915 36772 27916 36812
rect 27956 36772 27957 36812
rect 27915 36763 27957 36772
rect 27724 36728 27764 36737
rect 27627 36644 27669 36653
rect 27627 36604 27628 36644
rect 27668 36604 27669 36644
rect 27627 36595 27669 36604
rect 27724 36569 27764 36688
rect 27916 36678 27956 36763
rect 28011 36644 28053 36653
rect 28011 36604 28012 36644
rect 28052 36604 28053 36644
rect 28011 36595 28053 36604
rect 27051 36560 27093 36569
rect 27051 36520 27052 36560
rect 27092 36520 27093 36560
rect 27051 36511 27093 36520
rect 27723 36560 27765 36569
rect 27723 36520 27724 36560
rect 27764 36520 27765 36560
rect 27723 36511 27765 36520
rect 27051 36392 27093 36401
rect 27051 36352 27052 36392
rect 27092 36352 27093 36392
rect 27051 36343 27093 36352
rect 26764 36184 26900 36224
rect 26764 35216 26804 36184
rect 26764 35167 26804 35176
rect 26860 35888 26900 35897
rect 26571 34712 26613 34721
rect 26571 34672 26572 34712
rect 26612 34672 26613 34712
rect 26571 34663 26613 34672
rect 26860 34553 26900 35848
rect 27052 35216 27092 36343
rect 28012 36140 28052 36595
rect 28684 36569 28724 37192
rect 28780 36905 28820 37267
rect 28779 36896 28821 36905
rect 28779 36856 28780 36896
rect 28820 36856 28821 36896
rect 28779 36847 28821 36856
rect 28972 36812 29012 38284
rect 29260 38240 29300 38359
rect 29260 38191 29300 38200
rect 29451 38240 29493 38249
rect 29451 38200 29452 38240
rect 29492 38200 29493 38240
rect 29451 38191 29493 38200
rect 31467 38240 31509 38249
rect 31467 38200 31468 38240
rect 31508 38200 31509 38240
rect 31467 38191 31509 38200
rect 38476 38240 38516 38249
rect 29452 38106 29492 38191
rect 29356 37988 29396 37997
rect 29356 37400 29396 37948
rect 29356 37351 29396 37360
rect 29451 37400 29493 37409
rect 29451 37360 29452 37400
rect 29492 37360 29493 37400
rect 29451 37351 29493 37360
rect 30316 37400 30356 37409
rect 29452 37266 29492 37351
rect 29932 37316 29972 37325
rect 29740 37232 29780 37241
rect 29932 37232 29972 37276
rect 29780 37192 29972 37232
rect 29740 37183 29780 37192
rect 30316 36905 30356 37360
rect 31180 37400 31220 37409
rect 29451 36896 29493 36905
rect 29451 36856 29452 36896
rect 29492 36856 29493 36896
rect 29451 36847 29493 36856
rect 30315 36896 30357 36905
rect 30315 36856 30316 36896
rect 30356 36856 30357 36896
rect 30315 36847 30357 36856
rect 29068 36812 29108 36821
rect 28972 36772 29068 36812
rect 29068 36763 29108 36772
rect 29452 36728 29492 36847
rect 31180 36737 31220 37360
rect 31468 36896 31508 38191
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 32331 37400 32373 37409
rect 32331 37360 32332 37400
rect 32372 37360 32373 37400
rect 32331 37351 32373 37360
rect 33675 37400 33717 37409
rect 33675 37360 33676 37400
rect 33716 37360 33717 37400
rect 33675 37351 33717 37360
rect 36651 37400 36693 37409
rect 36651 37360 36652 37400
rect 36692 37360 36693 37400
rect 36651 37351 36693 37360
rect 38188 37400 38228 37409
rect 32332 37232 32372 37351
rect 32332 37183 32372 37192
rect 31468 36847 31508 36856
rect 33676 36737 33716 37351
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 29452 36679 29492 36688
rect 30315 36728 30357 36737
rect 30315 36688 30316 36728
rect 30356 36688 30357 36728
rect 30315 36679 30357 36688
rect 31179 36728 31221 36737
rect 31179 36688 31180 36728
rect 31220 36688 31221 36728
rect 31179 36679 31221 36688
rect 32428 36728 32468 36737
rect 32812 36728 32852 36737
rect 30316 36594 30356 36679
rect 28683 36560 28725 36569
rect 28683 36520 28684 36560
rect 28724 36520 28725 36560
rect 28683 36511 28725 36520
rect 28012 36091 28052 36100
rect 32236 36140 32276 36149
rect 32428 36140 32468 36688
rect 32276 36100 32468 36140
rect 32716 36688 32812 36728
rect 32236 36091 32276 36100
rect 31084 35972 31124 35981
rect 31124 35932 31220 35972
rect 31084 35923 31124 35932
rect 27531 35720 27573 35729
rect 27531 35680 27532 35720
rect 27572 35680 27573 35720
rect 27531 35671 27573 35680
rect 30123 35720 30165 35729
rect 30123 35680 30124 35720
rect 30164 35680 30165 35720
rect 30123 35671 30165 35680
rect 27243 35384 27285 35393
rect 27243 35344 27244 35384
rect 27284 35344 27285 35384
rect 27243 35335 27285 35344
rect 27244 35250 27284 35335
rect 27052 35167 27092 35176
rect 27532 35132 27572 35671
rect 28395 35468 28437 35477
rect 28395 35428 28396 35468
rect 28436 35428 28437 35468
rect 28395 35419 28437 35428
rect 29259 35468 29301 35477
rect 29259 35428 29260 35468
rect 29300 35428 29301 35468
rect 29259 35419 29301 35428
rect 27723 35384 27765 35393
rect 27723 35344 27724 35384
rect 27764 35344 27765 35384
rect 27723 35335 27765 35344
rect 28011 35384 28053 35393
rect 28011 35344 28012 35384
rect 28052 35344 28053 35384
rect 28011 35335 28053 35344
rect 27724 35250 27764 35335
rect 28012 35216 28052 35335
rect 28396 35300 28436 35419
rect 28971 35384 29013 35393
rect 28971 35344 28972 35384
rect 29012 35344 29013 35384
rect 28971 35335 29013 35344
rect 28396 35251 28436 35260
rect 28012 35167 28052 35176
rect 28300 35216 28340 35225
rect 28300 35132 28340 35176
rect 28972 35216 29012 35335
rect 28300 35092 28820 35132
rect 27532 35083 27572 35092
rect 28684 34964 28724 34973
rect 28012 34924 28684 34964
rect 26859 34544 26901 34553
rect 26859 34504 26860 34544
rect 26900 34504 26901 34544
rect 26859 34495 26901 34504
rect 27052 34460 27092 34471
rect 27052 34385 27092 34420
rect 27051 34376 27093 34385
rect 27051 34336 27052 34376
rect 27092 34336 27093 34376
rect 27051 34327 27093 34336
rect 28012 34376 28052 34924
rect 28684 34915 28724 34924
rect 28395 34460 28437 34469
rect 28395 34420 28396 34460
rect 28436 34420 28437 34460
rect 28395 34411 28437 34420
rect 28012 34327 28052 34336
rect 28396 34376 28436 34411
rect 28780 34385 28820 35092
rect 28972 34637 29012 35176
rect 29260 35216 29300 35419
rect 29355 35384 29397 35393
rect 29355 35344 29356 35384
rect 29396 35344 29397 35384
rect 29355 35335 29397 35344
rect 29356 35300 29396 35335
rect 29356 35249 29396 35260
rect 29260 34712 29300 35176
rect 29836 35216 29876 35225
rect 29644 35048 29684 35057
rect 29836 35048 29876 35176
rect 29684 35008 29876 35048
rect 29644 34999 29684 35008
rect 29260 34672 29396 34712
rect 28971 34628 29013 34637
rect 28971 34588 28972 34628
rect 29012 34588 29013 34628
rect 28971 34579 29013 34588
rect 29259 34544 29301 34553
rect 29259 34504 29260 34544
rect 29300 34504 29301 34544
rect 29259 34495 29301 34504
rect 28396 34325 28436 34336
rect 28779 34376 28821 34385
rect 28779 34336 28780 34376
rect 28820 34336 28821 34376
rect 28779 34327 28821 34336
rect 29260 34376 29300 34495
rect 29356 34469 29396 34672
rect 29355 34460 29397 34469
rect 29355 34420 29356 34460
rect 29396 34420 29397 34460
rect 29355 34411 29397 34420
rect 29835 34460 29877 34469
rect 29835 34420 29836 34460
rect 29876 34420 29877 34460
rect 29835 34411 29877 34420
rect 29260 34327 29300 34336
rect 29547 34376 29589 34385
rect 29547 34336 29548 34376
rect 29588 34336 29589 34376
rect 29547 34327 29589 34336
rect 26091 32528 26133 32537
rect 26091 32488 26092 32528
rect 26132 32488 26133 32528
rect 26091 32479 26133 32488
rect 29548 31772 29588 34327
rect 29836 31772 29876 34411
rect 18796 31732 18849 31772
rect 19372 31732 19617 31772
rect 23404 31732 23841 31772
rect 23980 31732 24033 31772
rect 29548 31732 29601 31772
rect 17355 31688 17397 31697
rect 17355 31648 17356 31688
rect 17396 31648 17397 31688
rect 17355 31639 17397 31648
rect 18040 31688 18082 31697
rect 18040 31648 18041 31688
rect 18081 31648 18082 31688
rect 18040 31639 18082 31648
rect 18267 31688 18309 31697
rect 18267 31648 18268 31688
rect 18308 31648 18309 31688
rect 18267 31639 18309 31648
rect 18699 31688 18741 31697
rect 18699 31648 18700 31688
rect 18740 31648 18741 31688
rect 18699 31639 18741 31648
rect 11211 31520 11253 31529
rect 11211 31480 11212 31520
rect 11252 31480 11253 31520
rect 11211 31471 11253 31480
rect 15160 31520 15202 31529
rect 15160 31480 15161 31520
rect 15201 31480 15202 31520
rect 15160 31471 15202 31480
rect 15915 31520 15957 31529
rect 15915 31480 15916 31520
rect 15956 31480 15957 31520
rect 15915 31471 15957 31480
rect 15161 31374 15201 31471
rect 16312 31380 16354 31389
rect 16312 31340 16313 31380
rect 16353 31340 16354 31380
rect 18041 31374 18081 31639
rect 18268 31379 18308 31639
rect 18809 31374 18849 31732
rect 19577 31374 19617 31732
rect 23801 31374 23841 31732
rect 23993 31374 24033 31732
rect 29561 31374 29601 31732
rect 29791 31732 29876 31772
rect 30124 31772 30164 35671
rect 30219 35552 30261 35561
rect 30219 35512 30220 35552
rect 30260 35512 30261 35552
rect 30219 35503 30261 35512
rect 30220 35216 30260 35503
rect 30220 35167 30260 35176
rect 31084 35216 31124 35225
rect 31084 34553 31124 35176
rect 31180 34637 31220 35932
rect 31275 35888 31317 35897
rect 31275 35848 31276 35888
rect 31316 35848 31317 35888
rect 31275 35839 31317 35848
rect 31563 35888 31605 35897
rect 31563 35848 31564 35888
rect 31604 35848 31605 35888
rect 31563 35839 31605 35848
rect 31852 35888 31892 35897
rect 31276 35720 31316 35839
rect 31467 35804 31509 35813
rect 31467 35764 31468 35804
rect 31508 35764 31509 35804
rect 31467 35755 31509 35764
rect 31179 34628 31221 34637
rect 31179 34588 31180 34628
rect 31220 34588 31221 34628
rect 31179 34579 31221 34588
rect 31083 34544 31125 34553
rect 31083 34504 31084 34544
rect 31124 34504 31125 34544
rect 31083 34495 31125 34504
rect 30411 34460 30453 34469
rect 30411 34420 30412 34460
rect 30452 34420 30453 34460
rect 30411 34411 30453 34420
rect 30412 34326 30452 34411
rect 31276 34376 31316 35680
rect 31276 34327 31316 34336
rect 31468 31772 31508 35755
rect 31564 35754 31604 35839
rect 31852 35393 31892 35848
rect 31947 35804 31989 35813
rect 31947 35764 31948 35804
rect 31988 35764 31989 35804
rect 31947 35755 31989 35764
rect 31948 35670 31988 35755
rect 32716 35561 32756 36688
rect 32812 36679 32852 36688
rect 33675 36728 33717 36737
rect 33675 36688 33676 36728
rect 33716 36688 33717 36728
rect 33675 36679 33717 36688
rect 35116 36728 35156 36737
rect 35404 36728 35444 36737
rect 33676 36594 33716 36679
rect 34828 36476 34868 36485
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 34443 36056 34485 36065
rect 34443 36016 34444 36056
rect 34484 36016 34485 36056
rect 34443 36007 34485 36016
rect 34444 35888 34484 36007
rect 34444 35839 34484 35848
rect 34828 35813 34868 36436
rect 35116 35981 35156 36688
rect 35308 36688 35404 36728
rect 35115 35972 35157 35981
rect 35115 35932 35116 35972
rect 35156 35932 35157 35972
rect 35115 35923 35157 35932
rect 34827 35804 34869 35813
rect 34827 35764 34828 35804
rect 34868 35764 34869 35804
rect 34827 35755 34869 35764
rect 32908 35720 32948 35729
rect 32523 35552 32565 35561
rect 32523 35512 32524 35552
rect 32564 35512 32565 35552
rect 32523 35503 32565 35512
rect 32715 35552 32757 35561
rect 32715 35512 32716 35552
rect 32756 35512 32757 35552
rect 32715 35503 32757 35512
rect 31851 35384 31893 35393
rect 31851 35344 31852 35384
rect 31892 35344 31893 35384
rect 31851 35335 31893 35344
rect 32235 35384 32277 35393
rect 32235 35344 32236 35384
rect 32276 35344 32277 35384
rect 32235 35335 32277 35344
rect 32236 35250 32276 35335
rect 32236 34964 32276 34973
rect 31948 34544 31988 34553
rect 31988 34504 32180 34544
rect 31948 34495 31988 34504
rect 31564 34376 31604 34385
rect 31564 34217 31604 34336
rect 32140 34376 32180 34504
rect 32140 34327 32180 34336
rect 31660 34292 31700 34301
rect 31563 34208 31605 34217
rect 31563 34168 31564 34208
rect 31604 34168 31605 34208
rect 31563 34159 31605 34168
rect 31660 34133 31700 34252
rect 31659 34124 31701 34133
rect 31659 34084 31660 34124
rect 31700 34084 31701 34124
rect 31659 34075 31701 34084
rect 32236 31772 32276 34924
rect 32524 34376 32564 35503
rect 32908 34385 32948 35680
rect 35019 35636 35061 35645
rect 35019 35596 35020 35636
rect 35060 35596 35061 35636
rect 35019 35587 35061 35596
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 33867 35300 33909 35309
rect 33867 35260 33868 35300
rect 33908 35260 33909 35300
rect 33867 35251 33909 35260
rect 33483 35216 33525 35225
rect 33483 35176 33484 35216
rect 33524 35176 33525 35216
rect 33483 35167 33525 35176
rect 33484 35082 33524 35167
rect 33772 34964 33812 34973
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 33387 34544 33429 34553
rect 33387 34504 33388 34544
rect 33428 34504 33429 34544
rect 33387 34495 33429 34504
rect 32524 34327 32564 34336
rect 32907 34376 32949 34385
rect 32907 34336 32908 34376
rect 32948 34336 32949 34376
rect 32907 34327 32949 34336
rect 33388 34376 33428 34495
rect 33388 34327 33428 34336
rect 33003 34208 33045 34217
rect 33003 34168 33004 34208
rect 33044 34168 33045 34208
rect 33003 34159 33045 34168
rect 32907 33956 32949 33965
rect 32907 33916 32908 33956
rect 32948 33916 32949 33956
rect 32907 33907 32949 33916
rect 32908 31772 32948 33907
rect 30124 31732 30177 31772
rect 31468 31732 31521 31772
rect 29791 31374 29831 31732
rect 30137 31374 30177 31732
rect 31481 31374 31521 31732
rect 32095 31732 32276 31772
rect 32863 31732 32948 31772
rect 33004 31772 33044 34159
rect 33772 32453 33812 34924
rect 33868 34721 33908 35251
rect 34635 35216 34677 35225
rect 34635 35176 34636 35216
rect 34676 35176 34677 35216
rect 34635 35167 34677 35176
rect 35020 35216 35060 35587
rect 35020 35167 35060 35176
rect 34636 35082 34676 35167
rect 33867 34712 33909 34721
rect 35116 34712 35156 35923
rect 35308 35813 35348 36688
rect 35404 36679 35444 36688
rect 35500 36728 35540 36737
rect 35307 35804 35349 35813
rect 35307 35764 35308 35804
rect 35348 35764 35349 35804
rect 35307 35755 35349 35764
rect 35404 35804 35444 35813
rect 35404 35552 35444 35764
rect 35500 35729 35540 36688
rect 35788 36476 35828 36485
rect 35692 36436 35788 36476
rect 35499 35720 35541 35729
rect 35499 35680 35500 35720
rect 35540 35680 35541 35720
rect 35499 35671 35541 35680
rect 35692 35552 35732 36436
rect 35788 36427 35828 36436
rect 35788 35888 35828 35897
rect 35788 35813 35828 35848
rect 36652 35888 36692 37351
rect 37803 37316 37845 37325
rect 37803 37276 37804 37316
rect 37844 37276 37845 37316
rect 37803 37267 37845 37276
rect 37804 37182 37844 37267
rect 38188 36905 38228 37360
rect 38476 37241 38516 38200
rect 38763 38240 38805 38249
rect 38763 38200 38764 38240
rect 38804 38200 38805 38240
rect 38763 38191 38805 38200
rect 38860 38240 38900 38249
rect 38764 38106 38804 38191
rect 38860 37460 38900 38200
rect 39819 38240 39861 38249
rect 39819 38200 39820 38240
rect 39860 38200 39861 38240
rect 39819 38191 39861 38200
rect 41068 38240 41108 38249
rect 39148 37988 39188 37997
rect 38860 37420 38996 37460
rect 38475 37232 38517 37241
rect 38380 37192 38476 37232
rect 38516 37192 38517 37232
rect 38187 36896 38229 36905
rect 38187 36856 38188 36896
rect 38228 36856 38229 36896
rect 38187 36847 38229 36856
rect 36652 35839 36692 35848
rect 38188 35813 38228 36847
rect 38380 35981 38420 37192
rect 38475 37183 38517 37192
rect 38859 36896 38901 36905
rect 38859 36856 38860 36896
rect 38900 36856 38901 36896
rect 38859 36847 38901 36856
rect 38476 36728 38516 36737
rect 38476 36149 38516 36688
rect 38571 36728 38613 36737
rect 38571 36688 38572 36728
rect 38612 36688 38613 36728
rect 38571 36679 38613 36688
rect 38860 36728 38900 36847
rect 38860 36679 38900 36688
rect 38475 36140 38517 36149
rect 38475 36100 38476 36140
rect 38516 36100 38517 36140
rect 38475 36091 38517 36100
rect 38379 35972 38421 35981
rect 38379 35932 38380 35972
rect 38420 35932 38421 35972
rect 38379 35923 38421 35932
rect 38476 35888 38516 35897
rect 35787 35804 35829 35813
rect 35787 35764 35788 35804
rect 35828 35764 35829 35804
rect 35787 35755 35829 35764
rect 37899 35804 37941 35813
rect 37899 35764 37900 35804
rect 37940 35764 37941 35804
rect 37899 35755 37941 35764
rect 38187 35804 38229 35813
rect 38187 35764 38188 35804
rect 38228 35764 38229 35804
rect 38187 35755 38229 35764
rect 35788 35645 35828 35755
rect 37803 35720 37845 35729
rect 37803 35680 37804 35720
rect 37844 35680 37845 35720
rect 37803 35671 37845 35680
rect 35787 35636 35829 35645
rect 35787 35596 35788 35636
rect 35828 35596 35829 35636
rect 35787 35587 35829 35596
rect 37804 35586 37844 35671
rect 35404 35512 35732 35552
rect 35499 35216 35541 35225
rect 35499 35176 35500 35216
rect 35540 35176 35541 35216
rect 35499 35167 35541 35176
rect 35883 35216 35925 35225
rect 35883 35176 35884 35216
rect 35924 35176 35925 35216
rect 35883 35167 35925 35176
rect 37612 35216 37652 35225
rect 33867 34672 33868 34712
rect 33908 34672 33909 34712
rect 33867 34663 33909 34672
rect 34828 34672 35156 34712
rect 34828 34376 34868 34672
rect 35500 34628 35540 35167
rect 35500 34579 35540 34588
rect 35884 34553 35924 35167
rect 37612 35057 37652 35176
rect 37611 35048 37653 35057
rect 37611 35008 37612 35048
rect 37652 35008 37653 35048
rect 37611 34999 37653 35008
rect 37036 34964 37076 34973
rect 35883 34544 35925 34553
rect 35883 34504 35884 34544
rect 35924 34504 35925 34544
rect 35883 34495 35925 34504
rect 34828 34327 34868 34336
rect 35116 34376 35156 34385
rect 34444 34252 34580 34292
rect 34444 34133 34484 34252
rect 34540 34208 34580 34252
rect 34540 34159 34580 34168
rect 34443 34124 34485 34133
rect 34443 34084 34444 34124
rect 34484 34084 34485 34124
rect 34443 34075 34485 34084
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 35116 33965 35156 34336
rect 35212 34292 35252 34303
rect 35212 34217 35252 34252
rect 37036 34217 37076 34924
rect 37804 34964 37844 34973
rect 37323 34628 37365 34637
rect 37323 34588 37324 34628
rect 37364 34588 37365 34628
rect 37323 34579 37365 34588
rect 37324 34376 37364 34579
rect 37804 34544 37844 34924
rect 37324 34327 37364 34336
rect 37612 34504 37844 34544
rect 35211 34208 35253 34217
rect 35211 34168 35212 34208
rect 35252 34168 35253 34208
rect 35211 34159 35253 34168
rect 37035 34208 37077 34217
rect 37035 34168 37036 34208
rect 37076 34168 37077 34208
rect 37035 34159 37077 34168
rect 35115 33956 35157 33965
rect 35115 33916 35116 33956
rect 35156 33916 35157 33956
rect 35115 33907 35157 33916
rect 37612 33881 37652 34504
rect 37708 34376 37748 34385
rect 37900 34376 37940 35755
rect 38476 35645 38516 35848
rect 38475 35636 38517 35645
rect 38475 35596 38476 35636
rect 38516 35596 38517 35636
rect 38475 35587 38517 35596
rect 38476 35309 38516 35587
rect 38475 35300 38517 35309
rect 38475 35260 38476 35300
rect 38516 35260 38517 35300
rect 38475 35251 38517 35260
rect 38091 35048 38133 35057
rect 38091 35008 38092 35048
rect 38132 35008 38133 35048
rect 38091 34999 38133 35008
rect 38092 34553 38132 34999
rect 38091 34544 38133 34553
rect 38091 34504 38092 34544
rect 38132 34504 38133 34544
rect 38091 34495 38133 34504
rect 37748 34336 37940 34376
rect 38572 34376 38612 36679
rect 38667 35972 38709 35981
rect 38667 35932 38668 35972
rect 38708 35932 38709 35972
rect 38667 35923 38709 35932
rect 38668 35216 38708 35923
rect 38764 35888 38804 35899
rect 38956 35897 38996 37420
rect 39051 37400 39093 37409
rect 39051 37360 39052 37400
rect 39092 37360 39093 37400
rect 39051 37351 39093 37360
rect 39052 37266 39092 37351
rect 39148 37325 39188 37948
rect 39147 37316 39189 37325
rect 39147 37276 39148 37316
rect 39188 37276 39189 37316
rect 39147 37267 39189 37276
rect 39723 36728 39765 36737
rect 39723 36688 39724 36728
rect 39764 36688 39765 36728
rect 39723 36679 39765 36688
rect 39724 36594 39764 36679
rect 39147 36140 39189 36149
rect 39147 36100 39148 36140
rect 39188 36100 39189 36140
rect 39147 36091 39189 36100
rect 39148 36006 39188 36091
rect 38764 35813 38804 35848
rect 38860 35888 38900 35897
rect 38955 35888 38997 35897
rect 38900 35848 38956 35888
rect 38996 35848 38997 35888
rect 38860 35839 38900 35848
rect 38955 35839 38997 35848
rect 39532 35888 39572 35899
rect 38763 35804 38805 35813
rect 38763 35764 38764 35804
rect 38804 35764 38805 35804
rect 38763 35755 38805 35764
rect 38956 35754 38996 35839
rect 39532 35813 39572 35848
rect 39820 35888 39860 38191
rect 41068 37241 41108 38200
rect 41356 38240 41396 38249
rect 41260 37400 41300 37409
rect 40204 37232 40244 37241
rect 40108 37192 40204 37232
rect 40108 35897 40148 37192
rect 40204 37183 40244 37192
rect 40587 37232 40629 37241
rect 40587 37192 40588 37232
rect 40628 37192 40629 37232
rect 40587 37183 40629 37192
rect 41067 37232 41109 37241
rect 41067 37192 41068 37232
rect 41108 37192 41109 37232
rect 41067 37183 41109 37192
rect 40204 36056 40244 36065
rect 40204 35972 40244 36016
rect 40299 35972 40341 35981
rect 40204 35932 40300 35972
rect 40340 35932 40341 35972
rect 40299 35923 40341 35932
rect 39820 35839 39860 35848
rect 39915 35888 39957 35897
rect 39915 35848 39916 35888
rect 39956 35848 39957 35888
rect 39915 35839 39957 35848
rect 40107 35888 40149 35897
rect 40107 35848 40108 35888
rect 40148 35848 40149 35888
rect 40107 35839 40149 35848
rect 40395 35888 40437 35897
rect 40395 35848 40396 35888
rect 40436 35848 40437 35888
rect 40395 35839 40437 35848
rect 39531 35804 39573 35813
rect 39531 35764 39532 35804
rect 39572 35764 39573 35804
rect 39531 35755 39573 35764
rect 39916 35754 39956 35839
rect 38764 35216 38804 35225
rect 38668 35176 38764 35216
rect 38764 35167 38804 35176
rect 39052 35216 39092 35225
rect 39052 35057 39092 35176
rect 39148 35216 39188 35225
rect 39051 35048 39093 35057
rect 39051 35008 39052 35048
rect 39092 35008 39093 35048
rect 39051 34999 39093 35008
rect 37708 34327 37748 34336
rect 38572 34327 38612 34336
rect 39148 33965 39188 35176
rect 40396 35216 40436 35839
rect 40396 35167 40436 35176
rect 40588 35216 40628 37183
rect 41067 36812 41109 36821
rect 41067 36772 41068 36812
rect 41108 36772 41109 36812
rect 41067 36763 41109 36772
rect 41068 36678 41108 36763
rect 40876 36476 40916 36485
rect 40876 35897 40916 36436
rect 41260 36224 41300 37360
rect 41356 37241 41396 38200
rect 41451 38240 41493 38249
rect 41451 38200 41452 38240
rect 41492 38200 41493 38240
rect 41451 38191 41493 38200
rect 43467 38240 43509 38249
rect 43467 38200 43468 38240
rect 43508 38200 43509 38240
rect 43467 38191 43509 38200
rect 70348 38240 70388 38249
rect 41452 38106 41492 38191
rect 41740 37988 41780 37997
rect 41548 37400 41588 37409
rect 41355 37232 41397 37241
rect 41355 37192 41356 37232
rect 41396 37192 41397 37232
rect 41355 37183 41397 37192
rect 41451 36896 41493 36905
rect 41451 36856 41452 36896
rect 41492 36856 41493 36896
rect 41451 36847 41493 36856
rect 41452 36728 41492 36847
rect 41452 36679 41492 36688
rect 41548 36224 41588 37360
rect 41644 37316 41684 37327
rect 41644 37241 41684 37276
rect 41643 37232 41685 37241
rect 41643 37192 41644 37232
rect 41684 37192 41685 37232
rect 41643 37183 41685 37192
rect 41740 36821 41780 37948
rect 41932 37568 41972 37577
rect 41932 37460 41972 37528
rect 41932 37420 42164 37460
rect 42124 37400 42164 37420
rect 42124 37351 42164 37360
rect 42508 37400 42548 37409
rect 42219 37232 42261 37241
rect 42219 37192 42220 37232
rect 42260 37192 42261 37232
rect 42219 37183 42261 37192
rect 41739 36812 41781 36821
rect 41739 36772 41740 36812
rect 41780 36772 41781 36812
rect 41739 36763 41781 36772
rect 41260 36184 41492 36224
rect 41548 36184 41684 36224
rect 41356 35972 41396 35981
rect 40875 35888 40917 35897
rect 40875 35848 40876 35888
rect 40916 35848 40917 35888
rect 40875 35839 40917 35848
rect 41163 35384 41205 35393
rect 41163 35344 41164 35384
rect 41204 35344 41205 35384
rect 41163 35335 41205 35344
rect 40588 35167 40628 35176
rect 40780 35216 40820 35225
rect 40780 35048 40820 35176
rect 41164 35216 41204 35335
rect 41164 35167 41204 35176
rect 40780 35008 41204 35048
rect 39436 34964 39476 34973
rect 39436 34721 39476 34924
rect 40588 34964 40628 34973
rect 40628 34924 41108 34964
rect 40588 34915 40628 34924
rect 39435 34712 39477 34721
rect 39435 34672 39436 34712
rect 39476 34672 39477 34712
rect 39435 34663 39477 34672
rect 41068 34376 41108 34924
rect 41068 34327 41108 34336
rect 41164 34292 41204 35008
rect 41356 34973 41396 35932
rect 41452 35720 41492 36184
rect 41644 35813 41684 36184
rect 41835 35888 41877 35897
rect 41835 35848 41836 35888
rect 41876 35848 41877 35888
rect 41835 35839 41877 35848
rect 42123 35888 42165 35897
rect 42123 35848 42124 35888
rect 42164 35848 42165 35888
rect 42123 35839 42165 35848
rect 42220 35888 42260 37183
rect 42508 36905 42548 37360
rect 43372 37400 43412 37409
rect 42795 37148 42837 37157
rect 42795 37108 42796 37148
rect 42836 37108 42837 37148
rect 42795 37099 42837 37108
rect 42507 36896 42549 36905
rect 42507 36856 42508 36896
rect 42548 36856 42549 36896
rect 42507 36847 42549 36856
rect 42315 36728 42357 36737
rect 42315 36688 42316 36728
rect 42356 36688 42357 36728
rect 42315 36679 42357 36688
rect 42316 36594 42356 36679
rect 42220 35839 42260 35848
rect 41643 35804 41685 35813
rect 41643 35764 41644 35804
rect 41684 35764 41685 35804
rect 41643 35755 41685 35764
rect 41836 35754 41876 35839
rect 42124 35754 42164 35839
rect 41548 35720 41588 35729
rect 41452 35680 41548 35720
rect 41548 35477 41588 35680
rect 42508 35678 42548 35687
rect 41547 35468 41589 35477
rect 41547 35428 41548 35468
rect 41588 35428 41589 35468
rect 41547 35419 41589 35428
rect 42027 35300 42069 35309
rect 42027 35260 42028 35300
rect 42068 35260 42069 35300
rect 42027 35251 42069 35260
rect 42028 35216 42068 35251
rect 42028 35165 42068 35176
rect 41355 34964 41397 34973
rect 41355 34924 41356 34964
rect 41396 34924 41397 34964
rect 41355 34915 41397 34924
rect 41355 34796 41397 34805
rect 41355 34756 41356 34796
rect 41396 34756 41397 34796
rect 41355 34747 41397 34756
rect 41164 34243 41204 34252
rect 41260 34376 41300 34385
rect 39724 34208 39764 34217
rect 39724 33965 39764 34168
rect 41260 34133 41300 34336
rect 41356 34376 41396 34747
rect 41356 34327 41396 34336
rect 41644 34376 41684 34385
rect 41644 34133 41684 34336
rect 41836 34376 41876 34385
rect 41740 34208 41780 34217
rect 41259 34124 41301 34133
rect 41259 34084 41260 34124
rect 41300 34084 41301 34124
rect 41259 34075 41301 34084
rect 41643 34124 41685 34133
rect 41643 34084 41644 34124
rect 41684 34084 41685 34124
rect 41643 34075 41685 34084
rect 39147 33956 39189 33965
rect 39147 33916 39148 33956
rect 39188 33916 39189 33956
rect 39147 33907 39189 33916
rect 39723 33956 39765 33965
rect 39723 33916 39724 33956
rect 39764 33916 39765 33956
rect 39723 33907 39765 33916
rect 37611 33872 37653 33881
rect 37611 33832 37612 33872
rect 37652 33832 37653 33872
rect 37611 33823 37653 33832
rect 41740 32873 41780 34168
rect 41836 33461 41876 34336
rect 42220 34376 42260 34385
rect 42220 33713 42260 34336
rect 42315 34208 42357 34217
rect 42315 34168 42316 34208
rect 42356 34168 42357 34208
rect 42315 34159 42357 34168
rect 42316 34074 42356 34159
rect 42219 33704 42261 33713
rect 42219 33664 42220 33704
rect 42260 33664 42261 33704
rect 42219 33655 42261 33664
rect 42508 33461 42548 35638
rect 42796 35057 42836 37099
rect 43372 35309 43412 37360
rect 43468 36896 43508 38191
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 44523 37232 44565 37241
rect 44523 37192 44524 37232
rect 44564 37192 44565 37232
rect 44523 37183 44565 37192
rect 44524 37098 44564 37183
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 43468 36847 43508 36856
rect 44908 36772 45524 36812
rect 44908 36644 44948 36772
rect 44908 36595 44948 36604
rect 45292 36644 45332 36653
rect 45100 36476 45140 36485
rect 44236 36056 44276 36065
rect 43564 35888 43604 35897
rect 43564 35645 43604 35848
rect 43851 35888 43893 35897
rect 43851 35848 43852 35888
rect 43892 35848 43893 35888
rect 44236 35888 44276 36016
rect 44428 35888 44468 35897
rect 44236 35848 44428 35888
rect 43851 35839 43893 35848
rect 44428 35839 44468 35848
rect 44812 35888 44852 35897
rect 45100 35888 45140 36436
rect 45292 36233 45332 36604
rect 45484 36476 45524 36772
rect 45291 36224 45333 36233
rect 45291 36184 45292 36224
rect 45332 36184 45333 36224
rect 45291 36175 45333 36184
rect 44852 35848 45140 35888
rect 43563 35636 43605 35645
rect 43563 35596 43564 35636
rect 43604 35596 43605 35636
rect 43563 35587 43605 35596
rect 43852 35561 43892 35839
rect 43948 35804 43988 35813
rect 43948 35645 43988 35764
rect 43947 35636 43989 35645
rect 43947 35596 43948 35636
rect 43988 35596 43989 35636
rect 43947 35587 43989 35596
rect 43851 35552 43893 35561
rect 43851 35512 43852 35552
rect 43892 35512 43893 35552
rect 43851 35503 43893 35512
rect 43564 35384 43604 35393
rect 44427 35384 44469 35393
rect 43604 35344 43892 35384
rect 43564 35335 43604 35344
rect 43371 35300 43413 35309
rect 43371 35260 43372 35300
rect 43412 35260 43413 35300
rect 43852 35300 43892 35344
rect 44427 35344 44428 35384
rect 44468 35344 44469 35384
rect 44427 35335 44469 35344
rect 44044 35300 44084 35309
rect 43852 35260 44044 35300
rect 43371 35251 43413 35260
rect 44044 35251 44084 35260
rect 43468 35216 43508 35225
rect 42795 35048 42837 35057
rect 42795 35008 42796 35048
rect 42836 35008 42837 35048
rect 42795 34999 42837 35008
rect 42700 34376 42740 34385
rect 42796 34376 42836 34999
rect 43180 34964 43220 34973
rect 42891 34712 42933 34721
rect 42891 34672 42892 34712
rect 42932 34672 42933 34712
rect 42891 34663 42933 34672
rect 42892 34544 42932 34663
rect 42892 34495 42932 34504
rect 42892 34376 42932 34385
rect 42796 34336 42892 34376
rect 42700 34049 42740 34336
rect 42892 34327 42932 34336
rect 42699 34040 42741 34049
rect 42699 34000 42700 34040
rect 42740 34000 42741 34040
rect 42699 33991 42741 34000
rect 43180 33713 43220 34924
rect 43468 34721 43508 35176
rect 43660 35216 43700 35225
rect 43467 34712 43509 34721
rect 43467 34672 43468 34712
rect 43508 34672 43509 34712
rect 43467 34663 43509 34672
rect 43371 34544 43413 34553
rect 43660 34544 43700 35176
rect 43756 35216 43796 35225
rect 43756 35057 43796 35176
rect 44428 35216 44468 35335
rect 44428 35167 44468 35176
rect 44812 35057 44852 35848
rect 45484 35393 45524 36436
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 47979 36056 48021 36065
rect 47979 36016 47980 36056
rect 48020 36016 48021 36056
rect 47979 36007 48021 36016
rect 52972 36056 53012 36065
rect 47980 35922 48020 36007
rect 45676 35888 45716 35897
rect 45483 35384 45525 35393
rect 45483 35344 45484 35384
rect 45524 35344 45525 35384
rect 45483 35335 45525 35344
rect 45676 35309 45716 35848
rect 49516 35888 49556 35897
rect 46828 35720 46868 35729
rect 46828 35561 46868 35680
rect 47019 35720 47061 35729
rect 47019 35680 47020 35720
rect 47060 35680 47061 35720
rect 47019 35671 47061 35680
rect 46827 35552 46869 35561
rect 46827 35512 46828 35552
rect 46868 35512 46869 35552
rect 46827 35503 46869 35512
rect 45291 35300 45333 35309
rect 45291 35260 45292 35300
rect 45332 35260 45333 35300
rect 45291 35251 45333 35260
rect 45675 35300 45717 35309
rect 45675 35260 45676 35300
rect 45716 35260 45717 35300
rect 45675 35251 45717 35260
rect 45292 35216 45332 35251
rect 45292 35165 45332 35176
rect 46732 35216 46772 35225
rect 43755 35048 43797 35057
rect 43755 35008 43756 35048
rect 43796 35008 43797 35048
rect 43755 34999 43797 35008
rect 44811 35048 44853 35057
rect 44811 35008 44812 35048
rect 44852 35008 44853 35048
rect 44811 34999 44853 35008
rect 46732 34973 46772 35176
rect 47020 35216 47060 35671
rect 47595 35468 47637 35477
rect 47595 35428 47596 35468
rect 47636 35428 47637 35468
rect 47595 35419 47637 35428
rect 48267 35468 48309 35477
rect 48267 35428 48268 35468
rect 48308 35428 48309 35468
rect 48267 35419 48309 35428
rect 47020 35167 47060 35176
rect 47116 35216 47156 35225
rect 46923 35132 46965 35141
rect 46923 35092 46924 35132
rect 46964 35092 46965 35132
rect 46923 35083 46965 35092
rect 46444 34964 46484 34973
rect 46444 34553 46484 34924
rect 46539 34964 46581 34973
rect 46539 34924 46540 34964
rect 46580 34924 46581 34964
rect 46539 34915 46581 34924
rect 46731 34964 46773 34973
rect 46731 34924 46732 34964
rect 46772 34924 46773 34964
rect 46731 34915 46773 34924
rect 43371 34504 43372 34544
rect 43412 34504 43413 34544
rect 43371 34495 43413 34504
rect 43564 34504 43700 34544
rect 46443 34544 46485 34553
rect 46443 34504 46444 34544
rect 46484 34504 46485 34544
rect 43372 34410 43412 34495
rect 43564 34217 43604 34504
rect 46443 34495 46485 34504
rect 43756 34376 43796 34385
rect 43756 34217 43796 34336
rect 45196 34376 45236 34385
rect 43563 34208 43605 34217
rect 43563 34168 43564 34208
rect 43604 34168 43605 34208
rect 43563 34159 43605 34168
rect 43755 34208 43797 34217
rect 43755 34168 43756 34208
rect 43796 34168 43797 34208
rect 43755 34159 43797 34168
rect 45196 33881 45236 34336
rect 46444 34049 46484 34495
rect 46540 34376 46580 34915
rect 46924 34889 46964 35083
rect 46923 34880 46965 34889
rect 46923 34840 46924 34880
rect 46964 34840 46965 34880
rect 46923 34831 46965 34840
rect 46540 34327 46580 34336
rect 46828 34376 46868 34385
rect 46443 34040 46485 34049
rect 46443 34000 46444 34040
rect 46484 34000 46485 34040
rect 46443 33991 46485 34000
rect 45195 33872 45237 33881
rect 45195 33832 45196 33872
rect 45236 33832 45237 33872
rect 45195 33823 45237 33832
rect 43179 33704 43221 33713
rect 43179 33664 43180 33704
rect 43220 33664 43221 33704
rect 43179 33655 43221 33664
rect 46828 33629 46868 34336
rect 46924 34376 46964 34831
rect 46924 34327 46964 34336
rect 46827 33620 46869 33629
rect 46827 33580 46828 33620
rect 46868 33580 46869 33620
rect 46827 33571 46869 33580
rect 47116 33545 47156 35176
rect 47596 35132 47636 35419
rect 47980 35216 48020 35225
rect 47596 35083 47636 35092
rect 47883 35132 47925 35141
rect 47883 35092 47884 35132
rect 47924 35092 47925 35132
rect 47883 35083 47925 35092
rect 47404 34964 47444 34973
rect 47211 34628 47253 34637
rect 47211 34588 47212 34628
rect 47252 34588 47253 34628
rect 47211 34579 47253 34588
rect 47212 34494 47252 34579
rect 47404 34376 47444 34924
rect 47787 34964 47829 34973
rect 47787 34924 47788 34964
rect 47828 34924 47829 34964
rect 47787 34915 47829 34924
rect 47788 34830 47828 34915
rect 47404 34327 47444 34336
rect 47788 34376 47828 34385
rect 47884 34376 47924 35083
rect 47980 34637 48020 35176
rect 48075 34880 48117 34889
rect 48075 34840 48076 34880
rect 48116 34840 48117 34880
rect 48075 34831 48117 34840
rect 47979 34628 48021 34637
rect 47979 34588 47980 34628
rect 48020 34588 48021 34628
rect 47979 34579 48021 34588
rect 47828 34336 47924 34376
rect 47788 34327 47828 34336
rect 47499 33620 47541 33629
rect 47499 33580 47500 33620
rect 47540 33580 47541 33620
rect 47499 33571 47541 33580
rect 47115 33536 47157 33545
rect 47115 33496 47116 33536
rect 47156 33496 47157 33536
rect 47115 33487 47157 33496
rect 41835 33452 41877 33461
rect 41835 33412 41836 33452
rect 41876 33412 41877 33452
rect 41835 33403 41877 33412
rect 42507 33452 42549 33461
rect 42507 33412 42508 33452
rect 42548 33412 42549 33452
rect 42507 33403 42549 33412
rect 47500 33377 47540 33571
rect 47499 33368 47541 33377
rect 47499 33328 47500 33368
rect 47540 33328 47541 33368
rect 47499 33319 47541 33328
rect 41739 32864 41781 32873
rect 41739 32824 41740 32864
rect 41780 32824 41781 32864
rect 41739 32815 41781 32824
rect 33771 32444 33813 32453
rect 33771 32404 33772 32444
rect 33812 32404 33813 32444
rect 33771 32395 33813 32404
rect 48076 31772 48116 34831
rect 48268 32789 48308 35419
rect 49228 35309 49268 35340
rect 49227 35300 49269 35309
rect 49227 35260 49228 35300
rect 49268 35260 49269 35300
rect 49227 35251 49269 35260
rect 48364 35216 48404 35227
rect 48364 35141 48404 35176
rect 49228 35216 49268 35251
rect 48363 35132 48405 35141
rect 48363 35092 48364 35132
rect 48404 35092 48405 35132
rect 48363 35083 48405 35092
rect 49228 34805 49268 35176
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 49227 34796 49269 34805
rect 49227 34756 49228 34796
rect 49268 34756 49269 34796
rect 49227 34747 49269 34756
rect 48651 34628 48693 34637
rect 48651 34588 48652 34628
rect 48692 34588 48693 34628
rect 48651 34579 48693 34588
rect 48652 34376 48692 34579
rect 48843 34544 48885 34553
rect 48843 34504 48844 34544
rect 48884 34504 48885 34544
rect 48843 34495 48885 34504
rect 49131 34544 49173 34553
rect 49131 34504 49132 34544
rect 49172 34504 49173 34544
rect 49131 34495 49173 34504
rect 48652 34327 48692 34336
rect 48844 33629 48884 34495
rect 48843 33620 48885 33629
rect 48843 33580 48844 33620
rect 48884 33580 48885 33620
rect 48843 33571 48885 33580
rect 49132 33545 49172 34495
rect 48939 33536 48981 33545
rect 48939 33496 48940 33536
rect 48980 33496 48981 33536
rect 48939 33487 48981 33496
rect 49131 33536 49173 33545
rect 49131 33496 49132 33536
rect 49172 33496 49173 33536
rect 49131 33487 49173 33496
rect 48267 32780 48309 32789
rect 48267 32740 48268 32780
rect 48308 32740 48309 32780
rect 48267 32731 48309 32740
rect 33004 31732 33057 31772
rect 32095 31374 32135 31732
rect 32863 31374 32903 31732
rect 33017 31374 33057 31732
rect 47993 31732 48116 31772
rect 48940 31772 48980 33487
rect 49131 33368 49173 33377
rect 49131 33328 49132 33368
rect 49172 33328 49173 33368
rect 49131 33319 49173 33328
rect 49132 31772 49172 33319
rect 49516 33125 49556 35848
rect 52300 35888 52340 35897
rect 52300 35729 52340 35848
rect 52588 35888 52628 35897
rect 50187 35720 50229 35729
rect 50187 35680 50188 35720
rect 50228 35680 50229 35720
rect 50187 35671 50229 35680
rect 52299 35720 52341 35729
rect 52299 35680 52300 35720
rect 52340 35680 52341 35720
rect 52299 35671 52341 35680
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 50188 34973 50228 35671
rect 50572 35216 50612 35225
rect 50187 34964 50229 34973
rect 50187 34924 50188 34964
rect 50228 34924 50229 34964
rect 50187 34915 50229 34924
rect 50379 34964 50421 34973
rect 50379 34924 50380 34964
rect 50420 34924 50421 34964
rect 50379 34915 50421 34924
rect 49803 34544 49845 34553
rect 49803 34504 49804 34544
rect 49844 34504 49845 34544
rect 49803 34495 49845 34504
rect 49804 34410 49844 34495
rect 50092 34376 50132 34385
rect 50188 34376 50228 34915
rect 50380 34830 50420 34915
rect 50572 34628 50612 35176
rect 50956 35216 50996 35227
rect 50956 35141 50996 35176
rect 51820 35216 51860 35225
rect 50955 35132 50997 35141
rect 50955 35092 50956 35132
rect 50996 35092 50997 35132
rect 50955 35083 50997 35092
rect 51820 34721 51860 35176
rect 52588 34964 52628 35848
rect 52683 35804 52725 35813
rect 52683 35764 52684 35804
rect 52724 35764 52725 35804
rect 52683 35755 52725 35764
rect 52684 35670 52724 35755
rect 52972 35468 53012 36016
rect 53932 36056 53972 36065
rect 53260 35888 53300 35897
rect 53260 35729 53300 35848
rect 53548 35888 53588 35897
rect 53548 35813 53588 35848
rect 53547 35804 53589 35813
rect 53547 35764 53548 35804
rect 53588 35764 53589 35804
rect 53547 35755 53589 35764
rect 53644 35804 53684 35813
rect 53259 35720 53301 35729
rect 53259 35680 53260 35720
rect 53300 35680 53301 35720
rect 53259 35671 53301 35680
rect 52972 35428 53204 35468
rect 53164 35300 53204 35428
rect 53548 35384 53588 35755
rect 53644 35468 53684 35764
rect 53644 35428 53876 35468
rect 53548 35344 53780 35384
rect 53164 35251 53204 35260
rect 53548 35216 53588 35225
rect 53548 35141 53588 35176
rect 53547 35132 53589 35141
rect 53547 35092 53548 35132
rect 53588 35092 53589 35132
rect 53547 35083 53589 35092
rect 52972 34964 53012 34973
rect 52588 34924 52972 34964
rect 51915 34796 51957 34805
rect 51915 34756 51916 34796
rect 51956 34756 51957 34796
rect 51915 34747 51957 34756
rect 51819 34712 51861 34721
rect 51819 34672 51820 34712
rect 51860 34672 51861 34712
rect 51819 34663 51861 34672
rect 50764 34628 50804 34637
rect 50572 34588 50764 34628
rect 50764 34579 50804 34588
rect 51916 34628 51956 34747
rect 51916 34579 51956 34588
rect 50379 34544 50421 34553
rect 50379 34504 50380 34544
rect 50420 34504 50421 34544
rect 50379 34495 50421 34504
rect 51531 34544 51573 34553
rect 51531 34504 51532 34544
rect 51572 34504 51573 34544
rect 51531 34495 51573 34504
rect 52779 34544 52821 34553
rect 52779 34504 52780 34544
rect 52820 34504 52821 34544
rect 52779 34495 52821 34504
rect 50132 34336 50228 34376
rect 50380 34376 50420 34495
rect 50092 34327 50132 34336
rect 50380 34327 50420 34336
rect 51532 34376 51572 34495
rect 50476 34292 50516 34301
rect 50476 34208 50516 34252
rect 51532 34217 51572 34336
rect 52780 34376 52820 34495
rect 52780 34327 52820 34336
rect 50380 34168 50516 34208
rect 51531 34208 51573 34217
rect 51531 34168 51532 34208
rect 51572 34168 51573 34208
rect 50380 34049 50420 34168
rect 51531 34159 51573 34168
rect 52491 34208 52533 34217
rect 52491 34168 52492 34208
rect 52532 34168 52533 34208
rect 52491 34159 52533 34168
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 50379 34040 50421 34049
rect 50379 34000 50380 34040
rect 50420 34000 50421 34040
rect 50379 33991 50421 34000
rect 52492 33629 52532 34159
rect 52972 34049 53012 34924
rect 53548 34133 53588 35083
rect 53740 34973 53780 35344
rect 53739 34964 53781 34973
rect 53739 34924 53740 34964
rect 53780 34924 53781 34964
rect 53739 34915 53781 34924
rect 53643 34712 53685 34721
rect 53643 34672 53644 34712
rect 53684 34672 53685 34712
rect 53643 34663 53685 34672
rect 53644 34376 53684 34663
rect 53644 34327 53684 34336
rect 53547 34124 53589 34133
rect 53547 34084 53548 34124
rect 53588 34084 53589 34124
rect 53547 34075 53589 34084
rect 52971 34040 53013 34049
rect 52971 34000 52972 34040
rect 53012 34000 53013 34040
rect 52971 33991 53013 34000
rect 52491 33620 52533 33629
rect 52491 33580 52492 33620
rect 52532 33580 52533 33620
rect 52491 33571 52533 33580
rect 49515 33116 49557 33125
rect 49515 33076 49516 33116
rect 49556 33076 49557 33116
rect 49515 33067 49557 33076
rect 52972 31772 53012 33991
rect 53740 31772 53780 34915
rect 53836 34049 53876 35428
rect 53932 34376 53972 36016
rect 65259 35972 65301 35981
rect 65259 35932 65260 35972
rect 65300 35932 65301 35972
rect 65259 35923 65301 35932
rect 65260 35561 65300 35923
rect 70348 35897 70388 38200
rect 70540 37988 70580 37997
rect 70580 37948 70676 37988
rect 70540 37939 70580 37948
rect 70636 37409 70676 37948
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 70635 37400 70677 37409
rect 70635 37360 70636 37400
rect 70676 37360 70677 37400
rect 70635 37351 70677 37360
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 93328 36896 93370 36905
rect 93328 36856 93329 36896
rect 93369 36856 93370 36896
rect 93328 36847 93370 36856
rect 91216 36812 91258 36821
rect 91216 36772 91217 36812
rect 91257 36772 91258 36812
rect 91216 36763 91258 36772
rect 74091 36728 74133 36737
rect 74091 36688 74092 36728
rect 74132 36688 74133 36728
rect 74091 36679 74133 36688
rect 83499 36728 83541 36737
rect 83499 36688 83500 36728
rect 83540 36688 83541 36728
rect 83499 36679 83541 36688
rect 65931 35888 65973 35897
rect 65931 35848 65932 35888
rect 65972 35848 65973 35888
rect 65931 35839 65973 35848
rect 70347 35888 70389 35897
rect 70347 35848 70348 35888
rect 70388 35848 70389 35888
rect 70347 35839 70389 35848
rect 72267 35888 72309 35897
rect 72267 35848 72268 35888
rect 72308 35848 72309 35888
rect 72267 35839 72309 35848
rect 73899 35888 73941 35897
rect 73899 35848 73900 35888
rect 73940 35848 73941 35888
rect 73899 35839 73941 35848
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 65259 35552 65301 35561
rect 65259 35512 65260 35552
rect 65300 35512 65301 35552
rect 65259 35503 65301 35512
rect 54412 35216 54452 35225
rect 54412 34721 54452 35176
rect 55563 34964 55605 34973
rect 55563 34924 55564 34964
rect 55604 34924 55605 34964
rect 55563 34915 55605 34924
rect 55564 34830 55604 34915
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 54411 34712 54453 34721
rect 54411 34672 54412 34712
rect 54452 34672 54453 34712
rect 54411 34663 54453 34672
rect 55371 34712 55413 34721
rect 55371 34672 55372 34712
rect 55412 34672 55413 34712
rect 55371 34663 55413 34672
rect 54124 34376 54164 34385
rect 53932 34336 54124 34376
rect 54124 34327 54164 34336
rect 54508 34376 54548 34385
rect 54508 34133 54548 34336
rect 55372 34376 55412 34663
rect 65932 34553 65972 35839
rect 72268 35754 72308 35839
rect 72652 35720 72692 35729
rect 72652 35225 72692 35680
rect 72651 35216 72693 35225
rect 72651 35176 72652 35216
rect 72692 35176 72693 35216
rect 72651 35167 72693 35176
rect 61515 34544 61557 34553
rect 61515 34504 61516 34544
rect 61556 34504 61557 34544
rect 61515 34495 61557 34504
rect 65931 34544 65973 34553
rect 65931 34504 65932 34544
rect 65972 34504 65973 34544
rect 65931 34495 65973 34504
rect 54507 34124 54549 34133
rect 54507 34084 54508 34124
rect 54548 34084 54549 34124
rect 54507 34075 54549 34084
rect 53835 34040 53877 34049
rect 53835 34000 53836 34040
rect 53876 34000 53877 34040
rect 53835 33991 53877 34000
rect 53836 33377 53876 33991
rect 53835 33368 53877 33377
rect 53835 33328 53836 33368
rect 53876 33328 53877 33368
rect 53835 33319 53877 33328
rect 55372 32453 55412 34336
rect 61516 34376 61556 34495
rect 61516 34327 61556 34336
rect 62476 34376 62516 34385
rect 56524 34208 56564 34217
rect 56524 34049 56564 34168
rect 56523 34040 56565 34049
rect 56523 34000 56524 34040
rect 56564 34000 56565 34040
rect 56523 33991 56565 34000
rect 62476 32453 62516 34336
rect 63340 34376 63380 34385
rect 63340 33125 63380 34336
rect 64683 34376 64725 34385
rect 64683 34336 64684 34376
rect 64724 34336 64725 34376
rect 64683 34327 64725 34336
rect 65932 34376 65972 34495
rect 65932 34327 65972 34336
rect 66892 34376 66932 34385
rect 64684 34242 64724 34327
rect 66892 34217 66932 34336
rect 66891 34208 66933 34217
rect 66891 34168 66892 34208
rect 66932 34168 66933 34208
rect 66891 34159 66933 34168
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 63339 33116 63381 33125
rect 63339 33076 63340 33116
rect 63380 33076 63381 33116
rect 63339 33067 63381 33076
rect 63340 32621 63380 33067
rect 63339 32612 63381 32621
rect 63339 32572 63340 32612
rect 63380 32572 63381 32612
rect 63339 32563 63381 32572
rect 55371 32444 55413 32453
rect 55371 32404 55372 32444
rect 55412 32404 55413 32444
rect 55371 32395 55413 32404
rect 62475 32444 62517 32453
rect 62475 32404 62476 32444
rect 62516 32404 62517 32444
rect 62475 32395 62517 32404
rect 48940 31732 48993 31772
rect 49132 31732 49185 31772
rect 52972 31732 53025 31772
rect 53740 31732 53793 31772
rect 47993 31374 48033 31732
rect 48953 31374 48993 31732
rect 49145 31374 49185 31732
rect 52985 31374 53025 31732
rect 53753 31374 53793 31732
rect 16312 31331 16354 31340
rect 73900 24464 73940 35839
rect 74092 24632 74132 36679
rect 83307 36644 83349 36653
rect 83307 36604 83308 36644
rect 83348 36604 83349 36644
rect 83307 36595 83349 36604
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 79563 35636 79605 35645
rect 79563 35596 79564 35636
rect 79604 35596 79605 35636
rect 79563 35587 79605 35596
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 79564 33797 79604 35587
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 81771 35384 81813 35393
rect 81771 35344 81772 35384
rect 81812 35344 81813 35384
rect 81771 35335 81813 35344
rect 81196 34376 81236 34385
rect 80812 34292 80852 34301
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 79563 33788 79605 33797
rect 79563 33748 79564 33788
rect 79604 33748 79605 33788
rect 79563 33739 79605 33748
rect 80139 33788 80181 33797
rect 80139 33748 80140 33788
rect 80180 33748 80181 33788
rect 80139 33739 80181 33748
rect 79755 33704 79797 33713
rect 79755 33664 79756 33704
rect 79796 33664 79797 33704
rect 79755 33655 79797 33664
rect 80044 33704 80084 33715
rect 79756 33570 79796 33655
rect 80044 33629 80084 33664
rect 80140 33654 80180 33739
rect 80715 33704 80757 33713
rect 80715 33664 80716 33704
rect 80756 33664 80757 33704
rect 80715 33655 80757 33664
rect 80043 33620 80085 33629
rect 80043 33580 80044 33620
rect 80084 33580 80085 33620
rect 80043 33571 80085 33580
rect 80427 33536 80469 33545
rect 80427 33496 80428 33536
rect 80468 33496 80469 33536
rect 80427 33487 80469 33496
rect 80428 33402 80468 33487
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 80428 32948 80468 32957
rect 80428 32789 80468 32908
rect 77355 32780 77397 32789
rect 77355 32740 77356 32780
rect 77396 32740 77397 32780
rect 77355 32731 77397 32740
rect 80427 32780 80469 32789
rect 80427 32740 80428 32780
rect 80468 32740 80469 32780
rect 80427 32731 80469 32740
rect 76107 32612 76149 32621
rect 76107 32572 76108 32612
rect 76148 32572 76149 32612
rect 76107 32563 76149 32572
rect 74764 28328 74804 28337
rect 76108 28328 76148 32563
rect 74804 28288 75572 28328
rect 74764 28279 74804 28288
rect 74132 24592 74420 24632
rect 74092 24583 74132 24592
rect 73900 24424 74228 24464
rect 74188 23792 74228 24424
rect 74188 23120 74228 23752
rect 74188 23071 74228 23080
rect 74380 22868 74420 24592
rect 74668 23624 74708 23633
rect 74476 22868 74516 22877
rect 74380 22828 74476 22868
rect 18617 7220 18657 7434
rect 20537 7220 20577 7434
rect 22841 7220 22881 7434
rect 23225 7220 23265 7434
rect 18412 7180 18657 7220
rect 20524 7180 20577 7220
rect 22444 7180 22881 7220
rect 23212 7180 23265 7220
rect 23452 7220 23492 7421
rect 23609 7220 23649 7434
rect 23801 7220 23841 7434
rect 23993 7220 24033 7434
rect 25721 7220 25761 7434
rect 25913 7220 25953 7434
rect 23452 7180 23540 7220
rect 16587 7160 16629 7169
rect 16587 7120 16588 7160
rect 16628 7120 16629 7160
rect 16587 7111 16629 7120
rect 15819 7076 15861 7085
rect 15819 7036 15820 7076
rect 15860 7036 15861 7076
rect 15819 7027 15861 7036
rect 12363 5396 12405 5405
rect 12363 5356 12364 5396
rect 12404 5356 12405 5396
rect 12363 5347 12405 5356
rect 12364 5153 12404 5347
rect 12363 5144 12405 5153
rect 12363 5104 12364 5144
rect 12404 5104 12405 5144
rect 12363 5095 12405 5104
rect 15820 4649 15860 7027
rect 16588 6665 16628 7111
rect 16395 6656 16437 6665
rect 16395 6616 16396 6656
rect 16436 6616 16437 6656
rect 16395 6607 16437 6616
rect 16587 6656 16629 6665
rect 16587 6616 16588 6656
rect 16628 6616 16629 6656
rect 16587 6607 16629 6616
rect 17163 6656 17205 6665
rect 17163 6616 17164 6656
rect 17204 6616 17205 6656
rect 17163 6607 17205 6616
rect 16012 4976 16052 4985
rect 15819 4640 15861 4649
rect 15819 4600 15820 4640
rect 15860 4600 15861 4640
rect 15819 4591 15861 4600
rect 16012 4397 16052 4936
rect 16396 4976 16436 6607
rect 16875 5816 16917 5825
rect 16875 5776 16876 5816
rect 16916 5776 16917 5816
rect 16875 5767 16917 5776
rect 16011 4388 16053 4397
rect 16011 4348 16012 4388
rect 16052 4348 16053 4388
rect 16011 4339 16053 4348
rect 16396 4229 16436 4936
rect 16587 4640 16629 4649
rect 16587 4600 16588 4640
rect 16628 4600 16629 4640
rect 16587 4591 16629 4600
rect 16395 4220 16437 4229
rect 16395 4180 16396 4220
rect 16436 4180 16437 4220
rect 16395 4171 16437 4180
rect 16588 4136 16628 4591
rect 16876 4136 16916 5767
rect 16971 5312 17013 5321
rect 16971 5272 16972 5312
rect 17012 5272 17013 5312
rect 16971 5263 17013 5272
rect 16628 4096 16820 4136
rect 16588 4087 16628 4096
rect 16780 3464 16820 4096
rect 16876 4087 16916 4096
rect 16972 4136 17012 5263
rect 17164 4556 17204 6607
rect 18412 5321 18452 7180
rect 19947 6656 19989 6665
rect 19947 6616 19948 6656
rect 19988 6616 19989 6656
rect 19947 6607 19989 6616
rect 19948 5993 19988 6607
rect 19947 5984 19989 5993
rect 19947 5944 19948 5984
rect 19988 5944 19989 5984
rect 19947 5935 19989 5944
rect 18411 5312 18453 5321
rect 18411 5272 18412 5312
rect 18452 5272 18453 5312
rect 18411 5263 18453 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 18412 5144 18452 5263
rect 18412 5095 18452 5104
rect 17260 4965 17300 4974
rect 17260 4817 17300 4925
rect 17259 4808 17301 4817
rect 17259 4768 17260 4808
rect 17300 4768 17301 4808
rect 17259 4759 17301 4768
rect 18699 4808 18741 4817
rect 18699 4768 18700 4808
rect 18740 4768 18741 4808
rect 18699 4759 18741 4768
rect 18232 4556 18600 4565
rect 17164 4516 17396 4556
rect 17259 4388 17301 4397
rect 17259 4348 17260 4388
rect 17300 4348 17301 4388
rect 17259 4339 17301 4348
rect 17260 4254 17300 4339
rect 17012 4096 17204 4136
rect 16972 4087 17012 4096
rect 17164 3884 17204 4096
rect 17164 3844 17300 3884
rect 17260 3491 17300 3844
rect 17356 3548 17396 4516
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 17835 4220 17877 4229
rect 17835 4180 17836 4220
rect 17876 4180 17877 4220
rect 17835 4171 17877 4180
rect 17836 4136 17876 4171
rect 18700 4145 18740 4759
rect 19852 4304 19892 4313
rect 19948 4304 19988 5935
rect 20235 4640 20277 4649
rect 20235 4600 20236 4640
rect 20276 4600 20277 4640
rect 20235 4591 20277 4600
rect 19892 4264 19988 4304
rect 19852 4255 19892 4264
rect 17836 4085 17876 4096
rect 18699 4136 18741 4145
rect 18699 4096 18700 4136
rect 18740 4096 18741 4136
rect 18699 4087 18741 4096
rect 17452 4052 17492 4061
rect 17492 4012 17684 4052
rect 17452 4003 17492 4012
rect 17356 3499 17396 3508
rect 16972 3464 17012 3473
rect 16780 3424 16972 3464
rect 17260 3442 17300 3451
rect 16972 3415 17012 3424
rect 17644 3296 17684 4012
rect 18700 4002 18740 4087
rect 20044 4052 20084 4061
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 20044 3305 20084 4012
rect 20236 3464 20276 4591
rect 20427 4220 20469 4229
rect 20427 4180 20428 4220
rect 20468 4180 20469 4220
rect 20427 4171 20469 4180
rect 20428 4136 20468 4171
rect 20428 3473 20468 4096
rect 20524 3977 20564 7180
rect 21195 6572 21237 6581
rect 21195 6532 21196 6572
rect 21236 6532 21237 6572
rect 21195 6523 21237 6532
rect 20619 4220 20661 4229
rect 20619 4180 20620 4220
rect 20660 4180 20661 4220
rect 20619 4171 20661 4180
rect 20523 3968 20565 3977
rect 20523 3928 20524 3968
rect 20564 3928 20565 3968
rect 20523 3919 20565 3928
rect 20236 3415 20276 3424
rect 20427 3464 20469 3473
rect 20427 3424 20428 3464
rect 20468 3424 20469 3464
rect 20427 3415 20469 3424
rect 20524 3464 20564 3919
rect 20620 3548 20660 4171
rect 20620 3499 20660 3508
rect 20524 3415 20564 3424
rect 21196 3380 21236 6523
rect 21771 5312 21813 5321
rect 21771 5272 21772 5312
rect 21812 5272 21813 5312
rect 21771 5263 21813 5272
rect 21772 5060 21812 5263
rect 21388 4976 21428 4985
rect 21388 4649 21428 4936
rect 21676 4976 21716 4985
rect 21579 4724 21621 4733
rect 21579 4684 21580 4724
rect 21620 4684 21621 4724
rect 21579 4675 21621 4684
rect 21387 4640 21429 4649
rect 21387 4600 21388 4640
rect 21428 4600 21429 4640
rect 21387 4591 21429 4600
rect 21291 4136 21333 4145
rect 21291 4096 21292 4136
rect 21332 4096 21333 4136
rect 21291 4087 21333 4096
rect 21292 4002 21332 4087
rect 21580 3548 21620 4675
rect 21676 4229 21716 4936
rect 21675 4220 21717 4229
rect 21675 4180 21676 4220
rect 21716 4180 21717 4220
rect 21675 4171 21717 4180
rect 21580 3499 21620 3508
rect 21196 3331 21236 3340
rect 17644 3247 17684 3256
rect 20043 3296 20085 3305
rect 20043 3256 20044 3296
rect 20084 3256 20085 3296
rect 20043 3247 20085 3256
rect 20907 3296 20949 3305
rect 20907 3256 20908 3296
rect 20948 3256 20949 3296
rect 20907 3247 20949 3256
rect 20908 3162 20948 3247
rect 21388 3212 21428 3221
rect 21428 3172 21524 3212
rect 21388 3163 21428 3172
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 21484 2708 21524 3172
rect 21484 2549 21524 2668
rect 21483 2540 21525 2549
rect 21483 2500 21484 2540
rect 21524 2500 21525 2540
rect 21483 2491 21525 2500
rect 21676 2456 21716 2465
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 21676 2120 21716 2416
rect 21772 2372 21812 5020
rect 22059 4724 22101 4733
rect 22059 4684 22060 4724
rect 22100 4684 22101 4724
rect 22059 4675 22101 4684
rect 22060 4590 22100 4675
rect 22444 4388 22484 7180
rect 23212 5321 23252 7180
rect 23211 5312 23253 5321
rect 23211 5272 23212 5312
rect 23252 5272 23253 5312
rect 23211 5263 23253 5272
rect 23403 4724 23445 4733
rect 23403 4684 23404 4724
rect 23444 4684 23445 4724
rect 23403 4675 23445 4684
rect 22731 4640 22773 4649
rect 22731 4600 22732 4640
rect 22772 4600 22773 4640
rect 22731 4591 22773 4600
rect 22444 4229 22484 4348
rect 22443 4220 22485 4229
rect 22443 4180 22444 4220
rect 22484 4180 22485 4220
rect 22443 4171 22485 4180
rect 21963 3464 22005 3473
rect 21963 3424 21964 3464
rect 22004 3424 22005 3464
rect 21963 3415 22005 3424
rect 22251 3464 22293 3473
rect 22251 3424 22252 3464
rect 22292 3424 22293 3464
rect 22251 3415 22293 3424
rect 21964 3330 22004 3415
rect 22252 2624 22292 3415
rect 22252 2575 22292 2584
rect 21868 2540 21908 2549
rect 21908 2500 22196 2540
rect 21868 2491 21908 2500
rect 21772 2332 22100 2372
rect 21771 2120 21813 2129
rect 21676 2080 21772 2120
rect 21812 2080 21813 2120
rect 21771 2071 21813 2080
rect 8331 1952 8373 1961
rect 8331 1912 8332 1952
rect 8372 1912 8373 1952
rect 8331 1903 8373 1912
rect 21772 1952 21812 2071
rect 21772 1903 21812 1912
rect 22060 1952 22100 2332
rect 22156 2204 22196 2500
rect 22156 2164 22484 2204
rect 22155 2036 22197 2045
rect 22155 1996 22156 2036
rect 22196 1996 22197 2036
rect 22155 1987 22197 1996
rect 22060 1903 22100 1912
rect 22156 1902 22196 1987
rect 22444 1784 22484 2164
rect 22732 2129 22772 4591
rect 22827 4136 22869 4145
rect 22827 4096 22828 4136
rect 22868 4096 22869 4136
rect 22827 4087 22869 4096
rect 23404 4136 23444 4675
rect 23404 4087 23444 4096
rect 22828 3464 22868 4087
rect 22868 3424 23156 3464
rect 22828 3415 22868 3424
rect 23019 2708 23061 2717
rect 23019 2668 23020 2708
rect 23060 2668 23061 2708
rect 23019 2659 23061 2668
rect 22731 2120 22773 2129
rect 22731 2080 22732 2120
rect 22772 2080 22773 2120
rect 22731 2071 22773 2080
rect 22732 1952 22772 2071
rect 23020 2045 23060 2659
rect 23116 2624 23156 3424
rect 23500 2717 23540 7180
rect 23596 7180 23649 7220
rect 23788 7180 23841 7220
rect 23980 7180 24033 7220
rect 25708 7180 25761 7220
rect 25900 7180 25953 7220
rect 26332 7220 26372 7421
rect 31708 7220 31748 7421
rect 26332 7180 26384 7220
rect 31708 7180 31796 7220
rect 23499 2708 23541 2717
rect 23499 2668 23500 2708
rect 23540 2668 23541 2708
rect 23499 2659 23541 2668
rect 23116 2575 23156 2584
rect 23596 2129 23636 7180
rect 23788 6833 23828 7180
rect 23787 6824 23829 6833
rect 23787 6784 23788 6824
rect 23828 6784 23829 6824
rect 23787 6775 23829 6784
rect 23980 5993 24020 7180
rect 25708 6917 25748 7180
rect 25707 6908 25749 6917
rect 25707 6868 25708 6908
rect 25748 6868 25749 6908
rect 25707 6859 25749 6868
rect 23979 5984 24021 5993
rect 23979 5944 23980 5984
rect 24020 5944 24021 5984
rect 23979 5935 24021 5944
rect 23979 5312 24021 5321
rect 23979 5272 23980 5312
rect 24020 5272 24021 5312
rect 23979 5263 24021 5272
rect 24363 5312 24405 5321
rect 24363 5272 24364 5312
rect 24404 5272 24405 5312
rect 24363 5263 24405 5272
rect 23788 4136 23828 4145
rect 23788 3473 23828 4096
rect 23980 3632 24020 5263
rect 24076 4976 24116 4985
rect 24076 4649 24116 4936
rect 24364 4976 24404 5263
rect 24364 4927 24404 4936
rect 24460 4976 24500 4985
rect 24075 4640 24117 4649
rect 24075 4600 24076 4640
rect 24116 4600 24117 4640
rect 24075 4591 24117 4600
rect 24460 3977 24500 4936
rect 25708 4976 25748 4985
rect 25228 4892 25268 4901
rect 25228 4733 25268 4852
rect 25419 4808 25461 4817
rect 25419 4768 25420 4808
rect 25460 4768 25461 4808
rect 25419 4759 25461 4768
rect 24747 4724 24789 4733
rect 24747 4684 24748 4724
rect 24788 4684 24789 4724
rect 24747 4675 24789 4684
rect 25227 4724 25269 4733
rect 25227 4684 25228 4724
rect 25268 4684 25269 4724
rect 25227 4675 25269 4684
rect 24748 4590 24788 4675
rect 25420 4674 25460 4759
rect 25708 4649 25748 4936
rect 25707 4640 25749 4649
rect 25707 4600 25708 4640
rect 25748 4600 25749 4640
rect 25707 4591 25749 4600
rect 24651 4136 24693 4145
rect 24651 4096 24652 4136
rect 24692 4096 24693 4136
rect 24651 4087 24693 4096
rect 24652 4002 24692 4087
rect 24459 3968 24501 3977
rect 24459 3928 24460 3968
rect 24500 3928 24501 3968
rect 24459 3919 24501 3928
rect 25708 3893 25748 4591
rect 25803 3968 25845 3977
rect 25803 3928 25804 3968
rect 25844 3928 25845 3968
rect 25803 3919 25845 3928
rect 25707 3884 25749 3893
rect 25707 3844 25708 3884
rect 25748 3844 25749 3884
rect 25707 3835 25749 3844
rect 23980 3583 24020 3592
rect 23787 3464 23829 3473
rect 23787 3424 23788 3464
rect 23828 3424 23829 3464
rect 23787 3415 23829 3424
rect 23979 3464 24021 3473
rect 23979 3424 23980 3464
rect 24020 3424 24021 3464
rect 23979 3415 24021 3424
rect 23115 2120 23157 2129
rect 23115 2080 23116 2120
rect 23156 2080 23157 2120
rect 23115 2071 23157 2080
rect 23595 2120 23637 2129
rect 23595 2080 23596 2120
rect 23636 2080 23637 2120
rect 23595 2071 23637 2080
rect 23019 2036 23061 2045
rect 23019 1996 23020 2036
rect 23060 1996 23061 2036
rect 23019 1987 23061 1996
rect 23116 2036 23156 2071
rect 22732 1903 22772 1912
rect 23020 1952 23060 1987
rect 23116 1985 23156 1996
rect 23020 1902 23060 1912
rect 23596 1952 23636 1961
rect 22444 1735 22484 1744
rect 23404 1784 23444 1793
rect 23596 1784 23636 1912
rect 23980 1952 24020 3415
rect 24267 2708 24309 2717
rect 24267 2668 24268 2708
rect 24308 2668 24309 2708
rect 24267 2659 24309 2668
rect 24268 2574 24308 2659
rect 23980 1903 24020 1912
rect 24843 1952 24885 1961
rect 24843 1912 24844 1952
rect 24884 1912 24885 1952
rect 24843 1903 24885 1912
rect 24844 1818 24884 1903
rect 23444 1744 23636 1784
rect 23404 1735 23444 1744
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 25708 1112 25748 3835
rect 25804 3834 25844 3919
rect 25900 3473 25940 7180
rect 26344 7169 26384 7180
rect 26344 7160 26421 7169
rect 26344 7120 26380 7160
rect 26420 7120 26421 7160
rect 26379 7111 26421 7120
rect 30603 5564 30645 5573
rect 30603 5524 30604 5564
rect 30644 5524 30645 5564
rect 30603 5515 30645 5524
rect 28587 5480 28629 5489
rect 28587 5440 28588 5480
rect 28628 5440 28629 5480
rect 28587 5431 28629 5440
rect 26091 5312 26133 5321
rect 26091 5272 26092 5312
rect 26132 5272 26133 5312
rect 26091 5263 26133 5272
rect 27243 5312 27285 5321
rect 27243 5272 27244 5312
rect 27284 5272 27285 5312
rect 27243 5263 27285 5272
rect 26092 5060 26132 5263
rect 26571 5144 26613 5153
rect 26571 5104 26572 5144
rect 26612 5104 26613 5144
rect 26571 5095 26613 5104
rect 26092 5011 26132 5020
rect 25996 4976 26036 4985
rect 25996 4145 26036 4936
rect 26572 4892 26612 5095
rect 26572 4843 26612 4852
rect 26956 4892 26996 4903
rect 26956 4817 26996 4852
rect 26955 4808 26997 4817
rect 26955 4768 26956 4808
rect 26996 4768 26997 4808
rect 26955 4759 26997 4768
rect 26380 4724 26420 4733
rect 26188 4684 26380 4724
rect 25995 4136 26037 4145
rect 25995 4096 25996 4136
rect 26036 4096 26037 4136
rect 25995 4087 26037 4096
rect 26188 3548 26228 4684
rect 26380 4675 26420 4684
rect 26763 4724 26805 4733
rect 26763 4684 26764 4724
rect 26804 4684 26805 4724
rect 26763 4675 26805 4684
rect 26764 4481 26804 4675
rect 26956 4565 26996 4759
rect 27244 4733 27284 5263
rect 28588 4733 28628 5431
rect 30604 5237 30644 5515
rect 30603 5228 30645 5237
rect 30603 5188 30604 5228
rect 30644 5188 30645 5228
rect 30603 5179 30645 5188
rect 30316 4976 30356 4985
rect 27148 4724 27188 4733
rect 27051 4640 27093 4649
rect 27051 4600 27052 4640
rect 27092 4600 27093 4640
rect 27051 4591 27093 4600
rect 26955 4556 26997 4565
rect 26955 4516 26956 4556
rect 26996 4516 26997 4556
rect 26955 4507 26997 4516
rect 27052 4481 27092 4591
rect 26763 4472 26805 4481
rect 26763 4432 26764 4472
rect 26804 4432 26805 4472
rect 26763 4423 26805 4432
rect 27051 4472 27093 4481
rect 27051 4432 27052 4472
rect 27092 4432 27093 4472
rect 27051 4423 27093 4432
rect 27148 4388 27188 4684
rect 27243 4724 27285 4733
rect 27243 4684 27244 4724
rect 27284 4684 27285 4724
rect 27243 4675 27285 4684
rect 28587 4724 28629 4733
rect 28587 4684 28588 4724
rect 28628 4684 28629 4724
rect 28587 4675 28629 4684
rect 29547 4724 29589 4733
rect 29547 4684 29548 4724
rect 29588 4684 29589 4724
rect 29547 4675 29589 4684
rect 28011 4556 28053 4565
rect 28011 4516 28012 4556
rect 28052 4516 28053 4556
rect 28011 4507 28053 4516
rect 27148 4348 27476 4388
rect 27052 4304 27092 4313
rect 27436 4304 27476 4348
rect 27092 4264 27284 4304
rect 27436 4264 27572 4304
rect 27052 4255 27092 4264
rect 26188 3499 26228 3508
rect 26380 4136 26420 4145
rect 25899 3464 25941 3473
rect 25899 3424 25900 3464
rect 25940 3424 25941 3464
rect 25899 3415 25941 3424
rect 26380 2549 26420 4096
rect 26668 4136 26708 4145
rect 26571 3464 26613 3473
rect 26571 3424 26572 3464
rect 26612 3424 26613 3464
rect 26571 3415 26613 3424
rect 26379 2540 26421 2549
rect 26379 2500 26380 2540
rect 26420 2500 26421 2540
rect 26379 2491 26421 2500
rect 25995 2120 26037 2129
rect 25995 2080 25996 2120
rect 26036 2080 26037 2120
rect 25995 2071 26037 2080
rect 25996 1986 26036 2071
rect 26188 1952 26228 1961
rect 25996 1700 26036 1709
rect 25804 1112 25844 1121
rect 25708 1072 25804 1112
rect 25996 1112 26036 1660
rect 26091 1700 26133 1709
rect 26091 1660 26092 1700
rect 26132 1660 26133 1700
rect 26091 1651 26133 1660
rect 26092 1280 26132 1651
rect 26188 1364 26228 1912
rect 26572 1952 26612 3415
rect 26668 2717 26708 4096
rect 26763 4136 26805 4145
rect 26763 4096 26764 4136
rect 26804 4096 26805 4136
rect 26763 4087 26805 4096
rect 27244 4136 27284 4264
rect 27244 4087 27284 4096
rect 27435 4136 27477 4145
rect 27435 4096 27436 4136
rect 27476 4096 27477 4136
rect 27532 4136 27572 4264
rect 27628 4136 27668 4145
rect 27532 4096 27628 4136
rect 27435 4087 27477 4096
rect 26764 4002 26804 4087
rect 27436 3464 27476 4087
rect 27628 3473 27668 4096
rect 27436 3415 27476 3424
rect 27627 3464 27669 3473
rect 27627 3424 27628 3464
rect 27668 3424 27669 3464
rect 27627 3415 27669 3424
rect 26667 2708 26709 2717
rect 26667 2668 26668 2708
rect 26708 2668 26709 2708
rect 26667 2659 26709 2668
rect 27820 2624 27860 2635
rect 27820 2549 27860 2584
rect 27819 2540 27861 2549
rect 27819 2500 27820 2540
rect 27860 2500 27861 2540
rect 27819 2491 27861 2500
rect 26572 1903 26612 1912
rect 27436 1952 27476 1963
rect 27436 1877 27476 1912
rect 27435 1868 27477 1877
rect 27435 1828 27436 1868
rect 27476 1828 27477 1868
rect 27435 1819 27477 1828
rect 28012 1541 28052 4507
rect 28491 4136 28533 4145
rect 28491 4096 28492 4136
rect 28532 4096 28533 4136
rect 28491 4087 28533 4096
rect 28492 4002 28532 4087
rect 28588 3632 28628 4675
rect 29355 3884 29397 3893
rect 29355 3844 29356 3884
rect 29396 3844 29397 3884
rect 29355 3835 29397 3844
rect 28588 3583 28628 3592
rect 28492 2792 28532 2801
rect 28300 2752 28492 2792
rect 28203 2708 28245 2717
rect 28203 2668 28204 2708
rect 28244 2668 28245 2708
rect 28203 2659 28245 2668
rect 28107 2624 28149 2633
rect 28107 2584 28108 2624
rect 28148 2584 28149 2624
rect 28107 2575 28149 2584
rect 28108 2490 28148 2575
rect 28204 2540 28244 2659
rect 28204 2381 28244 2500
rect 28203 2372 28245 2381
rect 28203 2332 28204 2372
rect 28244 2332 28245 2372
rect 28203 2323 28245 2332
rect 28011 1532 28053 1541
rect 28011 1492 28012 1532
rect 28052 1492 28053 1532
rect 28011 1483 28053 1492
rect 26476 1364 26516 1373
rect 26188 1324 26476 1364
rect 26476 1315 26516 1324
rect 26092 1240 26228 1280
rect 26092 1112 26132 1121
rect 25996 1072 26092 1112
rect 25804 1063 25844 1072
rect 26092 1063 26132 1072
rect 26188 1112 26228 1240
rect 26188 1063 26228 1072
rect 28108 1112 28148 1121
rect 28300 1112 28340 2752
rect 28492 2743 28532 2752
rect 29356 2624 29396 3835
rect 29548 3548 29588 4675
rect 29643 4220 29685 4229
rect 29643 4180 29644 4220
rect 29684 4180 29685 4220
rect 29643 4171 29685 4180
rect 29644 3977 29684 4171
rect 30220 4136 30260 4145
rect 30316 4136 30356 4936
rect 30604 4976 30644 5179
rect 30604 4927 30644 4936
rect 30700 4976 30740 4985
rect 30700 4229 30740 4936
rect 30987 4724 31029 4733
rect 30987 4684 30988 4724
rect 31028 4684 31029 4724
rect 30987 4675 31029 4684
rect 30988 4590 31028 4675
rect 30892 4304 30932 4313
rect 30932 4264 31124 4304
rect 30892 4255 30932 4264
rect 30507 4220 30549 4229
rect 30507 4180 30508 4220
rect 30548 4180 30549 4220
rect 30507 4171 30549 4180
rect 30699 4220 30741 4229
rect 30699 4180 30700 4220
rect 30740 4180 30741 4220
rect 30699 4171 30741 4180
rect 30260 4096 30356 4136
rect 30508 4136 30548 4171
rect 29643 3968 29685 3977
rect 29643 3928 29644 3968
rect 29684 3928 29685 3968
rect 29643 3919 29685 3928
rect 29644 3834 29684 3919
rect 30220 3893 30260 4096
rect 30508 4085 30548 4096
rect 30795 4136 30837 4145
rect 30795 4096 30796 4136
rect 30836 4096 30837 4136
rect 30795 4087 30837 4096
rect 31084 4136 31124 4264
rect 31084 4087 31124 4096
rect 31468 4136 31508 4145
rect 30603 4052 30645 4061
rect 30603 4012 30604 4052
rect 30644 4012 30645 4052
rect 30603 4003 30645 4012
rect 30604 3918 30644 4003
rect 30219 3884 30261 3893
rect 30219 3844 30220 3884
rect 30260 3844 30261 3884
rect 30219 3835 30261 3844
rect 29548 3499 29588 3508
rect 29931 3464 29973 3473
rect 29931 3424 29932 3464
rect 29972 3424 29973 3464
rect 29931 3415 29973 3424
rect 30796 3464 30836 4087
rect 31468 3473 31508 4096
rect 31756 3557 31796 7180
rect 33785 7076 33825 7434
rect 33977 7076 34017 7434
rect 34361 7076 34401 7434
rect 34553 7076 34593 7434
rect 34764 7253 34804 7434
rect 34763 7244 34805 7253
rect 34763 7204 34764 7244
rect 34804 7204 34805 7244
rect 34763 7195 34805 7204
rect 34937 7076 34977 7434
rect 35129 7076 35169 7434
rect 35211 7244 35253 7253
rect 35211 7204 35212 7244
rect 35252 7204 35253 7244
rect 35211 7195 35253 7204
rect 33772 7036 33825 7076
rect 33964 7036 34017 7076
rect 34348 7036 34401 7076
rect 34540 7036 34593 7076
rect 34924 7036 34977 7076
rect 35020 7036 35169 7076
rect 33772 5573 33812 7036
rect 33771 5564 33813 5573
rect 33771 5524 33772 5564
rect 33812 5524 33813 5564
rect 33771 5515 33813 5524
rect 32715 5228 32757 5237
rect 32715 5188 32716 5228
rect 32756 5188 32757 5228
rect 32715 5179 32757 5188
rect 31947 5144 31989 5153
rect 31947 5104 31948 5144
rect 31988 5104 31989 5144
rect 31947 5095 31989 5104
rect 32139 5144 32181 5153
rect 32139 5104 32140 5144
rect 32180 5104 32181 5144
rect 32139 5095 32181 5104
rect 32331 5144 32373 5153
rect 32331 5104 32332 5144
rect 32372 5104 32373 5144
rect 32331 5095 32373 5104
rect 32716 5144 32756 5179
rect 31948 5010 31988 5095
rect 32140 5010 32180 5095
rect 32236 4976 32276 4985
rect 32332 4976 32372 5095
rect 32716 5093 32756 5104
rect 32276 4936 32372 4976
rect 32236 4927 32276 4936
rect 32332 4304 32372 4936
rect 32427 4808 32469 4817
rect 32427 4768 32428 4808
rect 32468 4768 32469 4808
rect 32427 4759 32469 4768
rect 32428 4674 32468 4759
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 32332 4264 32468 4304
rect 31947 4220 31989 4229
rect 31947 4180 31948 4220
rect 31988 4180 31989 4220
rect 31947 4171 31989 4180
rect 31948 3632 31988 4171
rect 32235 4136 32277 4145
rect 32235 4096 32236 4136
rect 32276 4096 32277 4136
rect 32235 4087 32277 4096
rect 32332 4136 32372 4145
rect 31948 3583 31988 3592
rect 31755 3548 31797 3557
rect 31755 3508 31756 3548
rect 31796 3508 31797 3548
rect 31755 3499 31797 3508
rect 32236 3473 32276 4087
rect 29932 3330 29972 3415
rect 30028 2792 30068 2801
rect 29356 2575 29396 2584
rect 29452 2752 30028 2792
rect 29452 2372 29492 2752
rect 30028 2743 30068 2752
rect 29164 2332 29492 2372
rect 29644 2624 29684 2633
rect 29164 2036 29204 2332
rect 29644 2213 29684 2584
rect 29739 2624 29781 2633
rect 29739 2584 29740 2624
rect 29780 2584 29781 2624
rect 29739 2575 29781 2584
rect 29740 2490 29780 2575
rect 30507 2372 30549 2381
rect 30507 2332 30508 2372
rect 30548 2332 30549 2372
rect 30507 2323 30549 2332
rect 29643 2204 29685 2213
rect 29643 2164 29644 2204
rect 29684 2164 29685 2204
rect 29643 2155 29685 2164
rect 29164 1987 29204 1996
rect 29548 1952 29588 1961
rect 29355 1868 29397 1877
rect 29355 1828 29356 1868
rect 29396 1828 29397 1868
rect 29355 1819 29397 1828
rect 28588 1700 28628 1711
rect 28588 1625 28628 1660
rect 28587 1616 28629 1625
rect 28587 1576 28588 1616
rect 28628 1576 28629 1616
rect 28587 1567 28629 1576
rect 28491 1532 28533 1541
rect 28491 1492 28492 1532
rect 28532 1492 28533 1532
rect 28491 1483 28533 1492
rect 28148 1072 28340 1112
rect 28492 1112 28532 1483
rect 28108 1063 28148 1072
rect 28492 1063 28532 1072
rect 29356 1112 29396 1819
rect 29548 1541 29588 1912
rect 30412 1952 30452 1963
rect 30412 1877 30452 1912
rect 30411 1868 30453 1877
rect 30411 1828 30412 1868
rect 30452 1828 30453 1868
rect 30411 1819 30453 1828
rect 29547 1532 29589 1541
rect 29547 1492 29548 1532
rect 29588 1492 29589 1532
rect 29547 1483 29589 1492
rect 30508 1364 30548 2323
rect 30796 1961 30836 3424
rect 31467 3464 31509 3473
rect 31467 3424 31468 3464
rect 31508 3424 31509 3464
rect 31467 3415 31509 3424
rect 32235 3464 32277 3473
rect 32235 3424 32236 3464
rect 32276 3424 32277 3464
rect 32235 3415 32277 3424
rect 32236 3330 32276 3415
rect 31563 2708 31605 2717
rect 31563 2668 31564 2708
rect 31604 2668 31605 2708
rect 31563 2659 31605 2668
rect 31467 2540 31509 2549
rect 31467 2500 31468 2540
rect 31508 2500 31509 2540
rect 31467 2491 31509 2500
rect 30795 1952 30837 1961
rect 30795 1912 30796 1952
rect 30836 1912 30837 1952
rect 30795 1903 30837 1912
rect 31468 1868 31508 2491
rect 31564 2120 31604 2659
rect 31755 2624 31797 2633
rect 31755 2584 31756 2624
rect 31796 2584 31797 2624
rect 31755 2575 31797 2584
rect 32235 2624 32277 2633
rect 32235 2584 32236 2624
rect 32276 2584 32277 2624
rect 32235 2575 32277 2584
rect 31756 2490 31796 2575
rect 32236 2490 32276 2575
rect 31660 2456 31700 2465
rect 31660 2129 31700 2416
rect 31947 2456 31989 2465
rect 31947 2416 31948 2456
rect 31988 2416 31989 2456
rect 31947 2407 31989 2416
rect 32139 2456 32181 2465
rect 32139 2416 32140 2456
rect 32180 2416 32181 2456
rect 32139 2407 32181 2416
rect 31948 2322 31988 2407
rect 32140 2322 32180 2407
rect 31564 2071 31604 2080
rect 31659 2120 31701 2129
rect 31659 2080 31660 2120
rect 31700 2080 31701 2120
rect 31659 2071 31701 2080
rect 31756 1952 31796 1961
rect 31468 1828 31604 1868
rect 30508 1315 30548 1324
rect 31564 1205 31604 1828
rect 31756 1364 31796 1912
rect 32140 1952 32180 1961
rect 32140 1541 32180 1912
rect 32332 1877 32372 4096
rect 32428 3632 32468 4264
rect 33964 4061 34004 7036
rect 34348 4229 34388 7036
rect 34540 5480 34580 7036
rect 34924 5489 34964 7036
rect 34444 5440 34580 5480
rect 34923 5480 34965 5489
rect 34923 5440 34924 5480
rect 34964 5440 34965 5480
rect 34444 5144 34484 5440
rect 34923 5431 34965 5440
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 34444 5104 34580 5144
rect 34347 4220 34389 4229
rect 34347 4180 34348 4220
rect 34388 4180 34389 4220
rect 34347 4171 34389 4180
rect 33483 4052 33525 4061
rect 33483 4012 33484 4052
rect 33524 4012 33525 4052
rect 33483 4003 33525 4012
rect 33963 4052 34005 4061
rect 33963 4012 33964 4052
rect 34004 4012 34005 4052
rect 33963 4003 34005 4012
rect 34251 4052 34293 4061
rect 34251 4012 34252 4052
rect 34292 4012 34293 4052
rect 34251 4003 34293 4012
rect 33484 3968 33524 4003
rect 33484 3917 33524 3928
rect 34252 3893 34292 4003
rect 34540 3968 34580 5104
rect 34635 4220 34677 4229
rect 34635 4180 34636 4220
rect 34676 4180 34677 4220
rect 34635 4171 34677 4180
rect 34348 3928 34580 3968
rect 34636 3968 34676 4171
rect 34732 4136 34772 4147
rect 35020 4136 35060 7036
rect 35212 5060 35252 7195
rect 35356 7076 35396 7421
rect 35548 7076 35588 7421
rect 36700 7076 36740 7421
rect 37433 7160 37473 7434
rect 37433 7120 37556 7160
rect 35356 7036 35444 7076
rect 35548 7036 35924 7076
rect 36700 7036 37460 7076
rect 35404 5144 35444 7036
rect 35404 5104 35636 5144
rect 35212 5020 35540 5060
rect 35403 4640 35445 4649
rect 35403 4600 35404 4640
rect 35444 4600 35445 4640
rect 35403 4591 35445 4600
rect 34732 4061 34772 4096
rect 34828 4096 35060 4136
rect 35115 4136 35157 4145
rect 35115 4096 35116 4136
rect 35156 4096 35157 4136
rect 34731 4052 34773 4061
rect 34731 4012 34732 4052
rect 34772 4012 34773 4052
rect 34731 4003 34773 4012
rect 34828 3977 34868 4096
rect 35115 4087 35157 4096
rect 35308 4136 35348 4147
rect 34251 3884 34293 3893
rect 34251 3844 34252 3884
rect 34292 3844 34293 3884
rect 34251 3835 34293 3844
rect 32523 3716 32565 3725
rect 32523 3676 32524 3716
rect 32564 3676 32565 3716
rect 32523 3667 32565 3676
rect 32428 3583 32468 3592
rect 32524 3464 32564 3667
rect 32524 3415 32564 3424
rect 32524 3212 32564 3221
rect 32427 2876 32469 2885
rect 32427 2836 32428 2876
rect 32468 2836 32469 2876
rect 32427 2827 32469 2836
rect 32428 2742 32468 2827
rect 32524 2633 32564 3172
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 34348 2717 34388 3928
rect 34636 3919 34676 3928
rect 34827 3968 34869 3977
rect 34827 3928 34828 3968
rect 34868 3928 34869 3968
rect 34827 3919 34869 3928
rect 34924 3968 34964 3977
rect 34964 3928 35060 3968
rect 34924 3919 34964 3928
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 34827 3632 34869 3641
rect 34827 3592 34828 3632
rect 34868 3592 34869 3632
rect 34827 3583 34869 3592
rect 34828 3464 34868 3583
rect 35020 3473 35060 3928
rect 35116 3725 35156 4087
rect 35308 4061 35348 4096
rect 35307 4052 35349 4061
rect 35307 4012 35308 4052
rect 35348 4012 35349 4052
rect 35307 4003 35349 4012
rect 35212 3968 35252 3977
rect 35212 3800 35252 3928
rect 35212 3760 35348 3800
rect 35115 3716 35157 3725
rect 35115 3676 35116 3716
rect 35156 3676 35157 3716
rect 35115 3667 35157 3676
rect 35115 3548 35157 3557
rect 35115 3508 35116 3548
rect 35156 3508 35157 3548
rect 35115 3499 35157 3508
rect 34828 3415 34868 3424
rect 35019 3464 35061 3473
rect 35019 3424 35020 3464
rect 35060 3424 35061 3464
rect 35019 3415 35061 3424
rect 34923 3380 34965 3389
rect 34923 3340 34924 3380
rect 34964 3340 34965 3380
rect 34923 3331 34965 3340
rect 35116 3380 35156 3499
rect 35211 3464 35253 3473
rect 35211 3424 35212 3464
rect 35252 3424 35253 3464
rect 35211 3415 35253 3424
rect 35116 3331 35156 3340
rect 34924 3246 34964 3331
rect 35212 3330 35252 3415
rect 35308 3389 35348 3760
rect 35307 3380 35349 3389
rect 35307 3340 35308 3380
rect 35348 3340 35349 3380
rect 35307 3331 35349 3340
rect 35020 3296 35060 3305
rect 35020 2900 35060 3256
rect 34828 2860 35060 2900
rect 34347 2708 34389 2717
rect 34347 2668 34348 2708
rect 34388 2668 34389 2708
rect 34347 2659 34389 2668
rect 32523 2624 32565 2633
rect 32523 2584 32524 2624
rect 32564 2584 32565 2624
rect 32523 2575 32565 2584
rect 34828 2624 34868 2860
rect 34923 2792 34965 2801
rect 34923 2752 34924 2792
rect 34964 2752 34965 2792
rect 34923 2743 34965 2752
rect 34924 2658 34964 2743
rect 34828 2575 34868 2584
rect 35020 2624 35060 2633
rect 35060 2584 35348 2624
rect 35020 2575 35060 2584
rect 32715 2456 32757 2465
rect 32715 2416 32716 2456
rect 32756 2416 32757 2456
rect 32715 2407 32757 2416
rect 32427 2204 32469 2213
rect 32427 2164 32428 2204
rect 32468 2164 32469 2204
rect 32427 2155 32469 2164
rect 32331 1868 32373 1877
rect 32331 1828 32332 1868
rect 32372 1828 32373 1868
rect 32331 1819 32373 1828
rect 32139 1532 32181 1541
rect 32139 1492 32140 1532
rect 32180 1492 32181 1532
rect 32139 1483 32181 1492
rect 32236 1364 32276 1373
rect 31756 1324 32236 1364
rect 32236 1315 32276 1324
rect 31563 1196 31605 1205
rect 31563 1156 31564 1196
rect 31604 1156 31605 1196
rect 31563 1147 31605 1156
rect 29356 1063 29396 1072
rect 31564 1112 31604 1147
rect 31564 1063 31604 1072
rect 31851 1112 31893 1121
rect 31851 1072 31852 1112
rect 31892 1072 31893 1112
rect 31851 1063 31893 1072
rect 31948 1112 31988 1121
rect 32428 1112 32468 2155
rect 32716 1457 32756 2407
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 34155 2204 34197 2213
rect 34155 2164 34156 2204
rect 34196 2164 34197 2204
rect 34155 2155 34197 2164
rect 34156 2120 34196 2155
rect 34156 2069 34196 2080
rect 34731 2036 34773 2045
rect 34731 1996 34732 2036
rect 34772 1996 34773 2036
rect 34731 1987 34773 1996
rect 33003 1952 33045 1961
rect 33003 1912 33004 1952
rect 33044 1912 33045 1952
rect 33003 1903 33045 1912
rect 34348 1952 34388 1961
rect 33004 1818 33044 1903
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 32715 1448 32757 1457
rect 32715 1408 32716 1448
rect 32756 1408 32757 1448
rect 32715 1399 32757 1408
rect 34348 1373 34388 1912
rect 34732 1952 34772 1987
rect 34732 1901 34772 1912
rect 35308 1700 35348 2584
rect 35404 2045 35444 4591
rect 35500 3977 35540 5020
rect 35499 3968 35541 3977
rect 35499 3928 35500 3968
rect 35540 3928 35541 3968
rect 35499 3919 35541 3928
rect 35596 2801 35636 5104
rect 35691 4136 35733 4145
rect 35691 4096 35692 4136
rect 35732 4096 35733 4136
rect 35691 4087 35733 4096
rect 35692 3053 35732 4087
rect 35691 3044 35733 3053
rect 35691 3004 35692 3044
rect 35732 3004 35733 3044
rect 35691 2995 35733 3004
rect 35595 2792 35637 2801
rect 35595 2752 35596 2792
rect 35636 2752 35637 2792
rect 35595 2743 35637 2752
rect 35884 2213 35924 7036
rect 37131 6656 37173 6665
rect 37131 6616 37132 6656
rect 37172 6616 37173 6656
rect 37131 6607 37173 6616
rect 36363 6488 36405 6497
rect 36363 6448 36364 6488
rect 36404 6448 36405 6488
rect 36363 6439 36405 6448
rect 35979 5144 36021 5153
rect 35979 5104 35980 5144
rect 36020 5104 36021 5144
rect 35979 5095 36021 5104
rect 35883 2204 35925 2213
rect 35883 2164 35884 2204
rect 35924 2164 35925 2204
rect 35883 2155 35925 2164
rect 35403 2036 35445 2045
rect 35403 1996 35404 2036
rect 35444 1996 35445 2036
rect 35403 1987 35445 1996
rect 35595 1952 35637 1961
rect 35595 1912 35596 1952
rect 35636 1912 35637 1952
rect 35595 1903 35637 1912
rect 35596 1818 35636 1903
rect 35308 1660 35828 1700
rect 35691 1532 35733 1541
rect 35691 1492 35692 1532
rect 35732 1492 35733 1532
rect 35691 1483 35733 1492
rect 34347 1364 34389 1373
rect 34347 1324 34348 1364
rect 34388 1324 34389 1364
rect 34347 1315 34389 1324
rect 34827 1364 34869 1373
rect 34827 1324 34828 1364
rect 34868 1324 34869 1364
rect 34827 1315 34869 1324
rect 34443 1280 34485 1289
rect 34443 1240 34444 1280
rect 34484 1240 34485 1280
rect 34443 1231 34485 1240
rect 34155 1196 34197 1205
rect 34155 1156 34156 1196
rect 34196 1156 34197 1196
rect 34155 1147 34197 1156
rect 31988 1072 32468 1112
rect 34156 1112 34196 1147
rect 31948 1063 31988 1072
rect 31852 978 31892 1063
rect 34156 1061 34196 1072
rect 34444 1112 34484 1231
rect 34828 1230 34868 1315
rect 34444 1063 34484 1072
rect 34539 1112 34581 1121
rect 34539 1072 34540 1112
rect 34580 1072 34581 1112
rect 34539 1063 34581 1072
rect 35692 1112 35732 1483
rect 35788 1364 35828 1660
rect 35980 1541 36020 5095
rect 36364 4304 36404 6439
rect 36939 5144 36981 5153
rect 36939 5104 36940 5144
rect 36980 5104 36981 5144
rect 36939 5095 36981 5104
rect 36940 4976 36980 5095
rect 36940 4927 36980 4936
rect 37132 4976 37172 6607
rect 37227 5396 37269 5405
rect 37227 5356 37228 5396
rect 37268 5356 37269 5396
rect 37227 5347 37269 5356
rect 37132 4927 37172 4936
rect 37036 4724 37076 4733
rect 36364 4255 36404 4264
rect 36460 4684 37036 4724
rect 36268 4136 36308 4145
rect 36268 3716 36308 4096
rect 36460 4136 36500 4684
rect 37036 4675 37076 4684
rect 36460 4087 36500 4096
rect 36268 3676 37172 3716
rect 36939 3464 36981 3473
rect 36939 3424 36940 3464
rect 36980 3424 36981 3464
rect 36939 3415 36981 3424
rect 36940 3330 36980 3415
rect 37035 3380 37077 3389
rect 37035 3340 37036 3380
rect 37076 3340 37077 3380
rect 37035 3331 37077 3340
rect 36747 3296 36789 3305
rect 36747 3256 36748 3296
rect 36788 3256 36789 3296
rect 36747 3247 36789 3256
rect 36459 2624 36501 2633
rect 36459 2584 36460 2624
rect 36500 2584 36501 2624
rect 36459 2575 36501 2584
rect 35979 1532 36021 1541
rect 35979 1492 35980 1532
rect 36020 1492 36021 1532
rect 35979 1483 36021 1492
rect 35788 1315 35828 1324
rect 36460 1205 36500 2575
rect 36651 2540 36693 2549
rect 36651 2500 36652 2540
rect 36692 2500 36693 2540
rect 36651 2491 36693 2500
rect 36555 1784 36597 1793
rect 36555 1744 36556 1784
rect 36596 1744 36597 1784
rect 36555 1735 36597 1744
rect 36459 1196 36501 1205
rect 36459 1156 36460 1196
rect 36500 1156 36501 1196
rect 36459 1147 36501 1156
rect 36556 1121 36596 1735
rect 36652 1532 36692 2491
rect 36748 1793 36788 3247
rect 37036 3246 37076 3331
rect 37132 3296 37172 3676
rect 37228 3380 37268 5347
rect 37323 3548 37365 3557
rect 37323 3508 37324 3548
rect 37364 3508 37365 3548
rect 37323 3499 37365 3508
rect 37324 3464 37364 3499
rect 37324 3413 37364 3424
rect 37228 3331 37268 3340
rect 37132 3247 37172 3256
rect 37420 2900 37460 7036
rect 37516 5741 37556 7120
rect 37625 7076 37665 7434
rect 37612 7036 37665 7076
rect 39580 7076 39620 7421
rect 39737 7076 39777 7434
rect 39929 7076 39969 7434
rect 39580 7036 39668 7076
rect 37515 5732 37557 5741
rect 37515 5692 37516 5732
rect 37556 5692 37557 5732
rect 37515 5683 37557 5692
rect 37612 5405 37652 7036
rect 38859 6572 38901 6581
rect 38859 6532 38860 6572
rect 38900 6532 38901 6572
rect 38859 6523 38901 6532
rect 38667 5732 38709 5741
rect 38667 5692 38668 5732
rect 38708 5692 38709 5732
rect 38667 5683 38709 5692
rect 37611 5396 37653 5405
rect 37611 5356 37612 5396
rect 37652 5356 37653 5396
rect 37611 5347 37653 5356
rect 38571 5144 38613 5153
rect 38571 5104 38572 5144
rect 38612 5104 38613 5144
rect 38571 5095 38613 5104
rect 38668 5144 38708 5683
rect 38763 5144 38805 5153
rect 38668 5104 38764 5144
rect 38804 5104 38805 5144
rect 38572 4976 38612 5095
rect 38572 4178 38612 4936
rect 38668 4892 38708 5104
rect 38763 5095 38805 5104
rect 38860 5060 38900 6523
rect 39243 5312 39285 5321
rect 39243 5272 39244 5312
rect 39284 5272 39285 5312
rect 39243 5263 39285 5272
rect 39244 5060 39284 5263
rect 38860 5020 38996 5060
rect 38956 4976 38996 5020
rect 39244 5011 39284 5020
rect 38668 4843 38708 4852
rect 38860 4892 38900 4901
rect 38763 4808 38805 4817
rect 38763 4768 38764 4808
rect 38804 4768 38805 4808
rect 38763 4759 38805 4768
rect 38667 4724 38709 4733
rect 38667 4684 38668 4724
rect 38708 4684 38709 4724
rect 38667 4675 38709 4684
rect 38668 4304 38708 4675
rect 38764 4674 38804 4759
rect 38668 4255 38708 4264
rect 38572 4138 38708 4178
rect 38571 3968 38613 3977
rect 38571 3928 38572 3968
rect 38612 3928 38613 3968
rect 38571 3919 38613 3928
rect 38475 3716 38517 3725
rect 38475 3676 38476 3716
rect 38516 3676 38517 3716
rect 38475 3667 38517 3676
rect 38284 3464 38324 3473
rect 38284 3137 38324 3424
rect 38379 3380 38421 3389
rect 38379 3340 38380 3380
rect 38420 3340 38421 3380
rect 38379 3331 38421 3340
rect 38380 3246 38420 3331
rect 38476 3296 38516 3667
rect 38572 3380 38612 3919
rect 38668 3464 38708 4138
rect 38668 3415 38708 3424
rect 38860 3389 38900 4852
rect 38956 4733 38996 4936
rect 39148 4976 39188 4985
rect 39148 4817 39188 4936
rect 39340 4976 39380 4985
rect 39340 4817 39380 4936
rect 39147 4808 39189 4817
rect 39147 4768 39148 4808
rect 39188 4768 39189 4808
rect 39147 4759 39189 4768
rect 39339 4808 39381 4817
rect 39339 4768 39340 4808
rect 39380 4768 39381 4808
rect 39339 4759 39381 4768
rect 38955 4724 38997 4733
rect 38955 4684 38956 4724
rect 38996 4684 38997 4724
rect 38955 4675 38997 4684
rect 38572 3331 38612 3340
rect 38859 3380 38901 3389
rect 38859 3340 38860 3380
rect 38900 3340 38901 3380
rect 38859 3331 38901 3340
rect 38476 3247 38516 3256
rect 38283 3128 38325 3137
rect 38283 3088 38284 3128
rect 38324 3088 38325 3128
rect 38283 3079 38325 3088
rect 37420 2860 37556 2900
rect 37516 2717 37556 2860
rect 39051 2876 39093 2885
rect 39051 2836 39052 2876
rect 39092 2836 39093 2876
rect 39051 2827 39093 2836
rect 38955 2792 38997 2801
rect 38955 2752 38956 2792
rect 38996 2752 38997 2792
rect 38955 2743 38997 2752
rect 37515 2708 37557 2717
rect 37515 2668 37516 2708
rect 37556 2668 37557 2708
rect 37515 2659 37557 2668
rect 38667 2624 38709 2633
rect 38667 2584 38668 2624
rect 38708 2584 38709 2624
rect 38667 2575 38709 2584
rect 38956 2624 38996 2743
rect 38956 2575 38996 2584
rect 39052 2624 39092 2827
rect 39340 2792 39380 2801
rect 38668 2490 38708 2575
rect 39052 2549 39092 2584
rect 39244 2752 39340 2792
rect 39051 2540 39093 2549
rect 39051 2500 39052 2540
rect 39092 2500 39093 2540
rect 39051 2491 39093 2500
rect 39052 2460 39092 2491
rect 39147 2204 39189 2213
rect 39147 2164 39148 2204
rect 39188 2164 39189 2204
rect 39147 2155 39189 2164
rect 37323 2036 37365 2045
rect 37323 1996 37324 2036
rect 37364 1996 37365 2036
rect 37323 1987 37365 1996
rect 36940 1952 36980 1961
rect 36747 1784 36789 1793
rect 36747 1744 36748 1784
rect 36788 1744 36789 1784
rect 36747 1735 36789 1744
rect 36748 1650 36788 1735
rect 36843 1532 36885 1541
rect 36652 1492 36788 1532
rect 36651 1196 36693 1205
rect 36651 1156 36652 1196
rect 36692 1156 36693 1196
rect 36651 1147 36693 1156
rect 35692 1063 35732 1072
rect 35884 1112 35924 1121
rect 34540 978 34580 1063
rect 35884 953 35924 1072
rect 36555 1112 36597 1121
rect 36555 1072 36556 1112
rect 36596 1072 36597 1112
rect 36555 1063 36597 1072
rect 36652 1112 36692 1147
rect 36748 1112 36788 1492
rect 36843 1492 36844 1532
rect 36884 1492 36885 1532
rect 36843 1483 36885 1492
rect 36844 1280 36884 1483
rect 36940 1364 36980 1912
rect 37324 1952 37364 1987
rect 37324 1793 37364 1912
rect 38187 1952 38229 1961
rect 38187 1912 38188 1952
rect 38228 1912 38229 1952
rect 38187 1903 38229 1912
rect 38188 1818 38228 1903
rect 39148 1793 39188 2155
rect 37323 1784 37365 1793
rect 37323 1744 37324 1784
rect 37364 1744 37365 1784
rect 37323 1735 37365 1744
rect 39147 1784 39189 1793
rect 39147 1744 39148 1784
rect 39188 1744 39189 1784
rect 39147 1735 39189 1744
rect 37324 1364 37364 1373
rect 36940 1324 37324 1364
rect 37324 1315 37364 1324
rect 36844 1240 37076 1280
rect 36940 1112 36980 1121
rect 36748 1072 36940 1112
rect 36652 1061 36692 1072
rect 36940 1063 36980 1072
rect 37036 1112 37076 1240
rect 37036 1063 37076 1072
rect 38763 1112 38805 1121
rect 38763 1072 38764 1112
rect 38804 1072 38805 1112
rect 38763 1063 38805 1072
rect 39148 1112 39188 1735
rect 39244 1121 39284 2752
rect 39340 2743 39380 2752
rect 39339 2288 39381 2297
rect 39339 2248 39340 2288
rect 39380 2248 39381 2288
rect 39339 2239 39381 2248
rect 39340 2120 39380 2239
rect 39340 2071 39380 2080
rect 39628 1205 39668 7036
rect 39724 7036 39777 7076
rect 39916 7036 39969 7076
rect 40156 7076 40196 7421
rect 40348 7076 40388 7421
rect 40540 7076 40580 7421
rect 40732 7076 40772 7421
rect 40889 7337 40929 7434
rect 40888 7328 40930 7337
rect 40888 7288 40889 7328
rect 40929 7288 40930 7328
rect 40888 7279 40930 7288
rect 43001 7076 43041 7434
rect 46876 7220 46916 7421
rect 47068 7220 47108 7421
rect 47225 7220 47265 7434
rect 47417 7220 47457 7434
rect 47609 7220 47649 7434
rect 74476 7220 74516 22828
rect 46876 7180 46964 7220
rect 47068 7180 47156 7220
rect 40156 7036 40244 7076
rect 40348 7036 40436 7076
rect 40540 7036 40628 7076
rect 40732 7036 40820 7076
rect 39724 1289 39764 7036
rect 39916 3305 39956 7036
rect 40012 4136 40052 4145
rect 40012 3389 40052 4096
rect 40108 4136 40148 4145
rect 40108 3557 40148 4096
rect 40107 3548 40149 3557
rect 40107 3508 40108 3548
rect 40148 3508 40149 3548
rect 40107 3499 40149 3508
rect 40011 3380 40053 3389
rect 40011 3340 40012 3380
rect 40052 3340 40053 3380
rect 40011 3331 40053 3340
rect 39915 3296 39957 3305
rect 39915 3256 39916 3296
rect 39956 3256 39957 3296
rect 39915 3247 39957 3256
rect 40204 2801 40244 7036
rect 40299 4808 40341 4817
rect 40299 4768 40300 4808
rect 40340 4768 40341 4808
rect 40299 4759 40341 4768
rect 40300 3968 40340 4759
rect 40300 3919 40340 3928
rect 40396 2876 40436 7036
rect 40588 2885 40628 7036
rect 40780 6497 40820 7036
rect 42124 7036 43041 7076
rect 40779 6488 40821 6497
rect 40779 6448 40780 6488
rect 40820 6448 40821 6488
rect 40779 6439 40821 6448
rect 41259 5396 41301 5405
rect 41259 5356 41260 5396
rect 41300 5356 41301 5396
rect 41259 5347 41301 5356
rect 41260 4397 41300 5347
rect 40683 4388 40725 4397
rect 40683 4348 40684 4388
rect 40724 4348 40725 4388
rect 40683 4339 40725 4348
rect 41259 4388 41301 4397
rect 41259 4348 41260 4388
rect 41300 4348 41301 4388
rect 41259 4339 41301 4348
rect 40684 4136 40724 4339
rect 40971 4304 41013 4313
rect 40971 4264 40972 4304
rect 41012 4264 41013 4304
rect 40971 4255 41013 4264
rect 41260 4304 41300 4339
rect 40684 4087 40724 4096
rect 40779 4136 40821 4145
rect 40779 4096 40780 4136
rect 40820 4096 40821 4136
rect 40779 4087 40821 4096
rect 40876 4136 40916 4145
rect 40780 4002 40820 4087
rect 40876 3725 40916 4096
rect 40972 4136 41012 4255
rect 41260 4254 41300 4264
rect 40972 4087 41012 4096
rect 41259 4136 41301 4145
rect 41259 4096 41260 4136
rect 41300 4096 41301 4136
rect 41259 4087 41301 4096
rect 40875 3716 40917 3725
rect 40875 3676 40876 3716
rect 40916 3676 40917 3716
rect 40875 3667 40917 3676
rect 41260 3632 41300 4087
rect 41260 3583 41300 3592
rect 40972 3464 41012 3473
rect 40972 3221 41012 3424
rect 41067 3464 41109 3473
rect 41067 3424 41068 3464
rect 41108 3424 41109 3464
rect 41067 3415 41109 3424
rect 41164 3464 41204 3473
rect 41259 3464 41301 3473
rect 41204 3424 41260 3464
rect 41300 3424 41301 3464
rect 41164 3415 41204 3424
rect 41259 3415 41301 3424
rect 41068 3305 41108 3415
rect 41067 3296 41109 3305
rect 41067 3256 41068 3296
rect 41108 3256 41109 3296
rect 41067 3247 41109 3256
rect 40971 3212 41013 3221
rect 40971 3172 40972 3212
rect 41012 3172 41013 3212
rect 40971 3163 41013 3172
rect 40587 2876 40629 2885
rect 40396 2836 40532 2876
rect 40203 2792 40245 2801
rect 40203 2752 40204 2792
rect 40244 2752 40436 2792
rect 40203 2743 40245 2752
rect 40204 2658 40244 2743
rect 40011 2624 40053 2633
rect 40011 2584 40012 2624
rect 40052 2584 40053 2624
rect 40011 2575 40053 2584
rect 40299 2624 40341 2633
rect 40299 2584 40300 2624
rect 40340 2584 40341 2624
rect 40299 2575 40341 2584
rect 40396 2624 40436 2752
rect 40012 2490 40052 2575
rect 40300 2372 40340 2575
rect 40396 2549 40436 2584
rect 40395 2540 40437 2549
rect 40395 2500 40396 2540
rect 40436 2500 40437 2540
rect 40395 2491 40437 2500
rect 40396 2460 40436 2491
rect 40204 2332 40340 2372
rect 39915 2036 39957 2045
rect 39915 1996 39916 2036
rect 39956 1996 39957 2036
rect 39915 1987 39957 1996
rect 39916 1902 39956 1987
rect 40011 1868 40053 1877
rect 40011 1828 40012 1868
rect 40052 1828 40053 1868
rect 40011 1819 40053 1828
rect 39723 1280 39765 1289
rect 39723 1240 39724 1280
rect 39764 1240 39765 1280
rect 39723 1231 39765 1240
rect 39627 1196 39669 1205
rect 39627 1156 39628 1196
rect 39668 1156 39669 1196
rect 39627 1147 39669 1156
rect 39148 1063 39188 1072
rect 39243 1112 39285 1121
rect 39243 1072 39244 1112
rect 39284 1072 39285 1112
rect 39243 1063 39285 1072
rect 40012 1112 40052 1819
rect 40204 1625 40244 2332
rect 40299 2204 40341 2213
rect 40299 2164 40300 2204
rect 40340 2164 40341 2204
rect 40299 2155 40341 2164
rect 40300 1952 40340 2155
rect 40300 1903 40340 1912
rect 40203 1616 40245 1625
rect 40203 1576 40204 1616
rect 40244 1576 40245 1616
rect 40203 1567 40245 1576
rect 40492 1121 40532 2836
rect 40587 2836 40588 2876
rect 40628 2836 40629 2876
rect 40587 2827 40629 2836
rect 41067 2876 41109 2885
rect 41067 2836 41068 2876
rect 41108 2836 41109 2876
rect 41067 2827 41109 2836
rect 40684 2792 40724 2801
rect 40684 2045 40724 2752
rect 40683 2036 40725 2045
rect 40683 1996 40684 2036
rect 40724 1996 40725 2036
rect 40683 1987 40725 1996
rect 41068 1364 41108 2827
rect 42124 2633 42164 7036
rect 42891 6488 42933 6497
rect 42891 6448 42892 6488
rect 42932 6448 42933 6488
rect 42891 6439 42933 6448
rect 42507 4304 42549 4313
rect 42507 4264 42508 4304
rect 42548 4264 42549 4304
rect 42507 4255 42549 4264
rect 42316 4136 42356 4145
rect 42220 4096 42316 4136
rect 42220 3221 42260 4096
rect 42316 4087 42356 4096
rect 42508 4136 42548 4255
rect 42796 4145 42836 4230
rect 42508 4087 42548 4096
rect 42795 4136 42837 4145
rect 42795 4096 42796 4136
rect 42836 4096 42837 4136
rect 42795 4087 42837 4096
rect 42892 4136 42932 6439
rect 45195 4976 45237 4985
rect 45195 4936 45196 4976
rect 45236 4936 45237 4976
rect 45195 4927 45237 4936
rect 43852 4892 43892 4901
rect 43852 4733 43892 4852
rect 45196 4842 45236 4927
rect 46827 4892 46869 4901
rect 46827 4852 46828 4892
rect 46868 4852 46869 4892
rect 46827 4843 46869 4852
rect 46828 4758 46868 4843
rect 43851 4724 43893 4733
rect 43851 4684 43852 4724
rect 43892 4684 43893 4724
rect 43851 4675 43893 4684
rect 43851 4304 43893 4313
rect 46540 4304 46580 4313
rect 43851 4264 43852 4304
rect 43892 4264 43893 4304
rect 43851 4255 43893 4264
rect 46348 4264 46540 4304
rect 42892 4087 42932 4096
rect 43276 4136 43316 4145
rect 42412 3968 42452 3977
rect 42452 3928 43028 3968
rect 42412 3919 42452 3928
rect 42315 3716 42357 3725
rect 42315 3676 42316 3716
rect 42356 3676 42357 3716
rect 42315 3667 42357 3676
rect 42219 3212 42261 3221
rect 42219 3172 42220 3212
rect 42260 3172 42261 3212
rect 42219 3163 42261 3172
rect 42316 2708 42356 3667
rect 42988 3464 43028 3928
rect 43179 3884 43221 3893
rect 43179 3844 43180 3884
rect 43220 3844 43221 3884
rect 43179 3835 43221 3844
rect 43083 3548 43125 3557
rect 43083 3508 43084 3548
rect 43124 3508 43125 3548
rect 43083 3499 43125 3508
rect 42988 3415 43028 3424
rect 43084 3414 43124 3499
rect 43180 3450 43220 3835
rect 43276 3632 43316 4096
rect 43371 4136 43413 4145
rect 43371 4096 43372 4136
rect 43412 4096 43413 4136
rect 43371 4087 43413 4096
rect 43852 4136 43892 4255
rect 43852 4087 43892 4096
rect 44332 4141 44372 4150
rect 43372 4002 43412 4087
rect 43276 3592 43412 3632
rect 43275 3464 43317 3473
rect 43275 3424 43276 3464
rect 43316 3424 43317 3464
rect 43275 3415 43317 3424
rect 43180 3221 43220 3410
rect 43276 3330 43316 3415
rect 43179 3212 43221 3221
rect 43179 3172 43180 3212
rect 43220 3172 43221 3212
rect 43179 3163 43221 3172
rect 42316 2659 42356 2668
rect 42123 2624 42165 2633
rect 42123 2584 42124 2624
rect 42164 2584 42165 2624
rect 42123 2575 42165 2584
rect 42315 2540 42357 2549
rect 42315 2500 42316 2540
rect 42356 2500 42357 2540
rect 42315 2491 42357 2500
rect 42316 2120 42356 2491
rect 42508 2456 42548 2465
rect 42316 2071 42356 2080
rect 42412 2416 42508 2456
rect 41163 1952 41205 1961
rect 41163 1912 41164 1952
rect 41204 1912 41205 1952
rect 41163 1903 41205 1912
rect 41164 1818 41204 1903
rect 42412 1541 42452 2416
rect 42508 2407 42548 2416
rect 42891 2204 42933 2213
rect 42891 2164 42892 2204
rect 42932 2164 42933 2204
rect 42891 2155 42933 2164
rect 42508 1952 42548 1961
rect 42411 1532 42453 1541
rect 42411 1492 42412 1532
rect 42452 1492 42453 1532
rect 42411 1483 42453 1492
rect 41164 1364 41204 1373
rect 41068 1324 41164 1364
rect 41164 1315 41204 1324
rect 40012 1063 40052 1072
rect 40491 1112 40533 1121
rect 40491 1072 40492 1112
rect 40532 1072 40533 1112
rect 40491 1063 40533 1072
rect 42220 1112 42260 1121
rect 42412 1112 42452 1483
rect 42508 1364 42548 1912
rect 42892 1952 42932 2155
rect 42892 1903 42932 1912
rect 43372 1625 43412 3592
rect 43947 3548 43989 3557
rect 43947 3508 43948 3548
rect 43988 3508 43989 3548
rect 43947 3499 43989 3508
rect 43948 3464 43988 3499
rect 43948 3413 43988 3424
rect 44332 3053 44372 4101
rect 45868 4136 45908 4145
rect 44523 3968 44565 3977
rect 44523 3928 44524 3968
rect 44564 3928 44565 3968
rect 44523 3919 44565 3928
rect 44524 3834 44564 3919
rect 45195 3632 45237 3641
rect 45195 3592 45196 3632
rect 45236 3592 45237 3632
rect 45195 3583 45237 3592
rect 45196 3464 45236 3583
rect 45387 3548 45429 3557
rect 45387 3508 45388 3548
rect 45428 3508 45429 3548
rect 45387 3499 45429 3508
rect 45196 3415 45236 3424
rect 45388 3414 45428 3499
rect 44331 3044 44373 3053
rect 44331 3004 44332 3044
rect 44372 3004 44373 3044
rect 44331 2995 44373 3004
rect 45483 2792 45525 2801
rect 45483 2752 45484 2792
rect 45524 2752 45525 2792
rect 45483 2743 45525 2752
rect 43755 1952 43797 1961
rect 43755 1912 43756 1952
rect 43796 1912 43797 1952
rect 43755 1903 43797 1912
rect 45100 1952 45140 1961
rect 43756 1818 43796 1903
rect 44908 1700 44948 1709
rect 43371 1616 43413 1625
rect 43371 1576 43372 1616
rect 43412 1576 43413 1616
rect 43371 1567 43413 1576
rect 44427 1532 44469 1541
rect 44427 1492 44428 1532
rect 44468 1492 44469 1532
rect 44427 1483 44469 1492
rect 42892 1364 42932 1373
rect 42508 1324 42892 1364
rect 42892 1315 42932 1324
rect 42507 1196 42549 1205
rect 42507 1156 42508 1196
rect 42548 1156 42549 1196
rect 42507 1147 42549 1156
rect 42260 1072 42452 1112
rect 42508 1112 42548 1147
rect 42220 1063 42260 1072
rect 38764 978 38804 1063
rect 42508 1061 42548 1072
rect 42603 1112 42645 1121
rect 42603 1072 42604 1112
rect 42644 1072 42645 1112
rect 42603 1063 42645 1072
rect 44428 1112 44468 1483
rect 44811 1280 44853 1289
rect 44811 1240 44812 1280
rect 44852 1240 44853 1280
rect 44811 1231 44853 1240
rect 44428 1063 44468 1072
rect 44715 1112 44757 1121
rect 44715 1072 44716 1112
rect 44756 1072 44757 1112
rect 44715 1063 44757 1072
rect 44812 1112 44852 1231
rect 44908 1121 44948 1660
rect 45100 1364 45140 1912
rect 45484 1952 45524 2743
rect 45868 2717 45908 4096
rect 46155 4136 46197 4145
rect 46155 4096 46156 4136
rect 46196 4096 46197 4136
rect 46155 4087 46197 4096
rect 46156 4002 46196 4087
rect 46251 4052 46293 4061
rect 46251 4012 46252 4052
rect 46292 4012 46293 4052
rect 46251 4003 46293 4012
rect 46252 3918 46292 4003
rect 46059 3548 46101 3557
rect 46059 3508 46060 3548
rect 46100 3508 46101 3548
rect 46059 3499 46101 3508
rect 46252 3548 46292 3557
rect 46348 3548 46388 4264
rect 46540 4255 46580 4264
rect 46292 3508 46388 3548
rect 46252 3499 46292 3508
rect 45867 2708 45909 2717
rect 45867 2668 45868 2708
rect 45908 2668 45909 2708
rect 45867 2659 45909 2668
rect 45484 1903 45524 1912
rect 45868 1541 45908 2659
rect 46060 2624 46100 3499
rect 46924 3473 46964 7180
rect 47116 4985 47156 7180
rect 47212 7180 47265 7220
rect 47404 7180 47457 7220
rect 47596 7180 47649 7220
rect 74092 7180 74516 7220
rect 47115 4976 47157 4985
rect 47115 4936 47116 4976
rect 47156 4936 47157 4976
rect 47115 4927 47157 4936
rect 47020 4724 47060 4733
rect 46636 3464 46676 3473
rect 46347 2876 46389 2885
rect 46347 2836 46348 2876
rect 46388 2836 46389 2876
rect 46347 2827 46389 2836
rect 46060 2575 46100 2584
rect 46348 1952 46388 2827
rect 46636 2801 46676 3424
rect 46923 3464 46965 3473
rect 46923 3424 46924 3464
rect 46964 3424 46965 3464
rect 46923 3415 46965 3424
rect 47020 2801 47060 4684
rect 47212 4229 47252 7180
rect 47404 6068 47444 7180
rect 47308 6028 47444 6068
rect 47211 4220 47253 4229
rect 47211 4180 47212 4220
rect 47252 4180 47253 4220
rect 47211 4171 47253 4180
rect 47116 4136 47156 4145
rect 46635 2792 46677 2801
rect 46635 2752 46636 2792
rect 46676 2752 46677 2792
rect 46635 2743 46677 2752
rect 47019 2792 47061 2801
rect 47019 2752 47020 2792
rect 47060 2752 47061 2792
rect 47019 2743 47061 2752
rect 47116 2717 47156 4096
rect 47308 4061 47348 6028
rect 47596 5984 47636 7180
rect 47404 5944 47636 5984
rect 47404 4145 47444 5944
rect 54603 5732 54645 5741
rect 54603 5692 54604 5732
rect 54644 5692 54645 5732
rect 54603 5683 54645 5692
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 51724 4976 51764 4985
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 47788 4304 47828 4313
rect 47828 4264 48020 4304
rect 47788 4255 47828 4264
rect 47499 4220 47541 4229
rect 47499 4180 47500 4220
rect 47540 4180 47541 4220
rect 47499 4178 47541 4180
rect 47499 4171 47500 4178
rect 47403 4136 47445 4145
rect 47403 4096 47404 4136
rect 47444 4096 47445 4136
rect 47403 4087 47445 4096
rect 47540 4171 47541 4178
rect 47307 4052 47349 4061
rect 47307 4012 47308 4052
rect 47348 4012 47349 4052
rect 47307 4003 47349 4012
rect 47404 4001 47444 4087
rect 47500 4085 47540 4138
rect 47980 4136 48020 4264
rect 50187 4220 50229 4229
rect 50187 4180 50188 4220
rect 50228 4180 50229 4220
rect 50187 4171 50229 4180
rect 50379 4220 50421 4229
rect 50379 4180 50380 4220
rect 50420 4180 50421 4220
rect 50379 4171 50421 4180
rect 47980 4087 48020 4096
rect 48364 4136 48404 4145
rect 48075 3632 48117 3641
rect 48075 3592 48076 3632
rect 48116 3592 48117 3632
rect 48075 3583 48117 3592
rect 47500 3453 47540 3462
rect 47403 3296 47445 3305
rect 47403 3256 47404 3296
rect 47444 3256 47445 3296
rect 47500 3296 47540 3413
rect 47500 3256 47636 3296
rect 47403 3247 47445 3256
rect 47115 2708 47157 2717
rect 47115 2668 47116 2708
rect 47156 2668 47157 2708
rect 47115 2659 47157 2668
rect 46348 1903 46388 1912
rect 47308 2624 47348 2633
rect 47308 1793 47348 2584
rect 47404 2540 47444 3247
rect 47596 2885 47636 3256
rect 47595 2876 47637 2885
rect 47595 2836 47596 2876
rect 47636 2836 47637 2876
rect 47595 2827 47637 2836
rect 47500 2540 47540 2549
rect 47404 2500 47500 2540
rect 47500 2472 47540 2500
rect 47787 2540 47829 2549
rect 47787 2500 47788 2540
rect 47828 2500 47829 2540
rect 47787 2491 47829 2500
rect 47788 1952 47828 2491
rect 47788 1903 47828 1912
rect 48076 1952 48116 3583
rect 48364 2801 48404 4096
rect 48651 4136 48693 4145
rect 48651 4096 48652 4136
rect 48692 4096 48693 4136
rect 48651 4087 48693 4096
rect 49228 4136 49268 4147
rect 48652 3632 48692 4087
rect 49228 4061 49268 4096
rect 49035 4052 49077 4061
rect 49035 4012 49036 4052
rect 49076 4012 49077 4052
rect 49035 4003 49077 4012
rect 49227 4052 49269 4061
rect 49227 4012 49228 4052
rect 49268 4012 49269 4052
rect 49227 4003 49269 4012
rect 49036 3809 49076 4003
rect 49035 3800 49077 3809
rect 49035 3760 49036 3800
rect 49076 3760 49077 3800
rect 49035 3751 49077 3760
rect 48652 3583 48692 3592
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 49228 2885 49268 4003
rect 49419 3968 49461 3977
rect 49419 3928 49420 3968
rect 49460 3928 49461 3968
rect 49419 3919 49461 3928
rect 49420 3809 49460 3919
rect 49419 3800 49461 3809
rect 49419 3760 49420 3800
rect 49460 3760 49461 3800
rect 49419 3751 49461 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 49227 2876 49269 2885
rect 49227 2836 49228 2876
rect 49268 2836 49269 2876
rect 49227 2827 49269 2836
rect 48363 2792 48405 2801
rect 48363 2752 48364 2792
rect 48404 2752 48405 2792
rect 48363 2743 48405 2752
rect 49035 2792 49077 2801
rect 49035 2752 49036 2792
rect 49076 2752 49077 2792
rect 49035 2743 49077 2752
rect 48076 1903 48116 1912
rect 48172 1952 48212 1961
rect 48172 1793 48212 1912
rect 48652 1952 48692 1961
rect 47307 1784 47349 1793
rect 47307 1744 47308 1784
rect 47348 1744 47349 1784
rect 47307 1735 47349 1744
rect 48171 1784 48213 1793
rect 48171 1744 48172 1784
rect 48212 1744 48213 1784
rect 48171 1735 48213 1744
rect 48460 1784 48500 1793
rect 48652 1784 48692 1912
rect 49036 1952 49076 2743
rect 49132 2624 49172 2635
rect 49132 2549 49172 2584
rect 49420 2624 49460 3751
rect 50188 3632 50228 4171
rect 50380 4086 50420 4171
rect 51724 4145 51764 4936
rect 52012 4976 52052 4985
rect 50956 4136 50996 4145
rect 50092 3592 50228 3632
rect 50572 4052 50612 4061
rect 49804 3464 49844 3473
rect 49708 3424 49804 3464
rect 49515 2708 49557 2717
rect 49515 2668 49516 2708
rect 49556 2668 49557 2708
rect 49515 2659 49557 2668
rect 49420 2575 49460 2584
rect 49516 2624 49556 2659
rect 49516 2573 49556 2584
rect 49708 2549 49748 3424
rect 49804 3415 49844 3424
rect 50092 3464 50132 3592
rect 50092 3415 50132 3424
rect 50187 3464 50229 3473
rect 50187 3424 50188 3464
rect 50228 3424 50229 3464
rect 50187 3415 50229 3424
rect 50188 3330 50228 3415
rect 50476 3296 50516 3305
rect 50572 3296 50612 4012
rect 50516 3256 50612 3296
rect 50476 3247 50516 3256
rect 50956 2801 50996 4096
rect 51723 4136 51765 4145
rect 51723 4096 51724 4136
rect 51764 4096 51765 4136
rect 51723 4087 51765 4096
rect 51820 4136 51860 4147
rect 51724 3725 51764 4087
rect 51820 4061 51860 4096
rect 51819 4052 51861 4061
rect 51819 4012 51820 4052
rect 51860 4012 51861 4052
rect 51819 4003 51861 4012
rect 51723 3716 51765 3725
rect 51723 3676 51724 3716
rect 51764 3676 51765 3716
rect 51723 3667 51765 3676
rect 49804 2792 49844 2801
rect 50379 2792 50421 2801
rect 49844 2752 50036 2792
rect 49804 2743 49844 2752
rect 49996 2624 50036 2752
rect 50379 2752 50380 2792
rect 50420 2752 50421 2792
rect 50379 2743 50421 2752
rect 50955 2792 50997 2801
rect 50955 2752 50956 2792
rect 50996 2752 50997 2792
rect 50955 2743 50997 2752
rect 49996 2575 50036 2584
rect 50380 2624 50420 2743
rect 51723 2708 51765 2717
rect 51723 2668 51724 2708
rect 51764 2668 51765 2708
rect 51723 2659 51765 2668
rect 50380 2575 50420 2584
rect 51243 2624 51285 2633
rect 51243 2584 51244 2624
rect 51284 2584 51285 2624
rect 51243 2575 51285 2584
rect 49131 2540 49173 2549
rect 49131 2500 49132 2540
rect 49172 2500 49173 2540
rect 49131 2491 49173 2500
rect 49707 2540 49749 2549
rect 49707 2500 49708 2540
rect 49748 2500 49749 2540
rect 49707 2491 49749 2500
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 51244 2045 51284 2575
rect 51435 2540 51477 2549
rect 51435 2500 51436 2540
rect 51476 2500 51477 2540
rect 51435 2491 51477 2500
rect 49899 2036 49941 2045
rect 49899 1996 49900 2036
rect 49940 1996 49941 2036
rect 49899 1987 49941 1996
rect 51243 2036 51285 2045
rect 51243 1996 51244 2036
rect 51284 1996 51285 2036
rect 51243 1987 51285 1996
rect 49036 1903 49076 1912
rect 49900 1952 49940 1987
rect 49900 1901 49940 1912
rect 48500 1744 48692 1784
rect 51051 1784 51093 1793
rect 51051 1744 51052 1784
rect 51092 1744 51093 1784
rect 48460 1735 48500 1744
rect 51051 1735 51093 1744
rect 47500 1700 47540 1709
rect 45867 1532 45909 1541
rect 45867 1492 45868 1532
rect 45908 1492 45909 1532
rect 45867 1483 45909 1492
rect 45100 1315 45140 1324
rect 47500 1289 47540 1660
rect 51052 1650 51092 1735
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 47499 1280 47541 1289
rect 47499 1240 47500 1280
rect 47540 1240 47541 1280
rect 47499 1231 47541 1240
rect 44812 1063 44852 1072
rect 44907 1112 44949 1121
rect 44907 1072 44908 1112
rect 44948 1072 44949 1112
rect 44907 1063 44949 1072
rect 51436 1112 51476 2491
rect 51436 1063 51476 1072
rect 51724 1112 51764 2659
rect 51820 2633 51860 4003
rect 52012 3473 52052 4936
rect 52107 4976 52149 4985
rect 52107 4936 52108 4976
rect 52148 4936 52149 4976
rect 52107 4927 52149 4936
rect 53643 4976 53685 4985
rect 53643 4936 53644 4976
rect 53684 4936 53685 4976
rect 53643 4927 53685 4936
rect 52108 4842 52148 4927
rect 52396 4724 52436 4733
rect 52300 3548 52340 3557
rect 52396 3548 52436 4684
rect 53644 4397 53684 4927
rect 54604 4901 54644 5683
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 54603 4892 54645 4901
rect 54603 4852 54604 4892
rect 54644 4852 54645 4892
rect 54603 4843 54645 4852
rect 53643 4388 53685 4397
rect 53643 4348 53644 4388
rect 53684 4348 53685 4388
rect 53643 4339 53685 4348
rect 53355 4136 53397 4145
rect 53355 4096 53356 4136
rect 53396 4096 53397 4136
rect 53355 4087 53397 4096
rect 53547 4136 53589 4145
rect 53547 4096 53548 4136
rect 53588 4096 53589 4136
rect 53547 4087 53589 4096
rect 53644 4136 53684 4339
rect 54028 4304 54068 4313
rect 54068 4264 54260 4304
rect 54028 4255 54068 4264
rect 53644 4087 53684 4096
rect 54220 4136 54260 4264
rect 54220 4087 54260 4096
rect 54604 4136 54644 4843
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 54699 4388 54741 4397
rect 54699 4348 54700 4388
rect 54740 4348 54741 4388
rect 54699 4339 54741 4348
rect 54604 4087 54644 4096
rect 52340 3508 52436 3548
rect 52972 3968 53012 3977
rect 52300 3499 52340 3508
rect 52972 3473 53012 3928
rect 53356 3893 53396 4087
rect 53355 3884 53397 3893
rect 53355 3844 53356 3884
rect 53396 3844 53397 3884
rect 53355 3835 53397 3844
rect 52011 3464 52053 3473
rect 52011 3424 52012 3464
rect 52052 3424 52053 3464
rect 52011 3415 52053 3424
rect 52684 3464 52724 3473
rect 52684 2801 52724 3424
rect 52971 3464 53013 3473
rect 53548 3464 53588 4087
rect 53740 4052 53780 4063
rect 53740 3977 53780 4012
rect 53739 3968 53781 3977
rect 53739 3928 53740 3968
rect 53780 3928 53781 3968
rect 53739 3919 53781 3928
rect 54700 3632 54740 4339
rect 55467 4136 55509 4145
rect 55467 4096 55468 4136
rect 55508 4096 55509 4136
rect 55467 4087 55509 4096
rect 55468 4002 55508 4087
rect 56619 3968 56661 3977
rect 56619 3928 56620 3968
rect 56660 3928 56661 3968
rect 56619 3919 56661 3928
rect 56620 3834 56660 3919
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 54700 3583 54740 3592
rect 52971 3424 52972 3464
rect 53012 3424 53013 3464
rect 52971 3415 53013 3424
rect 53260 3424 53548 3464
rect 52299 2792 52341 2801
rect 52299 2752 52300 2792
rect 52340 2752 52341 2792
rect 52299 2743 52341 2752
rect 52683 2792 52725 2801
rect 52683 2752 52684 2792
rect 52724 2752 52725 2792
rect 52683 2743 52725 2752
rect 51819 2624 51861 2633
rect 51819 2584 51820 2624
rect 51860 2584 51861 2624
rect 51819 2575 51861 2584
rect 52012 1952 52052 1961
rect 52300 1952 52340 2743
rect 52395 2708 52437 2717
rect 52395 2668 52396 2708
rect 52436 2668 52437 2708
rect 52395 2659 52437 2668
rect 52396 2574 52436 2659
rect 52396 1952 52436 1961
rect 52052 1912 52148 1952
rect 52300 1912 52396 1952
rect 52012 1903 52052 1912
rect 52108 1364 52148 1912
rect 52396 1903 52436 1912
rect 53260 1952 53300 3424
rect 53548 3415 53588 3424
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 74092 1961 74132 7180
rect 74668 4061 74708 23584
rect 75532 18005 75572 28288
rect 76108 28279 76148 28288
rect 75531 17996 75573 18005
rect 75531 17956 75532 17996
rect 75572 17956 75573 17996
rect 75531 17947 75573 17956
rect 77356 17072 77396 32731
rect 80620 32696 80660 32705
rect 80716 32696 80756 33655
rect 80812 33545 80852 34252
rect 81003 33704 81045 33713
rect 81003 33664 81004 33704
rect 81044 33664 81045 33704
rect 81003 33655 81045 33664
rect 81100 33704 81140 33715
rect 81004 33570 81044 33655
rect 81100 33629 81140 33664
rect 81099 33620 81141 33629
rect 81099 33580 81100 33620
rect 81140 33580 81141 33620
rect 81099 33571 81141 33580
rect 80811 33536 80853 33545
rect 80811 33496 80812 33536
rect 80852 33496 80853 33536
rect 80811 33487 80853 33496
rect 80811 32864 80853 32873
rect 80811 32824 80812 32864
rect 80852 32824 80853 32864
rect 80811 32815 80853 32824
rect 81196 32864 81236 34336
rect 81483 33704 81525 33713
rect 81483 33664 81484 33704
rect 81524 33664 81525 33704
rect 81483 33655 81525 33664
rect 81388 33452 81428 33461
rect 81388 32873 81428 33412
rect 80812 32730 80852 32815
rect 80660 32656 80756 32696
rect 80620 32647 80660 32656
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 80427 31688 80469 31697
rect 80427 31648 80428 31688
rect 80468 31648 80469 31688
rect 80427 31639 80469 31648
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 79947 30596 79989 30605
rect 79947 30556 79948 30596
rect 79988 30556 79989 30596
rect 79947 30547 79989 30556
rect 79948 30462 79988 30547
rect 80140 30428 80180 30437
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 79563 30092 79605 30101
rect 79563 30052 79564 30092
rect 79604 30052 79605 30092
rect 79563 30043 79605 30052
rect 79179 29840 79221 29849
rect 79179 29800 79180 29840
rect 79220 29800 79221 29840
rect 79179 29791 79221 29800
rect 79468 29840 79508 29849
rect 79180 29177 79220 29791
rect 79468 29261 79508 29800
rect 79564 29840 79604 30043
rect 79852 30008 79892 30017
rect 79892 29968 80084 30008
rect 79852 29959 79892 29968
rect 79467 29252 79509 29261
rect 79467 29212 79468 29252
rect 79508 29212 79509 29252
rect 79467 29203 79509 29212
rect 79179 29168 79221 29177
rect 79179 29128 79180 29168
rect 79220 29128 79221 29168
rect 79179 29119 79221 29128
rect 79371 29168 79413 29177
rect 79371 29128 79372 29168
rect 79412 29128 79413 29168
rect 79371 29119 79413 29128
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 78603 28664 78645 28673
rect 78603 28624 78604 28664
rect 78644 28624 78645 28664
rect 78603 28615 78645 28624
rect 77739 17156 77781 17165
rect 77739 17116 77740 17156
rect 77780 17116 77781 17156
rect 77739 17107 77781 17116
rect 77356 17023 77396 17032
rect 77644 17072 77684 17081
rect 77644 7001 77684 17032
rect 77740 17022 77780 17107
rect 78220 17072 78260 17081
rect 78028 16904 78068 16913
rect 78220 16904 78260 17032
rect 78604 17072 78644 28615
rect 79372 28328 79412 29119
rect 79564 28328 79604 29800
rect 80044 29840 80084 29968
rect 80140 29849 80180 30388
rect 80044 29791 80084 29800
rect 80139 29840 80181 29849
rect 80139 29800 80140 29840
rect 80180 29800 80181 29840
rect 80139 29791 80181 29800
rect 80428 29840 80468 31639
rect 80716 31352 80756 32656
rect 80812 32192 80852 32201
rect 80812 31604 80852 32152
rect 81196 32192 81236 32824
rect 81387 32864 81429 32873
rect 81387 32824 81388 32864
rect 81428 32824 81429 32864
rect 81387 32815 81429 32824
rect 81196 31781 81236 32152
rect 81195 31772 81237 31781
rect 81195 31732 81196 31772
rect 81236 31732 81237 31772
rect 81195 31723 81237 31732
rect 81388 31604 81428 31613
rect 80812 31564 81388 31604
rect 81388 31555 81428 31564
rect 80619 30680 80661 30689
rect 80619 30640 80620 30680
rect 80660 30640 80661 30680
rect 80619 30631 80661 30640
rect 80428 29791 80468 29800
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 80427 29252 80469 29261
rect 80427 29212 80428 29252
rect 80468 29212 80469 29252
rect 80427 29203 80469 29212
rect 80043 29168 80085 29177
rect 80043 29128 80044 29168
rect 80084 29128 80085 29168
rect 80043 29119 80085 29128
rect 80332 29168 80372 29177
rect 80044 29034 80084 29119
rect 80332 28841 80372 29128
rect 80428 29118 80468 29203
rect 80331 28832 80373 28841
rect 80331 28792 80332 28832
rect 80372 28792 80373 28832
rect 80331 28783 80373 28792
rect 80523 28832 80565 28841
rect 80523 28792 80524 28832
rect 80564 28792 80565 28832
rect 80523 28783 80565 28792
rect 79755 28580 79797 28589
rect 79755 28540 79756 28580
rect 79796 28540 79797 28580
rect 79755 28531 79797 28540
rect 79660 28328 79700 28337
rect 79564 28288 79660 28328
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 79372 26153 79412 28288
rect 79660 28279 79700 28288
rect 79756 28328 79796 28531
rect 80044 28496 80084 28505
rect 80084 28456 80276 28496
rect 80044 28447 80084 28456
rect 79756 28279 79796 28288
rect 80236 28328 80276 28456
rect 80236 28279 80276 28288
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 80524 27380 80564 28783
rect 80620 28328 80660 30631
rect 80716 30605 80756 31312
rect 81004 31352 81044 31361
rect 80812 30680 80852 30689
rect 80715 30596 80757 30605
rect 80715 30556 80716 30596
rect 80756 30556 80757 30596
rect 80715 30547 80757 30556
rect 80716 29000 80756 29009
rect 80812 29000 80852 30640
rect 81004 29336 81044 31312
rect 81100 31352 81140 31361
rect 81484 31352 81524 33655
rect 81772 33620 81812 35335
rect 82060 34376 82100 34385
rect 82060 34217 82100 34336
rect 82059 34208 82101 34217
rect 82059 34168 82060 34208
rect 82100 34168 82101 34208
rect 82059 34159 82101 34168
rect 83211 34208 83253 34217
rect 83211 34168 83212 34208
rect 83252 34168 83253 34208
rect 83211 34159 83253 34168
rect 81676 33580 81772 33620
rect 81579 32444 81621 32453
rect 81579 32404 81580 32444
rect 81620 32404 81621 32444
rect 81579 32395 81621 32404
rect 81140 31312 81524 31352
rect 81100 31303 81140 31312
rect 81195 30680 81237 30689
rect 81195 30640 81196 30680
rect 81236 30640 81237 30680
rect 81195 30631 81237 30640
rect 81196 30546 81236 30631
rect 81291 29840 81333 29849
rect 81291 29800 81292 29840
rect 81332 29800 81333 29840
rect 81291 29791 81333 29800
rect 81483 29840 81525 29849
rect 81483 29800 81484 29840
rect 81524 29800 81525 29840
rect 81483 29791 81525 29800
rect 81292 29706 81332 29791
rect 81004 29296 81428 29336
rect 81003 29168 81045 29177
rect 81003 29128 81004 29168
rect 81044 29128 81045 29168
rect 81003 29119 81045 29128
rect 81292 29168 81332 29177
rect 81004 29034 81044 29119
rect 80756 28960 80852 29000
rect 80716 28951 80756 28960
rect 81292 28589 81332 29128
rect 81388 29168 81428 29296
rect 81291 28580 81333 28589
rect 81291 28540 81292 28580
rect 81332 28540 81333 28580
rect 81291 28531 81333 28540
rect 80620 27488 80660 28288
rect 81388 27833 81428 29128
rect 81484 28328 81524 29791
rect 81484 28279 81524 28288
rect 81387 27824 81429 27833
rect 81387 27784 81388 27824
rect 81428 27784 81429 27824
rect 81387 27775 81429 27784
rect 80811 27740 80853 27749
rect 80811 27700 80812 27740
rect 80852 27700 80853 27740
rect 80811 27691 80853 27700
rect 80812 27606 80852 27691
rect 81196 27656 81236 27665
rect 81196 27488 81236 27616
rect 80620 27448 81236 27488
rect 80524 27340 80660 27380
rect 80428 26732 80468 26741
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 79371 26144 79413 26153
rect 79371 26104 79372 26144
rect 79412 26104 79413 26144
rect 79371 26095 79413 26104
rect 79947 26144 79989 26153
rect 79947 26104 79948 26144
rect 79988 26104 79989 26144
rect 79947 26095 79989 26104
rect 80235 26144 80277 26153
rect 80235 26104 80236 26144
rect 80276 26104 80277 26144
rect 80235 26095 80277 26104
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 79948 25304 79988 26095
rect 80236 26010 80276 26095
rect 80331 26060 80373 26069
rect 80331 26020 80332 26060
rect 80372 26020 80373 26060
rect 80331 26011 80373 26020
rect 80332 25892 80372 26011
rect 80428 25985 80468 26692
rect 80620 26228 80660 27340
rect 80620 26179 80660 26188
rect 80812 26816 80852 27448
rect 81580 26816 81620 32395
rect 81676 31436 81716 33580
rect 81772 33571 81812 33580
rect 81964 33452 82004 33461
rect 81964 31697 82004 33412
rect 82060 32864 82100 34159
rect 83212 34074 83252 34159
rect 83308 33713 83348 36595
rect 83403 34208 83445 34217
rect 83403 34168 83404 34208
rect 83444 34168 83445 34208
rect 83403 34159 83445 34168
rect 83404 33797 83444 34159
rect 83403 33788 83445 33797
rect 83403 33748 83404 33788
rect 83444 33748 83445 33788
rect 83403 33739 83445 33748
rect 83307 33704 83349 33713
rect 83307 33664 83308 33704
rect 83348 33664 83349 33704
rect 83307 33655 83349 33664
rect 83115 33620 83157 33629
rect 83115 33580 83116 33620
rect 83156 33580 83157 33620
rect 83115 33571 83157 33580
rect 82060 32192 82100 32824
rect 81963 31688 82005 31697
rect 81963 31648 81964 31688
rect 82004 31648 82005 31688
rect 81963 31639 82005 31648
rect 81716 31396 81812 31436
rect 81676 31387 81716 31396
rect 81676 28916 81716 28925
rect 81676 27749 81716 28876
rect 81772 28673 81812 31396
rect 81868 31184 81908 31193
rect 81868 30689 81908 31144
rect 81867 30680 81909 30689
rect 81867 30640 81868 30680
rect 81908 30640 81909 30680
rect 81867 30631 81909 30640
rect 82060 30680 82100 32152
rect 83116 32696 83156 33571
rect 83212 32696 83252 32705
rect 83116 32656 83212 32696
rect 83116 31277 83156 32656
rect 83212 32647 83252 32656
rect 83212 32360 83252 32369
rect 83308 32360 83348 33655
rect 83252 32320 83348 32360
rect 83212 32311 83252 32320
rect 83404 31445 83444 33739
rect 83403 31436 83445 31445
rect 83403 31396 83404 31436
rect 83444 31396 83445 31436
rect 83403 31387 83445 31396
rect 83115 31268 83157 31277
rect 83115 31228 83116 31268
rect 83156 31228 83157 31268
rect 83115 31219 83157 31228
rect 83212 30848 83252 30857
rect 83500 30848 83540 36679
rect 91217 36540 91257 36763
rect 92176 36728 92218 36737
rect 92176 36688 92177 36728
rect 92217 36688 92218 36728
rect 92176 36679 92218 36688
rect 92177 36540 92217 36679
rect 93329 36540 93369 36847
rect 97515 31909 97557 31918
rect 97515 31869 97516 31909
rect 97556 31869 97557 31909
rect 97515 31860 97557 31869
rect 83252 30808 83540 30848
rect 83212 30799 83252 30808
rect 82060 29849 82100 30640
rect 83212 30428 83252 30437
rect 82443 30092 82485 30101
rect 82443 30052 82444 30092
rect 82484 30052 82485 30092
rect 82443 30043 82485 30052
rect 82444 29958 82484 30043
rect 82059 29840 82101 29849
rect 82059 29800 82060 29840
rect 82100 29800 82101 29840
rect 82059 29791 82101 29800
rect 82923 29756 82965 29765
rect 82923 29716 82924 29756
rect 82964 29716 82965 29756
rect 82923 29707 82965 29716
rect 82924 28841 82964 29707
rect 83212 29261 83252 30388
rect 83211 29252 83253 29261
rect 83211 29212 83212 29252
rect 83252 29212 83253 29252
rect 83211 29203 83253 29212
rect 82923 28832 82965 28841
rect 82923 28792 82924 28832
rect 82964 28792 82965 28832
rect 82923 28783 82965 28792
rect 81771 28664 81813 28673
rect 81771 28624 81772 28664
rect 81812 28624 81813 28664
rect 81771 28615 81813 28624
rect 82635 28580 82677 28589
rect 82635 28540 82636 28580
rect 82676 28540 82677 28580
rect 82635 28531 82677 28540
rect 82636 28446 82676 28531
rect 82636 28160 82676 28169
rect 81675 27740 81717 27749
rect 81675 27700 81676 27740
rect 81716 27700 81717 27740
rect 81675 27691 81717 27700
rect 82060 27656 82100 27665
rect 82060 27380 82100 27616
rect 81772 27340 82100 27380
rect 81676 26816 81716 26825
rect 81772 26816 81812 27340
rect 81580 26776 81676 26816
rect 81716 26776 81812 26816
rect 80524 26144 80564 26153
rect 80427 25976 80469 25985
rect 80427 25936 80428 25976
rect 80468 25936 80469 25976
rect 80427 25927 80469 25936
rect 79948 25255 79988 25264
rect 80236 25852 80372 25892
rect 80236 25304 80276 25852
rect 80236 25255 80276 25264
rect 80332 25220 80372 25229
rect 80524 25220 80564 26104
rect 80372 25180 80564 25220
rect 80620 25472 80660 25481
rect 80812 25472 80852 26776
rect 81676 26767 81716 26776
rect 81676 26153 81716 26238
rect 81291 26144 81333 26153
rect 81291 26104 81292 26144
rect 81332 26104 81333 26144
rect 81291 26095 81333 26104
rect 81580 26144 81620 26153
rect 81292 25985 81332 26095
rect 80907 25976 80949 25985
rect 80907 25936 80908 25976
rect 80948 25936 80949 25976
rect 80907 25927 80949 25936
rect 81291 25976 81333 25985
rect 81291 25936 81292 25976
rect 81332 25936 81333 25976
rect 81291 25927 81333 25936
rect 80908 25842 80948 25927
rect 80812 25432 80948 25472
rect 80332 25171 80372 25180
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 80428 24557 80468 25180
rect 80524 24716 80564 24725
rect 80620 24716 80660 25432
rect 80811 25304 80853 25313
rect 80811 25264 80812 25304
rect 80852 25264 80853 25304
rect 80811 25255 80853 25264
rect 80812 25170 80852 25255
rect 80564 24676 80660 24716
rect 80524 24667 80564 24676
rect 80908 24641 80948 25432
rect 81196 25304 81236 25313
rect 81196 24641 81236 25264
rect 80907 24632 80949 24641
rect 80907 24592 80908 24632
rect 80948 24592 80949 24632
rect 80907 24583 80949 24592
rect 81195 24632 81237 24641
rect 81195 24592 81196 24632
rect 81236 24592 81237 24632
rect 81195 24583 81237 24592
rect 80427 24548 80469 24557
rect 80427 24508 80428 24548
rect 80468 24508 80469 24548
rect 80427 24499 80469 24508
rect 80908 24498 80948 24583
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 79467 21608 79509 21617
rect 79467 21568 79468 21608
rect 79508 21568 79509 21608
rect 79467 21559 79509 21568
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 78604 17023 78644 17032
rect 79468 17072 79508 21559
rect 81580 20861 81620 26104
rect 81675 26144 81717 26153
rect 81675 26104 81676 26144
rect 81716 26104 81717 26144
rect 81675 26095 81717 26104
rect 81675 25976 81717 25985
rect 81675 25936 81676 25976
rect 81716 25936 81717 25976
rect 81675 25927 81717 25936
rect 81579 20852 81621 20861
rect 81579 20812 81580 20852
rect 81620 20812 81621 20852
rect 81579 20803 81621 20812
rect 80619 20768 80661 20777
rect 80619 20728 80620 20768
rect 80660 20728 80661 20768
rect 80619 20719 80661 20728
rect 81676 20768 81716 25927
rect 81772 24632 81812 26776
rect 81964 25892 82004 25901
rect 81964 25313 82004 25852
rect 81963 25304 82005 25313
rect 81963 25264 81964 25304
rect 82004 25264 82005 25304
rect 81963 25255 82005 25264
rect 82060 25304 82100 25313
rect 82060 24632 82100 25264
rect 81812 24592 82100 24632
rect 81772 21617 81812 24592
rect 82636 24473 82676 28120
rect 82828 27068 82868 27077
rect 82924 27068 82964 28783
rect 83212 27824 83252 27835
rect 83212 27749 83252 27784
rect 83211 27740 83253 27749
rect 83211 27700 83212 27740
rect 83252 27700 83253 27740
rect 83211 27691 83253 27700
rect 97516 27380 97556 31860
rect 82868 27028 82964 27068
rect 97420 27340 97556 27380
rect 82828 27019 82868 27028
rect 83211 25976 83253 25985
rect 83211 25936 83212 25976
rect 83252 25936 83253 25976
rect 83211 25927 83253 25936
rect 83212 25556 83252 25927
rect 83212 25507 83252 25516
rect 85420 24641 85861 24674
rect 83115 24632 83157 24641
rect 83115 24592 83116 24632
rect 83156 24592 83157 24632
rect 83115 24583 83157 24592
rect 85419 24634 85861 24641
rect 85419 24632 85461 24634
rect 85419 24592 85420 24632
rect 85460 24592 85461 24632
rect 85419 24583 85461 24592
rect 82923 24548 82965 24557
rect 82923 24508 82924 24548
rect 82964 24508 82965 24548
rect 82923 24499 82965 24508
rect 82635 24464 82677 24473
rect 82635 24424 82636 24464
rect 82676 24424 82677 24464
rect 82635 24415 82677 24424
rect 82924 24414 82964 24499
rect 81771 21608 81813 21617
rect 81771 21568 81772 21608
rect 81812 21568 81813 21608
rect 81771 21559 81813 21568
rect 82732 21608 82772 21617
rect 82348 21020 82388 21029
rect 82732 21020 82772 21568
rect 83116 21608 83156 24583
rect 89297 24557 89337 24654
rect 89296 24548 89338 24557
rect 89296 24508 89297 24548
rect 89337 24508 89338 24548
rect 89296 24499 89338 24508
rect 91601 24473 91641 24654
rect 91600 24464 91642 24473
rect 91600 24424 91601 24464
rect 91641 24424 91642 24464
rect 91600 24415 91642 24424
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 83116 21559 83156 21568
rect 83979 21608 84021 21617
rect 83979 21568 83980 21608
rect 84020 21568 84021 21608
rect 83979 21559 84021 21568
rect 83980 21474 84020 21559
rect 97420 21365 97460 27340
rect 85131 21356 85173 21365
rect 85131 21316 85132 21356
rect 85172 21316 85173 21356
rect 85131 21307 85173 21316
rect 97419 21356 97461 21365
rect 97419 21316 97420 21356
rect 97460 21316 97461 21356
rect 97419 21307 97461 21316
rect 82388 20980 82772 21020
rect 82348 20971 82388 20980
rect 85132 20861 85172 21307
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 82059 20852 82101 20861
rect 82059 20812 82060 20852
rect 82100 20812 82101 20852
rect 82059 20803 82101 20812
rect 85131 20852 85173 20861
rect 85131 20812 85132 20852
rect 85172 20812 85173 20852
rect 85131 20803 85173 20812
rect 81676 20719 81716 20728
rect 81963 20768 82005 20777
rect 81963 20728 81964 20768
rect 82004 20728 82005 20768
rect 81963 20719 82005 20728
rect 82060 20768 82100 20803
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 80620 17240 80660 20719
rect 81964 20634 82004 20719
rect 82060 20717 82100 20728
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 82731 20096 82773 20105
rect 82731 20056 82732 20096
rect 82772 20056 82773 20096
rect 82731 20047 82773 20056
rect 98379 20096 98421 20105
rect 98379 20056 98380 20096
rect 98420 20056 98421 20096
rect 98379 20047 98421 20056
rect 80620 17165 80660 17200
rect 80619 17156 80661 17165
rect 80619 17116 80620 17156
rect 80660 17116 80661 17156
rect 80619 17107 80661 17116
rect 80620 17076 80660 17107
rect 79468 17023 79508 17032
rect 78068 16864 78260 16904
rect 78028 16855 78068 16864
rect 80620 16820 80660 16829
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 80620 9269 80660 16780
rect 80619 9260 80661 9269
rect 80619 9220 80620 9260
rect 80660 9220 80661 9260
rect 80619 9211 80661 9220
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 77643 6992 77685 7001
rect 77643 6952 77644 6992
rect 77684 6952 77685 6992
rect 77643 6943 77685 6952
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 80235 6488 80277 6497
rect 80235 6448 80236 6488
rect 80276 6448 80277 6488
rect 80235 6439 80277 6448
rect 78891 6404 78933 6413
rect 78891 6364 78892 6404
rect 78932 6364 78933 6404
rect 78891 6355 78933 6364
rect 78892 6270 78932 6355
rect 80236 6354 80276 6439
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 82732 5153 82772 20047
rect 98380 19962 98420 20047
rect 96843 19928 96885 19937
rect 96843 19888 96844 19928
rect 96884 19888 96885 19928
rect 96843 19879 96885 19888
rect 96844 19794 96884 19879
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 98859 17996 98901 18005
rect 98859 17956 98860 17996
rect 98900 17956 98901 17996
rect 98859 17947 98901 17956
rect 98860 9428 98900 17947
rect 98859 9419 98901 9428
rect 98859 9379 98860 9419
rect 98900 9379 98901 9419
rect 98859 9370 98901 9379
rect 82731 5144 82773 5153
rect 82731 5104 82732 5144
rect 82772 5104 82773 5144
rect 82731 5095 82773 5104
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 74667 4052 74709 4061
rect 74667 4012 74668 4052
rect 74708 4012 74709 4052
rect 74667 4003 74709 4012
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 81963 3128 82005 3137
rect 81963 3088 81964 3128
rect 82004 3088 82005 3128
rect 81963 3079 82005 3088
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 81964 1961 82004 3079
rect 53260 1903 53300 1912
rect 74091 1952 74133 1961
rect 74091 1912 74092 1952
rect 74132 1912 74133 1952
rect 74091 1903 74133 1912
rect 81963 1952 82005 1961
rect 81963 1912 81964 1952
rect 82004 1912 82005 1952
rect 81963 1903 82005 1912
rect 52108 1315 52148 1324
rect 54412 1700 54452 1709
rect 54412 1205 54452 1660
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 90728 1479 90786 1480
rect 90728 1439 90737 1479
rect 90777 1439 90786 1479
rect 90728 1438 90786 1439
rect 91112 1479 91170 1480
rect 91112 1439 91121 1479
rect 91161 1439 91170 1479
rect 91112 1438 91170 1439
rect 91304 1479 91362 1480
rect 91304 1439 91313 1479
rect 91353 1439 91362 1479
rect 91304 1438 91362 1439
rect 90537 1289 90577 1421
rect 90536 1280 90578 1289
rect 90536 1240 90537 1280
rect 90577 1240 90578 1280
rect 90536 1231 90578 1240
rect 51819 1196 51861 1205
rect 51819 1156 51820 1196
rect 51860 1156 51861 1196
rect 51819 1147 51861 1156
rect 54411 1196 54453 1205
rect 54411 1156 54412 1196
rect 54452 1156 54453 1196
rect 54411 1147 54453 1156
rect 51724 1063 51764 1072
rect 51820 1112 51860 1147
rect 42604 978 42644 1063
rect 44716 978 44756 1063
rect 51820 1061 51860 1072
rect 90921 1037 90961 1421
rect 90891 1028 90961 1037
rect 90891 988 90892 1028
rect 90932 988 90961 1028
rect 90891 979 90933 988
rect 35883 944 35925 953
rect 35883 904 35884 944
rect 35924 904 35925 944
rect 35883 895 35925 904
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 21004 38368 21044 38408
rect 22252 38368 22292 38408
rect 844 37948 884 37988
rect 5452 37948 5492 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 652 37528 692 37568
rect 748 37360 788 37400
rect 652 24928 692 24968
rect 652 24088 692 24128
rect 652 23248 692 23288
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 7084 36688 7124 36728
rect 17836 36688 17876 36728
rect 5452 36184 5492 36224
rect 2572 35848 2612 35888
rect 1132 33748 1172 33788
rect 844 25096 884 25136
rect 844 24004 884 24044
rect 652 22408 692 22448
rect 844 21568 884 21608
rect 844 20728 884 20768
rect 844 19888 884 19928
rect 844 19048 884 19088
rect 844 18208 884 18248
rect 844 18040 884 18080
rect 844 17368 884 17408
rect 1324 25096 1364 25136
rect 1132 24004 1172 24044
rect 1228 20056 1268 20096
rect 1228 17872 1268 17912
rect 844 15688 884 15728
rect 652 15436 692 15476
rect 844 14848 884 14888
rect 844 14008 884 14048
rect 748 13168 788 13208
rect 844 12832 884 12872
rect 652 12412 692 12452
rect 1228 16528 1268 16568
rect 1132 16024 1172 16064
rect 1228 14344 1268 14384
rect 1228 13336 1268 13376
rect 652 11740 692 11780
rect 844 11488 884 11528
rect 652 10900 692 10940
rect 844 10732 884 10772
rect 652 10228 692 10268
rect 940 10228 980 10268
rect 844 9808 884 9848
rect 556 5440 596 5480
rect 844 8968 884 9008
rect 748 8128 788 8168
rect 844 7288 884 7328
rect 844 6448 884 6488
rect 844 5608 884 5648
rect 652 4852 692 4892
rect 844 4768 884 4808
rect 844 3928 884 3968
rect 844 3088 884 3128
rect 1228 12328 1268 12368
rect 1228 11740 1268 11780
rect 1132 11572 1172 11612
rect 1132 10900 1172 10940
rect 1036 3508 1076 3548
rect 1228 4180 1268 4220
rect 2092 20812 2132 20852
rect 1612 20728 1652 20768
rect 2284 20056 2324 20096
rect 1996 19552 2036 19592
rect 1612 18628 1652 18668
rect 1612 18040 1652 18080
rect 2476 20644 2516 20684
rect 2476 20056 2516 20096
rect 2476 19300 2516 19340
rect 2380 19216 2420 19256
rect 2284 18460 2324 18500
rect 2092 18376 2132 18416
rect 1804 17872 1844 17912
rect 2284 18208 2324 18248
rect 1900 16024 1940 16064
rect 1612 15352 1652 15392
rect 1804 14848 1844 14888
rect 1516 14680 1556 14720
rect 2188 15352 2228 15392
rect 1996 14344 2036 14384
rect 1612 13840 1652 13880
rect 2188 13840 2228 13880
rect 2092 13168 2132 13208
rect 2188 12832 2228 12872
rect 1900 12244 1940 12284
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4972 34336 5012 34376
rect 4780 34168 4820 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 4396 32068 4436 32108
rect 3820 31900 3860 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 2668 31648 2708 31688
rect 4588 31900 4628 31940
rect 4396 31732 4436 31772
rect 3436 30472 3476 30512
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 3436 27616 3476 27656
rect 5260 34000 5300 34040
rect 4876 31312 4916 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 4492 30724 4532 30764
rect 4780 30640 4820 30680
rect 4876 30556 4916 30596
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 4780 28288 4820 28328
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7084 36016 7124 36056
rect 6412 35848 6452 35888
rect 5548 33832 5588 33872
rect 5260 30724 5300 30764
rect 5356 30640 5396 30680
rect 5164 30472 5204 30512
rect 5068 28288 5108 28328
rect 4972 28036 5012 28076
rect 4876 26692 4916 26732
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3436 25180 3476 25220
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 3436 23080 3476 23120
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 4780 24676 4820 24716
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 3724 22324 3764 22364
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 4396 23080 4436 23120
rect 3916 22324 3956 22364
rect 4204 22324 4244 22364
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 3340 20728 3380 20768
rect 3916 20812 3956 20852
rect 3820 20728 3860 20768
rect 4108 22240 4148 22280
rect 4588 22240 4628 22280
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 4780 20812 4820 20852
rect 4012 20644 4052 20684
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 4300 20140 4340 20180
rect 4108 20056 4148 20096
rect 3532 19888 3572 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4588 19888 4628 19928
rect 3628 19552 3668 19592
rect 4204 19552 4244 19592
rect 3532 19468 3572 19508
rect 3436 19384 3476 19424
rect 2668 19300 2708 19340
rect 2668 18460 2708 18500
rect 2764 18208 2804 18248
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 2476 17116 2516 17156
rect 1804 11656 1844 11696
rect 2092 11656 2132 11696
rect 1900 11572 1940 11612
rect 1996 10984 2036 11024
rect 2188 10648 2228 10688
rect 1900 9808 1940 9848
rect 2476 10648 2516 10688
rect 2380 9808 2420 9848
rect 2284 6616 2324 6656
rect 1324 3676 1364 3716
rect 1132 2836 1172 2876
rect 3724 18628 3764 18668
rect 3820 18376 3860 18416
rect 3436 17032 3476 17072
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 2860 15940 2900 15980
rect 3436 15520 3476 15560
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 3628 14680 3668 14720
rect 3532 14344 3572 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 2956 13336 2996 13376
rect 2764 12412 2804 12452
rect 2572 6868 2612 6908
rect 3436 13252 3476 13292
rect 3436 12496 3476 12536
rect 3244 12244 3284 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3436 10060 3476 10100
rect 3628 11572 3668 11612
rect 3628 10984 3668 11024
rect 3628 10228 3668 10268
rect 3532 9976 3572 10016
rect 3820 17116 3860 17156
rect 4684 19384 4724 19424
rect 4396 19216 4436 19256
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 4300 18628 4340 18668
rect 4012 17956 4052 17996
rect 4108 17872 4148 17912
rect 4876 19300 4916 19340
rect 4492 17956 4532 17996
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4012 16864 4052 16904
rect 4012 16024 4052 16064
rect 4012 14848 4052 14888
rect 5164 27616 5204 27656
rect 5260 27364 5300 27404
rect 5164 26692 5204 26732
rect 5068 25180 5108 25220
rect 5068 19468 5108 19508
rect 4684 16696 4724 16736
rect 4588 16192 4628 16232
rect 4780 15940 4820 15980
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4108 14680 4148 14720
rect 4684 14680 4724 14720
rect 3916 14344 3956 14384
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3820 13336 3860 13376
rect 4012 14008 4052 14048
rect 4012 11908 4052 11948
rect 3916 11824 3956 11864
rect 3916 11572 3956 11612
rect 3820 10984 3860 11024
rect 3820 10732 3860 10772
rect 4780 14008 4820 14048
rect 4300 13252 4340 13292
rect 4972 17032 5012 17072
rect 5068 16192 5108 16232
rect 4972 15520 5012 15560
rect 5068 14680 5108 14720
rect 4684 13168 4724 13208
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 4204 12748 4244 12788
rect 4588 12496 4628 12536
rect 4300 11824 4340 11864
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 4972 12496 5012 12536
rect 5644 33076 5684 33116
rect 5644 32068 5684 32108
rect 5740 31648 5780 31688
rect 5932 31480 5972 31520
rect 5836 31312 5876 31352
rect 5740 30556 5780 30596
rect 5548 28036 5588 28076
rect 5836 27364 5876 27404
rect 6028 25936 6068 25976
rect 5836 24676 5876 24716
rect 5932 22240 5972 22280
rect 5836 21904 5876 21944
rect 5356 21484 5396 21524
rect 5836 21484 5876 21524
rect 5932 20896 5972 20936
rect 5356 20644 5396 20684
rect 5260 20140 5300 20180
rect 6412 19300 6452 19340
rect 6028 19216 6068 19256
rect 5356 18880 5396 18920
rect 5836 16696 5876 16736
rect 5836 16528 5876 16568
rect 5836 16192 5876 16232
rect 5836 14008 5876 14048
rect 5740 12748 5780 12788
rect 5164 11908 5204 11948
rect 4972 11656 5012 11696
rect 4780 10984 4820 11024
rect 4108 10732 4148 10772
rect 3724 9556 3764 9596
rect 3628 9472 3668 9512
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 3436 7960 3476 8000
rect 4012 9556 4052 9596
rect 4204 10060 4244 10100
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4396 9472 4436 9512
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 5836 12664 5876 12704
rect 5836 12328 5876 12368
rect 5836 11824 5876 11864
rect 5836 10228 5876 10268
rect 5068 7960 5108 8000
rect 4780 7708 4820 7748
rect 4684 7120 4724 7160
rect 5740 7708 5780 7748
rect 4012 7036 4052 7076
rect 4396 7036 4436 7076
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 5932 6784 5972 6824
rect 6412 6532 6452 6572
rect 2764 6448 2804 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 2476 5356 2516 5396
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 13708 35848 13748 35888
rect 12268 35092 12308 35132
rect 12460 35092 12500 35132
rect 7372 34504 7412 34544
rect 7372 34336 7412 34376
rect 10924 34000 10964 34040
rect 8236 33916 8276 33956
rect 7852 31564 7892 31604
rect 7756 20812 7796 20852
rect 7756 16696 7796 16736
rect 7756 16360 7796 16400
rect 7948 16360 7988 16400
rect 7948 6952 7988 6992
rect 7852 5776 7892 5816
rect 7084 5104 7124 5144
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 8332 32488 8372 32528
rect 8236 4012 8276 4052
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 2380 2752 2420 2792
rect 940 2416 980 2456
rect 844 2248 884 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 11308 34252 11348 34292
rect 13036 34168 13076 34208
rect 14188 35176 14228 35216
rect 15532 35848 15572 35888
rect 14572 35764 14612 35804
rect 14668 35596 14708 35636
rect 16492 35848 16532 35888
rect 17452 35848 17492 35888
rect 17356 35764 17396 35804
rect 15628 35596 15668 35636
rect 16876 35596 16916 35636
rect 14668 35092 14708 35132
rect 13804 34924 13844 34964
rect 14476 34924 14516 34964
rect 13708 34252 13748 34292
rect 14188 34252 14228 34292
rect 15628 35176 15668 35216
rect 16684 34924 16724 34964
rect 15244 34168 15284 34208
rect 15532 34168 15572 34208
rect 13420 34000 13460 34040
rect 16012 34336 16052 34376
rect 17068 34504 17108 34544
rect 17644 35680 17684 35720
rect 18892 36688 18932 36728
rect 19084 36688 19124 36728
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 19372 37276 19412 37316
rect 20140 37276 20180 37316
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 19372 36772 19412 36812
rect 19180 36604 19220 36644
rect 18316 35848 18356 35888
rect 19372 36436 19412 36476
rect 18124 35512 18164 35552
rect 19756 35848 19796 35888
rect 20236 36604 20276 36644
rect 19948 35764 19988 35804
rect 19372 35512 19412 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 18700 35344 18740 35384
rect 18316 35176 18356 35216
rect 18604 35008 18644 35048
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 19852 35176 19892 35216
rect 19564 34840 19604 34880
rect 19852 34504 19892 34544
rect 18892 34336 18932 34376
rect 19372 34336 19412 34376
rect 20620 37192 20660 37232
rect 20908 37108 20948 37148
rect 20428 36772 20468 36812
rect 20716 36604 20756 36644
rect 21388 37360 21428 37400
rect 21292 37276 21332 37316
rect 21772 37276 21812 37316
rect 21484 37108 21524 37148
rect 21772 37108 21812 37148
rect 21388 36688 21428 36728
rect 21004 36436 21044 36476
rect 20620 35764 20660 35804
rect 21196 35848 21236 35888
rect 20812 35680 20852 35720
rect 21004 35680 21044 35720
rect 21292 35764 21332 35804
rect 20140 35008 20180 35048
rect 20140 34588 20180 34628
rect 20044 34336 20084 34376
rect 18796 34168 18836 34208
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 20812 34504 20852 34544
rect 21292 35008 21332 35048
rect 21292 34840 21332 34880
rect 21580 37024 21620 37064
rect 21580 36688 21620 36728
rect 21772 36688 21812 36728
rect 21676 36268 21716 36308
rect 22540 37024 22580 37064
rect 22924 36856 22964 36896
rect 21964 36268 22004 36308
rect 22348 36688 22388 36728
rect 23020 36688 23060 36728
rect 22444 36436 22484 36476
rect 23500 37024 23540 37064
rect 23308 36940 23348 36980
rect 23308 36772 23348 36812
rect 23500 36520 23540 36560
rect 23212 36268 23252 36308
rect 22828 35848 22868 35888
rect 23116 35848 23156 35888
rect 23788 37360 23828 37400
rect 23980 37360 24020 37400
rect 23692 36604 23732 36644
rect 23692 36436 23732 36476
rect 23884 36688 23924 36728
rect 23980 36520 24020 36560
rect 23884 36268 23924 36308
rect 23596 35512 23636 35552
rect 21580 35344 21620 35384
rect 23404 34588 23444 34628
rect 21388 34504 21428 34544
rect 22252 34504 22292 34544
rect 20236 31900 20276 31940
rect 25900 37444 25940 37484
rect 24364 37024 24404 37064
rect 25228 36940 25268 36980
rect 24460 36856 24500 36896
rect 24844 36856 24884 36896
rect 24652 36772 24692 36812
rect 25324 36856 25364 36896
rect 26380 37276 26420 37316
rect 26668 37276 26708 37316
rect 25228 36688 25268 36728
rect 25516 36604 25556 36644
rect 26092 36688 26132 36728
rect 25900 36520 25940 36560
rect 25516 36352 25556 36392
rect 26188 36352 26228 36392
rect 26860 38200 26900 38240
rect 26860 37444 26900 37484
rect 26476 36940 26516 36980
rect 26668 36856 26708 36896
rect 27052 37360 27092 37400
rect 28876 38368 28916 38408
rect 29260 38368 29300 38408
rect 27340 38200 27380 38240
rect 28492 38200 28532 38240
rect 26956 37108 26996 37148
rect 26764 36772 26804 36812
rect 26860 36688 26900 36728
rect 26572 36604 26612 36644
rect 25228 36268 25268 36308
rect 25996 36268 26036 36308
rect 26380 36268 26420 36308
rect 25900 35848 25940 35888
rect 24268 35764 24308 35804
rect 24172 35596 24212 35636
rect 25612 35344 25652 35384
rect 24460 35176 24500 35216
rect 25708 35176 25748 35216
rect 23980 34924 24020 34964
rect 24076 34336 24116 34376
rect 25900 34504 25940 34544
rect 25036 34420 25076 34460
rect 25996 34420 26036 34460
rect 24844 33916 24884 33956
rect 24172 33748 24212 33788
rect 27148 36940 27188 36980
rect 27436 38116 27476 38156
rect 27340 36688 27380 36728
rect 28876 37444 28916 37484
rect 28780 37276 28820 37316
rect 27532 36688 27572 36728
rect 27916 36772 27956 36812
rect 27628 36604 27668 36644
rect 28012 36604 28052 36644
rect 27052 36520 27092 36560
rect 27724 36520 27764 36560
rect 27052 36352 27092 36392
rect 26572 34672 26612 34712
rect 28780 36856 28820 36896
rect 29452 38200 29492 38240
rect 31468 38200 31508 38240
rect 29452 37360 29492 37400
rect 29452 36856 29492 36896
rect 30316 36856 30356 36896
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 32332 37360 32372 37400
rect 33676 37360 33716 37400
rect 36652 37360 36692 37400
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 30316 36688 30356 36728
rect 31180 36688 31220 36728
rect 28684 36520 28724 36560
rect 27532 35680 27572 35720
rect 30124 35680 30164 35720
rect 27244 35344 27284 35384
rect 28396 35428 28436 35468
rect 29260 35428 29300 35468
rect 27724 35344 27764 35384
rect 28012 35344 28052 35384
rect 28972 35344 29012 35384
rect 26860 34504 26900 34544
rect 27052 34336 27092 34376
rect 28396 34420 28436 34460
rect 29356 35344 29396 35384
rect 28972 34588 29012 34628
rect 29260 34504 29300 34544
rect 28780 34336 28820 34376
rect 29356 34420 29396 34460
rect 29836 34420 29876 34460
rect 29548 34336 29588 34376
rect 26092 32488 26132 32528
rect 17356 31648 17396 31688
rect 18041 31648 18081 31688
rect 18268 31648 18308 31688
rect 18700 31648 18740 31688
rect 11212 31480 11252 31520
rect 15161 31480 15201 31520
rect 15916 31480 15956 31520
rect 16313 31340 16353 31380
rect 30220 35512 30260 35552
rect 31276 35848 31316 35888
rect 31564 35848 31604 35888
rect 31468 35764 31508 35804
rect 31180 34588 31220 34628
rect 31084 34504 31124 34544
rect 30412 34420 30452 34460
rect 31948 35764 31988 35804
rect 33676 36688 33716 36728
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 34444 36016 34484 36056
rect 35116 35932 35156 35972
rect 34828 35764 34868 35804
rect 32524 35512 32564 35552
rect 32716 35512 32756 35552
rect 31852 35344 31892 35384
rect 32236 35344 32276 35384
rect 31564 34168 31604 34208
rect 31660 34084 31700 34124
rect 35020 35596 35060 35636
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 33868 35260 33908 35300
rect 33484 35176 33524 35216
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 33388 34504 33428 34544
rect 32908 34336 32948 34376
rect 33004 34168 33044 34208
rect 32908 33916 32948 33956
rect 34636 35176 34676 35216
rect 35308 35764 35348 35804
rect 35500 35680 35540 35720
rect 37804 37276 37844 37316
rect 38764 38200 38804 38240
rect 39820 38200 39860 38240
rect 38476 37192 38516 37232
rect 38188 36856 38228 36896
rect 38860 36856 38900 36896
rect 38572 36688 38612 36728
rect 38476 36100 38516 36140
rect 38380 35932 38420 35972
rect 35788 35764 35828 35804
rect 37900 35764 37940 35804
rect 38188 35764 38228 35804
rect 37804 35680 37844 35720
rect 35788 35596 35828 35636
rect 35500 35176 35540 35216
rect 35884 35176 35924 35216
rect 33868 34672 33908 34712
rect 37612 35008 37652 35048
rect 35884 34504 35924 34544
rect 34444 34084 34484 34124
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 37324 34588 37364 34628
rect 35212 34168 35252 34208
rect 37036 34168 37076 34208
rect 35116 33916 35156 33956
rect 38476 35596 38516 35636
rect 38476 35260 38516 35300
rect 38092 35008 38132 35048
rect 38092 34504 38132 34544
rect 38668 35932 38708 35972
rect 39052 37360 39092 37400
rect 39148 37276 39188 37316
rect 39724 36688 39764 36728
rect 39148 36100 39188 36140
rect 38956 35848 38996 35888
rect 38764 35764 38804 35804
rect 40588 37192 40628 37232
rect 41068 37192 41108 37232
rect 40300 35932 40340 35972
rect 39916 35848 39956 35888
rect 40108 35848 40148 35888
rect 40396 35848 40436 35888
rect 39532 35764 39572 35804
rect 39052 35008 39092 35048
rect 41068 36772 41108 36812
rect 41452 38200 41492 38240
rect 43468 38200 43508 38240
rect 41356 37192 41396 37232
rect 41452 36856 41492 36896
rect 41644 37192 41684 37232
rect 42220 37192 42260 37232
rect 41740 36772 41780 36812
rect 40876 35848 40916 35888
rect 41164 35344 41204 35384
rect 39436 34672 39476 34712
rect 41836 35848 41876 35888
rect 42124 35848 42164 35888
rect 42796 37108 42836 37148
rect 42508 36856 42548 36896
rect 42316 36688 42356 36728
rect 41644 35764 41684 35804
rect 41548 35428 41588 35468
rect 42028 35260 42068 35300
rect 41356 34924 41396 34964
rect 41356 34756 41396 34796
rect 41260 34084 41300 34124
rect 41644 34084 41684 34124
rect 39148 33916 39188 33956
rect 39724 33916 39764 33956
rect 37612 33832 37652 33872
rect 42316 34168 42356 34208
rect 42220 33664 42260 33704
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 44524 37192 44564 37232
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 43852 35848 43892 35888
rect 45292 36184 45332 36224
rect 43564 35596 43604 35636
rect 43948 35596 43988 35636
rect 43852 35512 43892 35552
rect 43372 35260 43412 35300
rect 44428 35344 44468 35384
rect 42796 35008 42836 35048
rect 42892 34672 42932 34712
rect 42700 34000 42740 34040
rect 43468 34672 43508 34712
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 47980 36016 48020 36056
rect 45484 35344 45524 35384
rect 47020 35680 47060 35720
rect 46828 35512 46868 35552
rect 45292 35260 45332 35300
rect 45676 35260 45716 35300
rect 43756 35008 43796 35048
rect 44812 35008 44852 35048
rect 47596 35428 47636 35468
rect 48268 35428 48308 35468
rect 46924 35092 46964 35132
rect 46540 34924 46580 34964
rect 46732 34924 46772 34964
rect 43372 34504 43412 34544
rect 46444 34504 46484 34544
rect 43564 34168 43604 34208
rect 43756 34168 43796 34208
rect 46924 34840 46964 34880
rect 46444 34000 46484 34040
rect 45196 33832 45236 33872
rect 43180 33664 43220 33704
rect 46828 33580 46868 33620
rect 47884 35092 47924 35132
rect 47212 34588 47252 34628
rect 47788 34924 47828 34964
rect 48076 34840 48116 34880
rect 47980 34588 48020 34628
rect 47500 33580 47540 33620
rect 47116 33496 47156 33536
rect 41836 33412 41876 33452
rect 42508 33412 42548 33452
rect 47500 33328 47540 33368
rect 41740 32824 41780 32864
rect 33772 32404 33812 32444
rect 49228 35260 49268 35300
rect 48364 35092 48404 35132
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 49228 34756 49268 34796
rect 48652 34588 48692 34628
rect 48844 34504 48884 34544
rect 49132 34504 49172 34544
rect 48844 33580 48884 33620
rect 48940 33496 48980 33536
rect 49132 33496 49172 33536
rect 48268 32740 48308 32780
rect 49132 33328 49172 33368
rect 50188 35680 50228 35720
rect 52300 35680 52340 35720
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 50188 34924 50228 34964
rect 50380 34924 50420 34964
rect 49804 34504 49844 34544
rect 50956 35092 50996 35132
rect 52684 35764 52724 35804
rect 53548 35764 53588 35804
rect 53260 35680 53300 35720
rect 53548 35092 53588 35132
rect 51916 34756 51956 34796
rect 51820 34672 51860 34712
rect 50380 34504 50420 34544
rect 51532 34504 51572 34544
rect 52780 34504 52820 34544
rect 51532 34168 51572 34208
rect 52492 34168 52532 34208
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 50380 34000 50420 34040
rect 53740 34924 53780 34964
rect 53644 34672 53684 34712
rect 53548 34084 53588 34124
rect 52972 34000 53012 34040
rect 52492 33580 52532 33620
rect 49516 33076 49556 33116
rect 65260 35932 65300 35972
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 70636 37360 70676 37400
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 93329 36856 93369 36896
rect 91217 36772 91257 36812
rect 74092 36688 74132 36728
rect 83500 36688 83540 36728
rect 65932 35848 65972 35888
rect 70348 35848 70388 35888
rect 72268 35848 72308 35888
rect 73900 35848 73940 35888
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 65260 35512 65300 35552
rect 55564 34924 55604 34964
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 54412 34672 54452 34712
rect 55372 34672 55412 34712
rect 72652 35176 72692 35216
rect 61516 34504 61556 34544
rect 65932 34504 65972 34544
rect 54508 34084 54548 34124
rect 53836 34000 53876 34040
rect 53836 33328 53876 33368
rect 56524 34000 56564 34040
rect 64684 34336 64724 34376
rect 66892 34168 66932 34208
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 63340 33076 63380 33116
rect 63340 32572 63380 32612
rect 55372 32404 55412 32444
rect 62476 32404 62516 32444
rect 83308 36604 83348 36644
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 79564 35596 79604 35636
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 81772 35344 81812 35384
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 79564 33748 79604 33788
rect 80140 33748 80180 33788
rect 79756 33664 79796 33704
rect 80716 33664 80756 33704
rect 80044 33580 80084 33620
rect 80428 33496 80468 33536
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 77356 32740 77396 32780
rect 80428 32740 80468 32780
rect 76108 32572 76148 32612
rect 16588 7120 16628 7160
rect 15820 7036 15860 7076
rect 12364 5356 12404 5396
rect 12364 5104 12404 5144
rect 16396 6616 16436 6656
rect 16588 6616 16628 6656
rect 17164 6616 17204 6656
rect 15820 4600 15860 4640
rect 16876 5776 16916 5816
rect 16012 4348 16052 4388
rect 16588 4600 16628 4640
rect 16396 4180 16436 4220
rect 16972 5272 17012 5312
rect 19948 6616 19988 6656
rect 19948 5944 19988 5984
rect 18412 5272 18452 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 17260 4768 17300 4808
rect 18700 4768 18740 4808
rect 17260 4348 17300 4388
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 17836 4180 17876 4220
rect 20236 4600 20276 4640
rect 18700 4096 18740 4136
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 20428 4180 20468 4220
rect 21196 6532 21236 6572
rect 20620 4180 20660 4220
rect 20524 3928 20564 3968
rect 20428 3424 20468 3464
rect 21772 5272 21812 5312
rect 21580 4684 21620 4724
rect 21388 4600 21428 4640
rect 21292 4096 21332 4136
rect 21676 4180 21716 4220
rect 20044 3256 20084 3296
rect 20908 3256 20948 3296
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 21484 2500 21524 2540
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 22060 4684 22100 4724
rect 23212 5272 23252 5312
rect 23404 4684 23444 4724
rect 22732 4600 22772 4640
rect 22444 4180 22484 4220
rect 21964 3424 22004 3464
rect 22252 3424 22292 3464
rect 21772 2080 21812 2120
rect 8332 1912 8372 1952
rect 22156 1996 22196 2036
rect 22828 4096 22868 4136
rect 23020 2668 23060 2708
rect 22732 2080 22772 2120
rect 23500 2668 23540 2708
rect 23788 6784 23828 6824
rect 25708 6868 25748 6908
rect 23980 5944 24020 5984
rect 23980 5272 24020 5312
rect 24364 5272 24404 5312
rect 24076 4600 24116 4640
rect 25420 4768 25460 4808
rect 24748 4684 24788 4724
rect 25228 4684 25268 4724
rect 25708 4600 25748 4640
rect 24652 4096 24692 4136
rect 24460 3928 24500 3968
rect 25804 3928 25844 3968
rect 25708 3844 25748 3884
rect 23788 3424 23828 3464
rect 23980 3424 24020 3464
rect 23116 2080 23156 2120
rect 23596 2080 23636 2120
rect 23020 1996 23060 2036
rect 24268 2668 24308 2708
rect 24844 1912 24884 1952
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 26380 7120 26420 7160
rect 30604 5524 30644 5564
rect 28588 5440 28628 5480
rect 26092 5272 26132 5312
rect 27244 5272 27284 5312
rect 26572 5104 26612 5144
rect 26956 4768 26996 4808
rect 25996 4096 26036 4136
rect 26764 4684 26804 4724
rect 30604 5188 30644 5228
rect 27052 4600 27092 4640
rect 26956 4516 26996 4556
rect 26764 4432 26804 4472
rect 27052 4432 27092 4472
rect 27244 4684 27284 4724
rect 28588 4684 28628 4724
rect 29548 4684 29588 4724
rect 28012 4516 28052 4556
rect 25900 3424 25940 3464
rect 26572 3424 26612 3464
rect 26380 2500 26420 2540
rect 25996 2080 26036 2120
rect 26092 1660 26132 1700
rect 26764 4096 26804 4136
rect 27436 4096 27476 4136
rect 27628 3424 27668 3464
rect 26668 2668 26708 2708
rect 27820 2500 27860 2540
rect 27436 1828 27476 1868
rect 28492 4096 28532 4136
rect 29356 3844 29396 3884
rect 28204 2668 28244 2708
rect 28108 2584 28148 2624
rect 28204 2332 28244 2372
rect 28012 1492 28052 1532
rect 29644 4180 29684 4220
rect 30988 4684 31028 4724
rect 30508 4180 30548 4220
rect 30700 4180 30740 4220
rect 29644 3928 29684 3968
rect 30796 4096 30836 4136
rect 30604 4012 30644 4052
rect 30220 3844 30260 3884
rect 29932 3424 29972 3464
rect 34764 7204 34804 7244
rect 35212 7204 35252 7244
rect 33772 5524 33812 5564
rect 32716 5188 32756 5228
rect 31948 5104 31988 5144
rect 32140 5104 32180 5144
rect 32332 5104 32372 5144
rect 32428 4768 32468 4808
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 31948 4180 31988 4220
rect 32236 4096 32276 4136
rect 31756 3508 31796 3548
rect 29740 2584 29780 2624
rect 30508 2332 30548 2372
rect 29644 2164 29684 2204
rect 29356 1828 29396 1868
rect 28588 1576 28628 1616
rect 28492 1492 28532 1532
rect 30412 1828 30452 1868
rect 29548 1492 29588 1532
rect 31468 3424 31508 3464
rect 32236 3424 32276 3464
rect 31564 2668 31604 2708
rect 31468 2500 31508 2540
rect 30796 1912 30836 1952
rect 31756 2584 31796 2624
rect 32236 2584 32276 2624
rect 31948 2416 31988 2456
rect 32140 2416 32180 2456
rect 31660 2080 31700 2120
rect 34924 5440 34964 5480
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 34348 4180 34388 4220
rect 33484 4012 33524 4052
rect 33964 4012 34004 4052
rect 34252 4012 34292 4052
rect 34636 4180 34676 4220
rect 35404 4600 35444 4640
rect 35116 4096 35156 4136
rect 34732 4012 34772 4052
rect 34252 3844 34292 3884
rect 32524 3676 32564 3716
rect 32428 2836 32468 2876
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 34828 3928 34868 3968
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 34828 3592 34868 3632
rect 35308 4012 35348 4052
rect 35116 3676 35156 3716
rect 35116 3508 35156 3548
rect 35020 3424 35060 3464
rect 34924 3340 34964 3380
rect 35212 3424 35252 3464
rect 35308 3340 35348 3380
rect 34348 2668 34388 2708
rect 32524 2584 32564 2624
rect 34924 2752 34964 2792
rect 32716 2416 32756 2456
rect 32428 2164 32468 2204
rect 32332 1828 32372 1868
rect 32140 1492 32180 1532
rect 31564 1156 31604 1196
rect 31852 1072 31892 1112
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 34156 2164 34196 2204
rect 34732 1996 34772 2036
rect 33004 1912 33044 1952
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 32716 1408 32756 1448
rect 35500 3928 35540 3968
rect 35692 4096 35732 4136
rect 35692 3004 35732 3044
rect 35596 2752 35636 2792
rect 37132 6616 37172 6656
rect 36364 6448 36404 6488
rect 35980 5104 36020 5144
rect 35884 2164 35924 2204
rect 35404 1996 35444 2036
rect 35596 1912 35636 1952
rect 35692 1492 35732 1532
rect 34348 1324 34388 1364
rect 34828 1324 34868 1364
rect 34444 1240 34484 1280
rect 34156 1156 34196 1196
rect 34540 1072 34580 1112
rect 36940 5104 36980 5144
rect 37228 5356 37268 5396
rect 36940 3424 36980 3464
rect 37036 3340 37076 3380
rect 36748 3256 36788 3296
rect 36460 2584 36500 2624
rect 35980 1492 36020 1532
rect 36652 2500 36692 2540
rect 36556 1744 36596 1784
rect 36460 1156 36500 1196
rect 37324 3508 37364 3548
rect 37516 5692 37556 5732
rect 38860 6532 38900 6572
rect 38668 5692 38708 5732
rect 37612 5356 37652 5396
rect 38572 5104 38612 5144
rect 38764 5104 38804 5144
rect 39244 5272 39284 5312
rect 38764 4768 38804 4808
rect 38668 4684 38708 4724
rect 38572 3928 38612 3968
rect 38476 3676 38516 3716
rect 38380 3340 38420 3380
rect 39148 4768 39188 4808
rect 39340 4768 39380 4808
rect 38956 4684 38996 4724
rect 38860 3340 38900 3380
rect 38284 3088 38324 3128
rect 39052 2836 39092 2876
rect 38956 2752 38996 2792
rect 37516 2668 37556 2708
rect 38668 2584 38708 2624
rect 39052 2500 39092 2540
rect 39148 2164 39188 2204
rect 37324 1996 37364 2036
rect 36748 1744 36788 1784
rect 36652 1156 36692 1196
rect 36556 1072 36596 1112
rect 36844 1492 36884 1532
rect 38188 1912 38228 1952
rect 37324 1744 37364 1784
rect 39148 1744 39188 1784
rect 38764 1072 38804 1112
rect 39340 2248 39380 2288
rect 40889 7288 40929 7328
rect 40108 3508 40148 3548
rect 40012 3340 40052 3380
rect 39916 3256 39956 3296
rect 40300 4768 40340 4808
rect 40780 6448 40820 6488
rect 41260 5356 41300 5396
rect 40684 4348 40724 4388
rect 41260 4348 41300 4388
rect 40972 4264 41012 4304
rect 40780 4096 40820 4136
rect 41260 4096 41300 4136
rect 40876 3676 40916 3716
rect 41068 3424 41108 3464
rect 41260 3424 41300 3464
rect 41068 3256 41108 3296
rect 40972 3172 41012 3212
rect 40204 2752 40244 2792
rect 40012 2584 40052 2624
rect 40300 2584 40340 2624
rect 40396 2500 40436 2540
rect 39916 1996 39956 2036
rect 40012 1828 40052 1868
rect 39724 1240 39764 1280
rect 39628 1156 39668 1196
rect 39244 1072 39284 1112
rect 40300 2164 40340 2204
rect 40204 1576 40244 1616
rect 40588 2836 40628 2876
rect 41068 2836 41108 2876
rect 40684 1996 40724 2036
rect 42892 6448 42932 6488
rect 42508 4264 42548 4304
rect 42796 4096 42836 4136
rect 45196 4936 45236 4976
rect 46828 4852 46868 4892
rect 43852 4684 43892 4724
rect 43852 4264 43892 4304
rect 42316 3676 42356 3716
rect 42220 3172 42260 3212
rect 43180 3844 43220 3884
rect 43084 3508 43124 3548
rect 43372 4096 43412 4136
rect 43276 3424 43316 3464
rect 43180 3172 43220 3212
rect 42124 2584 42164 2624
rect 42316 2500 42356 2540
rect 41164 1912 41204 1952
rect 42892 2164 42932 2204
rect 42412 1492 42452 1532
rect 40492 1072 40532 1112
rect 43948 3508 43988 3548
rect 44524 3928 44564 3968
rect 45196 3592 45236 3632
rect 45388 3508 45428 3548
rect 44332 3004 44372 3044
rect 45484 2752 45524 2792
rect 43756 1912 43796 1952
rect 43372 1576 43412 1616
rect 44428 1492 44468 1532
rect 42508 1156 42548 1196
rect 42604 1072 42644 1112
rect 44812 1240 44852 1280
rect 44716 1072 44756 1112
rect 46156 4096 46196 4136
rect 46252 4012 46292 4052
rect 46060 3508 46100 3548
rect 45868 2668 45908 2708
rect 47116 4936 47156 4976
rect 46348 2836 46388 2876
rect 46924 3424 46964 3464
rect 47212 4180 47252 4220
rect 46636 2752 46676 2792
rect 47020 2752 47060 2792
rect 54604 5692 54644 5732
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 47500 4180 47540 4220
rect 47404 4096 47444 4136
rect 47308 4012 47348 4052
rect 50188 4180 50228 4220
rect 50380 4180 50420 4220
rect 48076 3592 48116 3632
rect 47404 3256 47444 3296
rect 47116 2668 47156 2708
rect 47596 2836 47636 2876
rect 47788 2500 47828 2540
rect 48652 4096 48692 4136
rect 49036 4012 49076 4052
rect 49228 4012 49268 4052
rect 49036 3760 49076 3800
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 49420 3928 49460 3968
rect 49420 3760 49460 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 49228 2836 49268 2876
rect 48364 2752 48404 2792
rect 49036 2752 49076 2792
rect 47308 1744 47348 1784
rect 48172 1744 48212 1784
rect 49516 2668 49556 2708
rect 50188 3424 50228 3464
rect 51724 4096 51764 4136
rect 51820 4012 51860 4052
rect 51724 3676 51764 3716
rect 50380 2752 50420 2792
rect 50956 2752 50996 2792
rect 51724 2668 51764 2708
rect 51244 2584 51284 2624
rect 49132 2500 49172 2540
rect 49708 2500 49748 2540
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 51436 2500 51476 2540
rect 49900 1996 49940 2036
rect 51244 1996 51284 2036
rect 51052 1744 51092 1784
rect 45868 1492 45908 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 47500 1240 47540 1280
rect 44908 1072 44948 1112
rect 52108 4936 52148 4976
rect 53644 4936 53684 4976
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 54604 4852 54644 4892
rect 53644 4348 53684 4388
rect 53356 4096 53396 4136
rect 53548 4096 53588 4136
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 54700 4348 54740 4388
rect 53356 3844 53396 3884
rect 52012 3424 52052 3464
rect 53740 3928 53780 3968
rect 55468 4096 55508 4136
rect 56620 3928 56660 3968
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 52972 3424 53012 3464
rect 52300 2752 52340 2792
rect 52684 2752 52724 2792
rect 51820 2584 51860 2624
rect 52396 2668 52436 2708
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 75532 17956 75572 17996
rect 81004 33664 81044 33704
rect 81100 33580 81140 33620
rect 80812 33496 80852 33536
rect 80812 32824 80852 32864
rect 81484 33664 81524 33704
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 80428 31648 80468 31688
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 79948 30556 79988 30596
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 79564 30052 79604 30092
rect 79180 29800 79220 29840
rect 79468 29212 79508 29252
rect 79180 29128 79220 29168
rect 79372 29128 79412 29168
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 78604 28624 78644 28664
rect 77740 17116 77780 17156
rect 80140 29800 80180 29840
rect 81388 32824 81428 32864
rect 81196 31732 81236 31772
rect 80620 30640 80660 30680
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 80428 29212 80468 29252
rect 80044 29128 80084 29168
rect 80332 28792 80372 28832
rect 80524 28792 80564 28832
rect 79756 28540 79796 28580
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 80716 30556 80756 30596
rect 82060 34168 82100 34208
rect 83212 34168 83252 34208
rect 81580 32404 81620 32444
rect 81196 30640 81236 30680
rect 81292 29800 81332 29840
rect 81484 29800 81524 29840
rect 81004 29128 81044 29168
rect 81292 28540 81332 28580
rect 81388 27784 81428 27824
rect 80812 27700 80852 27740
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 79372 26104 79412 26144
rect 79948 26104 79988 26144
rect 80236 26104 80276 26144
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 80332 26020 80372 26060
rect 83404 34168 83444 34208
rect 83404 33748 83444 33788
rect 83308 33664 83348 33704
rect 83116 33580 83156 33620
rect 81964 31648 82004 31688
rect 81868 30640 81908 30680
rect 83404 31396 83444 31436
rect 83116 31228 83156 31268
rect 92177 36688 92217 36728
rect 97516 31869 97556 31909
rect 82444 30052 82484 30092
rect 82060 29800 82100 29840
rect 82924 29716 82964 29756
rect 83212 29212 83252 29252
rect 82924 28792 82964 28832
rect 81772 28624 81812 28664
rect 82636 28540 82676 28580
rect 81676 27700 81716 27740
rect 80428 25936 80468 25976
rect 81292 26104 81332 26144
rect 80908 25936 80948 25976
rect 81292 25936 81332 25976
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 80812 25264 80852 25304
rect 80908 24592 80948 24632
rect 81196 24592 81236 24632
rect 80428 24508 80468 24548
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 79468 21568 79508 21608
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 81676 26104 81716 26144
rect 81676 25936 81716 25976
rect 81580 20812 81620 20852
rect 80620 20728 80660 20768
rect 81964 25264 82004 25304
rect 83212 27700 83252 27740
rect 83212 25936 83252 25976
rect 83116 24592 83156 24632
rect 85420 24592 85460 24632
rect 82924 24508 82964 24548
rect 82636 24424 82676 24464
rect 81772 21568 81812 21608
rect 89297 24508 89337 24548
rect 91601 24424 91641 24464
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 83980 21568 84020 21608
rect 85132 21316 85172 21356
rect 97420 21316 97460 21356
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 82060 20812 82100 20852
rect 85132 20812 85172 20852
rect 81964 20728 82004 20768
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 82732 20056 82772 20096
rect 98380 20056 98420 20096
rect 80620 17116 80660 17156
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 80620 9220 80660 9260
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 77644 6952 77684 6992
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 80236 6448 80276 6488
rect 78892 6364 78932 6404
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 96844 19888 96884 19928
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 98860 17956 98900 17996
rect 98860 9379 98900 9419
rect 82732 5104 82772 5144
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 74668 4012 74708 4052
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 81964 3088 82004 3128
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 74092 1912 74132 1952
rect 81964 1912 82004 1952
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 90737 1439 90777 1479
rect 91121 1439 91161 1479
rect 91313 1439 91353 1479
rect 90537 1240 90577 1280
rect 51820 1156 51860 1196
rect 54412 1156 54452 1196
rect 90892 988 90932 1028
rect 35884 904 35924 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 20995 38368 21004 38408
rect 21044 38368 22252 38408
rect 22292 38368 22301 38408
rect 28867 38368 28876 38408
rect 28916 38368 29260 38408
rect 29300 38368 29309 38408
rect 26851 38200 26860 38240
rect 26900 38200 27340 38240
rect 27380 38200 27389 38240
rect 27436 38200 28492 38240
rect 28532 38200 29452 38240
rect 29492 38200 31468 38240
rect 31508 38200 31517 38240
rect 38755 38200 38764 38240
rect 38804 38200 39820 38240
rect 39860 38200 41452 38240
rect 41492 38200 43468 38240
rect 43508 38200 43517 38240
rect 27436 38156 27476 38200
rect 27427 38116 27436 38156
rect 27476 38116 27485 38156
rect 835 37948 844 37988
rect 884 37948 5452 37988
rect 5492 37948 5501 37988
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 0 37568 80 37588
rect 0 37528 652 37568
rect 692 37528 701 37568
rect 0 37508 80 37528
rect 25891 37444 25900 37484
rect 25940 37444 26860 37484
rect 26900 37444 28876 37484
rect 28916 37444 28925 37484
rect 739 37360 748 37400
rect 788 37360 7220 37400
rect 21379 37360 21388 37400
rect 21428 37360 23788 37400
rect 23828 37360 23980 37400
rect 24020 37360 24029 37400
rect 27043 37360 27052 37400
rect 27092 37360 29452 37400
rect 29492 37360 32332 37400
rect 32372 37360 32381 37400
rect 33667 37360 33676 37400
rect 33716 37360 36652 37400
rect 36692 37360 39052 37400
rect 39092 37360 70636 37400
rect 70676 37360 70685 37400
rect 7180 37316 7220 37360
rect 7180 37276 19372 37316
rect 19412 37276 19421 37316
rect 20131 37276 20140 37316
rect 20180 37276 21292 37316
rect 21332 37276 21341 37316
rect 21763 37276 21772 37316
rect 21812 37276 21821 37316
rect 26371 37276 26380 37316
rect 26420 37276 26668 37316
rect 26708 37276 28780 37316
rect 28820 37276 28829 37316
rect 37795 37276 37804 37316
rect 37844 37276 39148 37316
rect 39188 37276 39197 37316
rect 21772 37232 21812 37276
rect 20611 37192 20620 37232
rect 20660 37192 33140 37232
rect 38467 37192 38476 37232
rect 38516 37192 40588 37232
rect 40628 37192 41068 37232
rect 41108 37192 41117 37232
rect 41347 37192 41356 37232
rect 41396 37192 41644 37232
rect 41684 37192 42220 37232
rect 42260 37192 44524 37232
rect 44564 37192 44573 37232
rect 33100 37148 33140 37192
rect 20899 37108 20908 37148
rect 20948 37108 21484 37148
rect 21524 37108 21772 37148
rect 21812 37108 26956 37148
rect 26996 37108 27005 37148
rect 33100 37108 42796 37148
rect 42836 37108 42845 37148
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 21571 37024 21580 37064
rect 21620 37024 22540 37064
rect 22580 37024 23500 37064
rect 23540 37024 24364 37064
rect 24404 37024 24413 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 23299 36940 23308 36980
rect 23348 36940 25228 36980
rect 25268 36940 26476 36980
rect 26516 36940 27148 36980
rect 27188 36940 27197 36980
rect 22915 36856 22924 36896
rect 22964 36856 24460 36896
rect 24500 36856 24844 36896
rect 24884 36856 24893 36896
rect 25315 36856 25324 36896
rect 25364 36856 26668 36896
rect 26708 36856 26717 36896
rect 28771 36856 28780 36896
rect 28820 36856 29452 36896
rect 29492 36856 30316 36896
rect 30356 36856 30365 36896
rect 38179 36856 38188 36896
rect 38228 36856 38860 36896
rect 38900 36856 41452 36896
rect 41492 36856 42508 36896
rect 42548 36856 42557 36896
rect 87820 36856 93329 36896
rect 93369 36856 93378 36896
rect 25324 36812 25364 36856
rect 19363 36772 19372 36812
rect 19412 36772 20428 36812
rect 20468 36772 20477 36812
rect 22348 36772 23308 36812
rect 23348 36772 23357 36812
rect 24643 36772 24652 36812
rect 24692 36772 25364 36812
rect 26755 36772 26764 36812
rect 26804 36772 27916 36812
rect 27956 36772 27965 36812
rect 41059 36772 41068 36812
rect 41108 36772 41740 36812
rect 41780 36772 41789 36812
rect 0 36728 80 36748
rect 22348 36728 22388 36772
rect 87820 36728 87860 36856
rect 0 36688 7084 36728
rect 7124 36688 7133 36728
rect 17827 36688 17836 36728
rect 17876 36688 18892 36728
rect 18932 36688 18941 36728
rect 19075 36688 19084 36728
rect 19124 36688 21388 36728
rect 21428 36688 21437 36728
rect 21571 36688 21580 36728
rect 21620 36688 21772 36728
rect 21812 36688 21821 36728
rect 22339 36688 22348 36728
rect 22388 36688 22397 36728
rect 23011 36688 23020 36728
rect 23060 36688 23884 36728
rect 23924 36688 23933 36728
rect 25219 36688 25228 36728
rect 25268 36688 25844 36728
rect 26083 36688 26092 36728
rect 26132 36688 26860 36728
rect 26900 36688 27340 36728
rect 27380 36688 27389 36728
rect 27523 36688 27532 36728
rect 27572 36688 30316 36728
rect 30356 36688 31180 36728
rect 31220 36688 33676 36728
rect 33716 36688 33725 36728
rect 38563 36688 38572 36728
rect 38612 36688 39724 36728
rect 39764 36688 42316 36728
rect 42356 36688 74092 36728
rect 74132 36688 74141 36728
rect 83491 36688 83500 36728
rect 83540 36688 87860 36728
rect 89548 36772 91217 36812
rect 91257 36772 91266 36812
rect 0 36668 80 36688
rect 25804 36644 25844 36688
rect 27340 36644 27380 36688
rect 89548 36644 89588 36772
rect 19171 36604 19180 36644
rect 19220 36604 20236 36644
rect 20276 36604 20716 36644
rect 20756 36604 20765 36644
rect 23683 36604 23692 36644
rect 23732 36604 25516 36644
rect 25556 36604 25565 36644
rect 25804 36604 26572 36644
rect 26612 36604 26621 36644
rect 27340 36604 27628 36644
rect 27668 36604 28012 36644
rect 28052 36604 28061 36644
rect 83299 36604 83308 36644
rect 83348 36604 89588 36644
rect 90028 36688 92177 36728
rect 92217 36688 92226 36728
rect 23491 36520 23500 36560
rect 23540 36520 23980 36560
rect 24020 36520 24029 36560
rect 25891 36520 25900 36560
rect 25940 36520 27052 36560
rect 27092 36520 27724 36560
rect 27764 36520 28684 36560
rect 28724 36520 28733 36560
rect 71971 36476 72029 36477
rect 90028 36476 90068 36688
rect 19363 36436 19372 36476
rect 19412 36436 21004 36476
rect 21044 36436 21053 36476
rect 22435 36436 22444 36476
rect 22484 36436 23692 36476
rect 23732 36436 23741 36476
rect 71971 36436 71980 36476
rect 72020 36436 90068 36476
rect 71971 36435 72029 36436
rect 25507 36352 25516 36392
rect 25556 36352 26188 36392
rect 26228 36352 27052 36392
rect 27092 36352 27101 36392
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 21667 36268 21676 36308
rect 21716 36268 21964 36308
rect 22004 36268 23212 36308
rect 23252 36268 23884 36308
rect 23924 36268 25228 36308
rect 25268 36268 25277 36308
rect 25987 36268 25996 36308
rect 26036 36268 26380 36308
rect 26420 36268 26429 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 5443 36184 5452 36224
rect 5492 36184 45292 36224
rect 45332 36184 45341 36224
rect 38467 36100 38476 36140
rect 38516 36100 39148 36140
rect 39188 36100 39197 36140
rect 70627 36056 70685 36057
rect 71971 36056 72029 36057
rect 7075 36016 7084 36056
rect 7124 36016 34444 36056
rect 34484 36016 34493 36056
rect 47971 36016 47980 36056
rect 48020 36016 70636 36056
rect 70676 36016 71980 36056
rect 72020 36016 72029 36056
rect 70627 36015 70685 36016
rect 71971 36015 72029 36016
rect 35107 35932 35116 35972
rect 35156 35932 38380 35972
rect 38420 35932 38668 35972
rect 38708 35932 38717 35972
rect 40291 35932 40300 35972
rect 40340 35932 65260 35972
rect 65300 35932 65309 35972
rect 0 35888 80 35908
rect 35116 35888 35156 35932
rect 0 35848 2572 35888
rect 2612 35848 2621 35888
rect 6403 35848 6412 35888
rect 6452 35848 13708 35888
rect 13748 35848 13757 35888
rect 15523 35848 15532 35888
rect 15572 35848 16492 35888
rect 16532 35848 17452 35888
rect 17492 35848 17501 35888
rect 18307 35848 18316 35888
rect 18356 35848 19756 35888
rect 19796 35848 21196 35888
rect 21236 35848 21245 35888
rect 22819 35848 22828 35888
rect 22868 35848 23116 35888
rect 23156 35848 25900 35888
rect 25940 35848 25949 35888
rect 31267 35848 31276 35888
rect 31316 35848 31564 35888
rect 31604 35848 35156 35888
rect 38947 35848 38956 35888
rect 38996 35848 39916 35888
rect 39956 35848 40108 35888
rect 40148 35848 40157 35888
rect 40387 35848 40396 35888
rect 40436 35848 40876 35888
rect 40916 35848 41836 35888
rect 41876 35848 41885 35888
rect 42115 35848 42124 35888
rect 42164 35848 43852 35888
rect 43892 35848 43901 35888
rect 65923 35848 65932 35888
rect 65972 35848 70348 35888
rect 70388 35848 72268 35888
rect 72308 35848 73900 35888
rect 73940 35848 73949 35888
rect 0 35828 80 35848
rect 13708 35720 13748 35848
rect 24259 35804 24317 35805
rect 40396 35804 40436 35848
rect 42124 35804 42164 35848
rect 14563 35764 14572 35804
rect 14612 35764 17356 35804
rect 17396 35764 17684 35804
rect 19939 35764 19948 35804
rect 19988 35764 20620 35804
rect 20660 35764 21292 35804
rect 21332 35764 21341 35804
rect 24174 35764 24268 35804
rect 24308 35764 24317 35804
rect 31459 35764 31468 35804
rect 31508 35764 31948 35804
rect 31988 35764 34828 35804
rect 34868 35764 35308 35804
rect 35348 35764 35357 35804
rect 35779 35764 35788 35804
rect 35828 35764 37900 35804
rect 37940 35764 38188 35804
rect 38228 35764 38237 35804
rect 38755 35764 38764 35804
rect 38804 35764 39532 35804
rect 39572 35764 40436 35804
rect 41635 35764 41644 35804
rect 41684 35764 42164 35804
rect 52675 35764 52684 35804
rect 52724 35764 53548 35804
rect 53588 35764 53597 35804
rect 17644 35720 17684 35764
rect 24259 35763 24317 35764
rect 69187 35720 69245 35721
rect 13708 35680 17588 35720
rect 17635 35680 17644 35720
rect 17684 35680 17693 35720
rect 20803 35680 20812 35720
rect 20852 35680 21004 35720
rect 21044 35680 27532 35720
rect 27572 35680 27581 35720
rect 30115 35680 30124 35720
rect 30164 35680 35500 35720
rect 35540 35680 37460 35720
rect 37795 35680 37804 35720
rect 37844 35680 47020 35720
rect 47060 35680 47069 35720
rect 50179 35680 50188 35720
rect 50228 35680 52300 35720
rect 52340 35680 53260 35720
rect 53300 35680 69196 35720
rect 69236 35680 69245 35720
rect 17548 35636 17588 35680
rect 20812 35636 20852 35680
rect 37420 35636 37460 35680
rect 37804 35636 37844 35680
rect 69187 35679 69245 35680
rect 14659 35596 14668 35636
rect 14708 35596 15628 35636
rect 15668 35596 16876 35636
rect 16916 35596 17300 35636
rect 17548 35596 20852 35636
rect 24163 35596 24172 35636
rect 24212 35596 35020 35636
rect 35060 35596 35788 35636
rect 35828 35596 35837 35636
rect 37420 35596 37844 35636
rect 38467 35596 38476 35636
rect 38516 35596 43564 35636
rect 43604 35596 43613 35636
rect 43939 35596 43948 35636
rect 43988 35596 79564 35636
rect 79604 35596 79613 35636
rect 17260 35552 17300 35596
rect 69091 35552 69149 35553
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 17260 35512 18124 35552
rect 18164 35512 19372 35552
rect 19412 35512 19421 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 23587 35512 23596 35552
rect 23636 35512 30220 35552
rect 30260 35512 32524 35552
rect 32564 35512 32716 35552
rect 32756 35512 32765 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 43843 35512 43852 35552
rect 43892 35512 46828 35552
rect 46868 35512 46877 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 65251 35512 65260 35552
rect 65300 35512 69100 35552
rect 69140 35512 69149 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 69091 35511 69149 35512
rect 28387 35428 28396 35468
rect 28436 35428 29260 35468
rect 29300 35428 29309 35468
rect 41539 35428 41548 35468
rect 41588 35428 47596 35468
rect 47636 35428 48268 35468
rect 48308 35428 48317 35468
rect 41155 35384 41213 35385
rect 18691 35344 18700 35384
rect 18740 35344 21580 35384
rect 21620 35344 21629 35384
rect 25603 35344 25612 35384
rect 25652 35344 27244 35384
rect 27284 35344 27293 35384
rect 27715 35344 27724 35384
rect 27764 35344 28012 35384
rect 28052 35344 28972 35384
rect 29012 35344 29021 35384
rect 29347 35344 29356 35384
rect 29396 35344 31852 35384
rect 31892 35344 32236 35384
rect 32276 35344 32285 35384
rect 41070 35344 41164 35384
rect 41204 35344 41213 35384
rect 44419 35344 44428 35384
rect 44468 35344 45484 35384
rect 45524 35344 81772 35384
rect 81812 35344 81821 35384
rect 41155 35343 41213 35344
rect 33859 35260 33868 35300
rect 33908 35260 38476 35300
rect 38516 35260 38525 35300
rect 42019 35260 42028 35300
rect 42068 35260 43372 35300
rect 43412 35260 45292 35300
rect 45332 35260 45676 35300
rect 45716 35260 49228 35300
rect 49268 35260 49277 35300
rect 14179 35176 14188 35216
rect 14228 35176 15628 35216
rect 15668 35176 18316 35216
rect 18356 35176 18365 35216
rect 19843 35176 19852 35216
rect 19892 35176 24460 35216
rect 24500 35176 25708 35216
rect 25748 35176 33484 35216
rect 33524 35176 33533 35216
rect 34627 35176 34636 35216
rect 34676 35176 35500 35216
rect 35540 35176 35549 35216
rect 35875 35176 35884 35216
rect 35924 35176 72652 35216
rect 72692 35176 72701 35216
rect 12259 35132 12317 35133
rect 12174 35092 12268 35132
rect 12308 35092 12317 35132
rect 12451 35092 12460 35132
rect 12500 35092 14668 35132
rect 14708 35092 14717 35132
rect 12259 35091 12317 35092
rect 0 34988 80 35068
rect 33484 35048 33524 35176
rect 39052 35092 46924 35132
rect 46964 35092 46973 35132
rect 47875 35092 47884 35132
rect 47924 35092 48364 35132
rect 48404 35092 50956 35132
rect 50996 35092 53548 35132
rect 53588 35092 53597 35132
rect 39052 35048 39092 35092
rect 47884 35048 47924 35092
rect 18595 35008 18604 35048
rect 18644 35008 20140 35048
rect 20180 35008 20189 35048
rect 21283 35008 21292 35048
rect 21332 35008 33140 35048
rect 33484 35008 37612 35048
rect 37652 35008 38092 35048
rect 38132 35008 38141 35048
rect 39043 35008 39052 35048
rect 39092 35008 39101 35048
rect 42787 35008 42796 35048
rect 42836 35008 43756 35048
rect 43796 35008 43805 35048
rect 44803 35008 44812 35048
rect 44852 35008 47924 35048
rect 13795 34924 13804 34964
rect 13844 34924 14476 34964
rect 14516 34924 16684 34964
rect 16724 34924 23980 34964
rect 24020 34924 24029 34964
rect 33100 34880 33140 35008
rect 41347 34924 41356 34964
rect 41396 34924 41405 34964
rect 46531 34924 46540 34964
rect 46580 34924 46732 34964
rect 46772 34924 47788 34964
rect 47828 34924 50188 34964
rect 50228 34924 50237 34964
rect 50371 34924 50380 34964
rect 50420 34924 50429 34964
rect 53731 34924 53740 34964
rect 53780 34924 55564 34964
rect 55604 34924 55613 34964
rect 41356 34880 41396 34924
rect 50380 34880 50420 34924
rect 19555 34840 19564 34880
rect 19604 34840 21292 34880
rect 21332 34840 21341 34880
rect 33100 34840 41396 34880
rect 46915 34840 46924 34880
rect 46964 34840 48076 34880
rect 48116 34840 50420 34880
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 33964 34756 41356 34796
rect 41396 34756 41405 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 49036 34756 49228 34796
rect 49268 34756 51916 34796
rect 51956 34756 51965 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 26563 34672 26572 34712
rect 26612 34672 33868 34712
rect 33908 34672 33917 34712
rect 33964 34628 34004 34756
rect 37516 34672 39436 34712
rect 39476 34672 39485 34712
rect 42883 34672 42892 34712
rect 42932 34672 43468 34712
rect 43508 34672 43517 34712
rect 37516 34628 37556 34672
rect 49036 34628 49076 34756
rect 51811 34672 51820 34712
rect 51860 34672 53644 34712
rect 53684 34672 54412 34712
rect 54452 34672 55372 34712
rect 55412 34672 55421 34712
rect 20131 34588 20140 34628
rect 20180 34588 23404 34628
rect 23444 34588 23453 34628
rect 28963 34588 28972 34628
rect 29012 34588 31180 34628
rect 31220 34588 34004 34628
rect 37315 34588 37324 34628
rect 37364 34588 37556 34628
rect 47203 34588 47212 34628
rect 47252 34588 47980 34628
rect 48020 34588 48029 34628
rect 48643 34588 48652 34628
rect 48692 34588 49076 34628
rect 7363 34504 7372 34544
rect 7412 34504 17068 34544
rect 17108 34504 19852 34544
rect 19892 34504 19901 34544
rect 20803 34504 20812 34544
rect 20852 34504 21388 34544
rect 21428 34504 22252 34544
rect 22292 34504 22301 34544
rect 25891 34504 25900 34544
rect 25940 34504 26860 34544
rect 26900 34504 29260 34544
rect 29300 34504 31084 34544
rect 31124 34504 33388 34544
rect 33428 34504 35884 34544
rect 35924 34504 35933 34544
rect 38083 34504 38092 34544
rect 38132 34504 43372 34544
rect 43412 34504 43421 34544
rect 46435 34504 46444 34544
rect 46484 34504 48844 34544
rect 48884 34504 48893 34544
rect 49123 34504 49132 34544
rect 49172 34504 49804 34544
rect 49844 34504 50380 34544
rect 50420 34504 50429 34544
rect 51523 34504 51532 34544
rect 51572 34504 52780 34544
rect 52820 34504 61516 34544
rect 61556 34504 65932 34544
rect 65972 34504 65981 34544
rect 25027 34420 25036 34460
rect 25076 34420 25996 34460
rect 26036 34420 28396 34460
rect 28436 34420 28445 34460
rect 29347 34420 29356 34460
rect 29396 34420 29836 34460
rect 29876 34420 30412 34460
rect 30452 34420 30461 34460
rect 4963 34336 4972 34376
rect 5012 34336 7372 34376
rect 7412 34336 7421 34376
rect 16003 34336 16012 34376
rect 16052 34336 18892 34376
rect 18932 34336 19372 34376
rect 19412 34336 20044 34376
rect 20084 34336 20093 34376
rect 24067 34336 24076 34376
rect 24116 34336 27052 34376
rect 27092 34336 28780 34376
rect 28820 34336 29548 34376
rect 29588 34336 29597 34376
rect 32899 34336 32908 34376
rect 32948 34336 64684 34376
rect 64724 34336 64733 34376
rect 11299 34252 11308 34292
rect 11348 34252 13708 34292
rect 13748 34252 14188 34292
rect 14228 34252 17300 34292
rect 0 34148 80 34228
rect 17260 34208 17300 34252
rect 4771 34168 4780 34208
rect 4820 34168 13036 34208
rect 13076 34168 15244 34208
rect 15284 34168 15532 34208
rect 15572 34168 15581 34208
rect 17260 34168 18796 34208
rect 18836 34168 18845 34208
rect 31555 34168 31564 34208
rect 31604 34168 33004 34208
rect 33044 34168 35212 34208
rect 35252 34168 37036 34208
rect 37076 34168 37085 34208
rect 42307 34168 42316 34208
rect 42356 34168 43564 34208
rect 43604 34168 43613 34208
rect 43747 34168 43756 34208
rect 43796 34168 51532 34208
rect 51572 34168 51581 34208
rect 52483 34168 52492 34208
rect 52532 34168 62612 34208
rect 66883 34168 66892 34208
rect 66932 34168 82060 34208
rect 82100 34168 82109 34208
rect 83203 34168 83212 34208
rect 83252 34168 83404 34208
rect 83444 34168 83453 34208
rect 8419 34124 8477 34125
rect 42316 34124 42356 34168
rect 61027 34124 61085 34125
rect 8419 34084 8428 34124
rect 8468 34084 31660 34124
rect 31700 34084 34444 34124
rect 34484 34084 34493 34124
rect 41251 34084 41260 34124
rect 41300 34084 41644 34124
rect 41684 34084 42356 34124
rect 53539 34084 53548 34124
rect 53588 34084 54508 34124
rect 54548 34084 61036 34124
rect 61076 34084 61085 34124
rect 62572 34124 62612 34168
rect 69475 34124 69533 34125
rect 62572 34084 69484 34124
rect 69524 34084 69533 34124
rect 8419 34083 8477 34084
rect 61027 34083 61085 34084
rect 69475 34083 69533 34084
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 5251 34000 5260 34040
rect 5300 34000 10924 34040
rect 10964 34000 13420 34040
rect 13460 34000 13469 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 42691 34000 42700 34040
rect 42740 34000 46444 34040
rect 46484 34000 46493 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 50371 34000 50380 34040
rect 50420 34000 52972 34040
rect 53012 34000 53021 34040
rect 53827 34000 53836 34040
rect 53876 34000 56524 34040
rect 56564 34000 56573 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 8227 33916 8236 33956
rect 8276 33916 24844 33956
rect 24884 33916 24893 33956
rect 32899 33916 32908 33956
rect 32948 33916 35116 33956
rect 35156 33916 39148 33956
rect 39188 33916 39724 33956
rect 39764 33916 39773 33956
rect 68803 33872 68861 33873
rect 5539 33832 5548 33872
rect 5588 33832 37612 33872
rect 37652 33832 37661 33872
rect 45187 33832 45196 33872
rect 45236 33832 68812 33872
rect 68852 33832 68861 33872
rect 68803 33831 68861 33832
rect 1123 33748 1132 33788
rect 1172 33748 24172 33788
rect 24212 33748 24221 33788
rect 79555 33748 79564 33788
rect 79604 33748 80140 33788
rect 80180 33748 83404 33788
rect 83444 33748 83453 33788
rect 69379 33704 69437 33705
rect 42211 33664 42220 33704
rect 42260 33664 43180 33704
rect 43220 33664 69388 33704
rect 69428 33664 69437 33704
rect 79747 33664 79756 33704
rect 79796 33664 80716 33704
rect 80756 33664 80765 33704
rect 80995 33664 81004 33704
rect 81044 33664 81484 33704
rect 81524 33664 83308 33704
rect 83348 33664 83357 33704
rect 69379 33663 69437 33664
rect 46819 33580 46828 33620
rect 46868 33580 47500 33620
rect 47540 33580 47549 33620
rect 48835 33580 48844 33620
rect 48884 33580 52492 33620
rect 52532 33580 52541 33620
rect 80035 33580 80044 33620
rect 80084 33580 81100 33620
rect 81140 33580 83116 33620
rect 83156 33580 83165 33620
rect 69283 33536 69341 33537
rect 47107 33496 47116 33536
rect 47156 33496 48940 33536
rect 48980 33496 49132 33536
rect 49172 33496 49181 33536
rect 57580 33496 69292 33536
rect 69332 33496 69341 33536
rect 80419 33496 80428 33536
rect 80468 33496 80812 33536
rect 80852 33496 80861 33536
rect 57580 33452 57620 33496
rect 69283 33495 69341 33496
rect 41827 33412 41836 33452
rect 41876 33412 42508 33452
rect 42548 33412 57620 33452
rect 0 33308 80 33388
rect 85036 33370 85440 33410
rect 72643 33368 72701 33369
rect 85036 33368 85076 33370
rect 47491 33328 47500 33368
rect 47540 33328 49132 33368
rect 49172 33328 53836 33368
rect 53876 33328 53885 33368
rect 72643 33328 72652 33368
rect 72692 33328 85076 33368
rect 72643 33327 72701 33328
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 99811 33200 99869 33201
rect 99920 33200 100000 33220
rect 99811 33160 99820 33200
rect 99860 33160 100000 33200
rect 99811 33159 99869 33160
rect 99920 33140 100000 33160
rect 12259 33116 12317 33117
rect 5635 33076 5644 33116
rect 5684 33076 12268 33116
rect 12308 33076 12317 33116
rect 49507 33076 49516 33116
rect 49556 33076 63340 33116
rect 63380 33076 63389 33116
rect 12259 33075 12317 33076
rect 68995 32864 69053 32865
rect 41731 32824 41740 32864
rect 41780 32824 69004 32864
rect 69044 32824 69053 32864
rect 80803 32824 80812 32864
rect 80852 32824 81388 32864
rect 81428 32824 81437 32864
rect 68995 32823 69053 32824
rect 48259 32740 48268 32780
rect 48308 32740 77356 32780
rect 77396 32740 80428 32780
rect 80468 32740 80477 32780
rect 63331 32572 63340 32612
rect 63380 32572 76108 32612
rect 76148 32572 76157 32612
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 8323 32488 8332 32528
rect 8372 32488 26092 32528
rect 26132 32488 26141 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 8515 32444 8573 32445
rect 60739 32444 60797 32445
rect 8515 32404 8524 32444
rect 8564 32404 33772 32444
rect 33812 32404 33821 32444
rect 55363 32404 55372 32444
rect 55412 32404 60748 32444
rect 60788 32404 60797 32444
rect 62467 32404 62476 32444
rect 62516 32404 81580 32444
rect 81620 32404 81629 32444
rect 8515 32403 8573 32404
rect 60739 32403 60797 32404
rect 4387 32068 4396 32108
rect 4436 32068 5644 32108
rect 5684 32068 5693 32108
rect 3811 31900 3820 31940
rect 3860 31900 4588 31940
rect 4628 31900 20236 31940
rect 20276 31900 20285 31940
rect 97360 31869 97516 31909
rect 97556 31869 97565 31909
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 3628 31732 4396 31772
rect 4436 31732 4445 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 81187 31732 81196 31772
rect 81236 31732 81245 31772
rect 0 31628 80 31708
rect 3628 31688 3668 31732
rect 81196 31688 81236 31732
rect 2659 31648 2668 31688
rect 2708 31648 3668 31688
rect 5731 31648 5740 31688
rect 5780 31648 17356 31688
rect 17396 31648 18041 31688
rect 18081 31648 18090 31688
rect 18220 31648 18268 31688
rect 18308 31648 18700 31688
rect 18740 31648 18749 31688
rect 80419 31648 80428 31688
rect 80468 31648 81964 31688
rect 82004 31648 82013 31688
rect 18220 31604 18260 31648
rect 7843 31564 7852 31604
rect 7892 31564 18260 31604
rect 5923 31480 5932 31520
rect 5972 31480 11212 31520
rect 11252 31480 15161 31520
rect 15201 31480 15210 31520
rect 15907 31480 15916 31520
rect 15956 31480 15965 31520
rect 15916 31380 15956 31480
rect 83395 31396 83404 31436
rect 83444 31396 85421 31436
rect 15916 31352 16313 31380
rect 4867 31312 4876 31352
rect 4916 31312 5836 31352
rect 5876 31340 16313 31352
rect 16353 31340 16362 31380
rect 5876 31312 15956 31340
rect 83107 31228 83116 31268
rect 83156 31228 85421 31268
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 0 30788 80 30868
rect 4483 30724 4492 30764
rect 4532 30724 5260 30764
rect 5300 30724 5309 30764
rect 4771 30640 4780 30680
rect 4820 30640 5356 30680
rect 5396 30640 5405 30680
rect 80611 30640 80620 30680
rect 80660 30640 81196 30680
rect 81236 30640 81868 30680
rect 81908 30640 81917 30680
rect 4867 30556 4876 30596
rect 4916 30556 5740 30596
rect 5780 30556 5789 30596
rect 79939 30556 79948 30596
rect 79988 30556 80716 30596
rect 80756 30556 80765 30596
rect 3427 30472 3436 30512
rect 3476 30472 5164 30512
rect 5204 30472 5213 30512
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 83491 30092 83549 30093
rect 79555 30052 79564 30092
rect 79604 30052 82444 30092
rect 82484 30052 83500 30092
rect 83540 30052 83549 30092
rect 83491 30051 83549 30052
rect 97323 30091 97365 30100
rect 97323 30051 97324 30091
rect 97364 30051 97365 30091
rect 97323 30042 97365 30051
rect 0 29948 80 30028
rect 79171 29800 79180 29840
rect 79220 29800 80140 29840
rect 80180 29800 80189 29840
rect 81283 29800 81292 29840
rect 81332 29800 81484 29840
rect 81524 29800 82060 29840
rect 82100 29800 82109 29840
rect 82915 29716 82924 29756
rect 82964 29716 85421 29756
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 79459 29212 79468 29252
rect 79508 29212 80428 29252
rect 80468 29212 83212 29252
rect 83252 29212 83261 29252
rect 0 29108 80 29188
rect 79171 29128 79180 29168
rect 79220 29128 79372 29168
rect 79412 29128 80044 29168
rect 80084 29128 81004 29168
rect 81044 29128 81053 29168
rect 97323 29061 97365 29070
rect 97323 29021 97324 29061
rect 97364 29021 97365 29061
rect 97323 29012 97365 29021
rect 80323 28792 80332 28832
rect 80372 28792 80524 28832
rect 80564 28792 82924 28832
rect 82964 28792 82973 28832
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 78595 28624 78604 28664
rect 78644 28624 81772 28664
rect 81812 28624 81821 28664
rect 79747 28540 79756 28580
rect 79796 28540 81292 28580
rect 81332 28540 82636 28580
rect 82676 28540 82685 28580
rect 0 28268 80 28348
rect 4771 28288 4780 28328
rect 4820 28288 5068 28328
rect 5108 28288 5117 28328
rect 4963 28036 4972 28076
rect 5012 28036 5548 28076
rect 5588 28036 5597 28076
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 81379 27784 81388 27824
rect 81428 27784 83252 27824
rect 83212 27740 83252 27784
rect 80803 27700 80812 27740
rect 80852 27700 81676 27740
rect 81716 27700 81725 27740
rect 83203 27700 83212 27740
rect 83252 27700 85421 27740
rect 3427 27616 3436 27656
rect 3476 27616 5164 27656
rect 5204 27616 5213 27656
rect 0 27428 80 27508
rect 5251 27364 5260 27404
rect 5300 27364 5836 27404
rect 5876 27364 5885 27404
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 4867 26692 4876 26732
rect 4916 26692 5164 26732
rect 5204 26692 5213 26732
rect 0 26588 80 26668
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 79363 26104 79372 26144
rect 79412 26104 79948 26144
rect 79988 26104 80236 26144
rect 80276 26104 81292 26144
rect 81332 26104 81341 26144
rect 81667 26104 81676 26144
rect 81716 26104 83252 26144
rect 81676 26060 81716 26104
rect 80323 26020 80332 26060
rect 80372 26020 81716 26060
rect 83212 25976 83252 26104
rect 84931 25976 84989 25977
rect 6019 25936 6028 25976
rect 6068 25936 8021 25976
rect 80419 25936 80428 25976
rect 80468 25936 80908 25976
rect 80948 25936 80957 25976
rect 81283 25936 81292 25976
rect 81332 25936 81676 25976
rect 81716 25936 81725 25976
rect 83203 25936 83212 25976
rect 83252 25936 84940 25976
rect 84980 25936 84989 25976
rect 84931 25935 84989 25936
rect 0 25748 80 25828
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 80803 25264 80812 25304
rect 80852 25264 81964 25304
rect 82004 25264 82013 25304
rect 3427 25180 3436 25220
rect 3476 25180 5068 25220
rect 5108 25180 5117 25220
rect 835 25096 844 25136
rect 884 25096 1324 25136
rect 1364 25096 1373 25136
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 0 24908 80 24928
rect 4771 24676 4780 24716
rect 4820 24676 5836 24716
rect 5876 24676 5885 24716
rect 80899 24592 80908 24632
rect 80948 24592 81196 24632
rect 81236 24592 83116 24632
rect 83156 24592 85420 24632
rect 85460 24592 85469 24632
rect 80419 24508 80428 24548
rect 80468 24508 82924 24548
rect 82964 24508 89297 24548
rect 89337 24508 89346 24548
rect 82627 24424 82636 24464
rect 82676 24424 91601 24464
rect 91641 24424 91650 24464
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 0 24068 80 24088
rect 835 24004 844 24044
rect 884 24004 1132 24044
rect 1172 24004 1181 24044
rect 82915 23792 82973 23793
rect 99907 23792 99965 23793
rect 82915 23752 82924 23792
rect 82964 23752 99916 23792
rect 99956 23752 99965 23792
rect 82915 23751 82973 23752
rect 99907 23751 99965 23752
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 0 23288 80 23308
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 0 23228 80 23248
rect 3427 23080 3436 23120
rect 3476 23080 4396 23120
rect 4436 23080 4445 23120
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 0 22448 80 22468
rect 0 22408 652 22448
rect 692 22408 701 22448
rect 0 22388 80 22408
rect 3715 22324 3724 22364
rect 3764 22324 3916 22364
rect 3956 22324 4204 22364
rect 4244 22324 4253 22364
rect 4099 22240 4108 22280
rect 4148 22240 4588 22280
rect 4628 22240 5932 22280
rect 5972 22240 5981 22280
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 5827 21904 5836 21944
rect 5876 21904 8021 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 0 21608 80 21628
rect 0 21568 844 21608
rect 884 21568 893 21608
rect 79459 21568 79468 21608
rect 79508 21568 81772 21608
rect 81812 21568 83980 21608
rect 84020 21568 84029 21608
rect 0 21548 80 21568
rect 5347 21484 5356 21524
rect 5396 21484 5836 21524
rect 5876 21484 5885 21524
rect 85123 21316 85132 21356
rect 85172 21316 97420 21356
rect 97460 21316 97469 21356
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 5923 20896 5932 20936
rect 5972 20896 8021 20936
rect 2083 20812 2092 20852
rect 2132 20812 3916 20852
rect 3956 20812 3965 20852
rect 4771 20812 4780 20852
rect 4820 20812 7756 20852
rect 7796 20812 7805 20852
rect 81571 20812 81580 20852
rect 81620 20812 82060 20852
rect 82100 20812 85132 20852
rect 85172 20812 85181 20852
rect 0 20768 80 20788
rect 0 20728 844 20768
rect 884 20728 893 20768
rect 1603 20728 1612 20768
rect 1652 20728 3340 20768
rect 3380 20728 3820 20768
rect 3860 20728 3869 20768
rect 80611 20728 80620 20768
rect 80660 20728 81964 20768
rect 82004 20728 82013 20768
rect 0 20708 80 20728
rect 2467 20644 2476 20684
rect 2516 20644 4012 20684
rect 4052 20644 5356 20684
rect 5396 20644 5405 20684
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 4291 20140 4300 20180
rect 4340 20140 5260 20180
rect 5300 20140 5309 20180
rect 1219 20056 1228 20096
rect 1268 20056 2284 20096
rect 2324 20056 2333 20096
rect 2467 20056 2476 20096
rect 2516 20056 4108 20096
rect 4148 20056 4157 20096
rect 82723 20056 82732 20096
rect 82772 20056 98380 20096
rect 98420 20056 98429 20096
rect 0 19928 80 19948
rect 99920 19928 100000 19948
rect 0 19888 844 19928
rect 884 19888 893 19928
rect 3523 19888 3532 19928
rect 3572 19888 4588 19928
rect 4628 19888 4637 19928
rect 96835 19888 96844 19928
rect 96884 19888 100000 19928
rect 0 19868 80 19888
rect 99920 19868 100000 19888
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 1987 19552 1996 19592
rect 2036 19552 3628 19592
rect 3668 19552 4204 19592
rect 4244 19552 7700 19592
rect 3523 19468 3532 19508
rect 3572 19468 5068 19508
rect 5108 19468 5117 19508
rect 3427 19384 3436 19424
rect 3476 19384 4684 19424
rect 4724 19384 4733 19424
rect 2467 19300 2476 19340
rect 2516 19300 2668 19340
rect 2708 19300 2717 19340
rect 4867 19300 4876 19340
rect 4916 19300 6412 19340
rect 6452 19300 6461 19340
rect 2371 19216 2380 19256
rect 2420 19216 4396 19256
rect 4436 19216 6028 19256
rect 6068 19216 6077 19256
rect 7660 19130 7700 19552
rect 0 19088 80 19108
rect 7660 19090 8040 19130
rect 0 19048 844 19088
rect 884 19048 893 19088
rect 0 19028 80 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 5347 18880 5356 18920
rect 5396 18880 8021 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 1603 18628 1612 18668
rect 1652 18628 3724 18668
rect 3764 18628 4300 18668
rect 4340 18628 4349 18668
rect 2275 18460 2284 18500
rect 2324 18460 2668 18500
rect 2708 18460 2717 18500
rect 2083 18376 2092 18416
rect 2132 18376 3820 18416
rect 3860 18376 3869 18416
rect 0 18248 80 18268
rect 0 18208 844 18248
rect 884 18208 893 18248
rect 2275 18208 2284 18248
rect 2324 18208 2764 18248
rect 2804 18208 2813 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 835 18040 844 18080
rect 884 18040 1612 18080
rect 1652 18040 1661 18080
rect 4003 17956 4012 17996
rect 4052 17956 4492 17996
rect 4532 17956 4541 17996
rect 75523 17956 75532 17996
rect 75572 17956 98860 17996
rect 98900 17956 98909 17996
rect 1219 17872 1228 17912
rect 1268 17872 1804 17912
rect 1844 17872 4108 17912
rect 4148 17872 8021 17912
rect 0 17408 80 17428
rect 0 17368 844 17408
rect 884 17368 893 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 0 17348 80 17368
rect 2467 17116 2476 17156
rect 2516 17116 3820 17156
rect 3860 17116 3869 17156
rect 77731 17116 77740 17156
rect 77780 17116 80620 17156
rect 80660 17116 80669 17156
rect 3427 17032 3436 17072
rect 3476 17032 4972 17072
rect 5012 17032 5021 17072
rect 4003 16864 4012 16904
rect 4052 16864 8021 16904
rect 4675 16696 4684 16736
rect 4724 16696 5836 16736
rect 5876 16696 7756 16736
rect 7796 16696 8021 16736
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 0 16568 80 16588
rect 0 16528 1228 16568
rect 1268 16528 1277 16568
rect 5827 16528 5836 16568
rect 5876 16528 8021 16568
rect 0 16508 80 16528
rect 7747 16360 7756 16400
rect 7796 16360 7948 16400
rect 7988 16360 7997 16400
rect 4579 16192 4588 16232
rect 4628 16192 5068 16232
rect 5108 16192 5836 16232
rect 5876 16192 5885 16232
rect 1123 16024 1132 16064
rect 1172 16024 1900 16064
rect 1940 16024 4012 16064
rect 4052 16024 4061 16064
rect 2851 15940 2860 15980
rect 2900 15940 4780 15980
rect 4820 15940 4829 15980
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 0 15728 80 15748
rect 0 15688 844 15728
rect 884 15688 893 15728
rect 0 15668 80 15688
rect 3427 15520 3436 15560
rect 3476 15520 4972 15560
rect 5012 15520 5021 15560
rect 643 15476 701 15477
rect 558 15436 652 15476
rect 692 15436 701 15476
rect 643 15435 701 15436
rect 1603 15352 1612 15392
rect 1652 15352 2188 15392
rect 2228 15352 2237 15392
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 0 14888 80 14908
rect 0 14848 844 14888
rect 884 14848 893 14888
rect 1795 14848 1804 14888
rect 1844 14848 4012 14888
rect 4052 14848 8021 14888
rect 0 14828 80 14848
rect 1507 14680 1516 14720
rect 1556 14680 3628 14720
rect 3668 14680 4108 14720
rect 4148 14680 4157 14720
rect 4675 14680 4684 14720
rect 4724 14680 5068 14720
rect 5108 14680 5117 14720
rect 1219 14344 1228 14384
rect 1268 14344 1996 14384
rect 2036 14344 2045 14384
rect 3523 14344 3532 14384
rect 3572 14344 3916 14384
rect 3956 14344 3965 14384
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 0 14048 80 14068
rect 0 14008 844 14048
rect 884 14008 893 14048
rect 4003 14008 4012 14048
rect 4052 14008 4780 14048
rect 4820 14008 5836 14048
rect 5876 14008 5885 14048
rect 0 13988 80 14008
rect 1603 13840 1612 13880
rect 1652 13840 2188 13880
rect 2228 13840 2237 13880
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 1219 13336 1228 13376
rect 1268 13336 2956 13376
rect 2996 13336 3820 13376
rect 3860 13336 3869 13376
rect 3427 13252 3436 13292
rect 3476 13252 4300 13292
rect 4340 13252 4349 13292
rect 0 13208 80 13228
rect 0 13168 748 13208
rect 788 13168 797 13208
rect 2083 13168 2092 13208
rect 2132 13168 4684 13208
rect 4724 13168 4733 13208
rect 0 13148 80 13168
rect 835 12832 844 12872
rect 884 12832 2188 12872
rect 2228 12832 2237 12872
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 7660 12821 8040 12861
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 7660 12788 7700 12821
rect 4195 12748 4204 12788
rect 4244 12748 5740 12788
rect 5780 12748 7700 12788
rect 5827 12664 5836 12704
rect 5876 12664 8021 12704
rect 3427 12496 3436 12536
rect 3476 12496 4588 12536
rect 4628 12496 4637 12536
rect 4963 12496 4972 12536
rect 5012 12496 8021 12536
rect 643 12412 652 12452
rect 692 12412 2764 12452
rect 2804 12412 2813 12452
rect 0 12368 80 12388
rect 0 12328 1228 12368
rect 1268 12328 1277 12368
rect 5827 12328 5836 12368
rect 5876 12328 8021 12368
rect 0 12308 80 12328
rect 1891 12244 1900 12284
rect 1940 12244 3244 12284
rect 3284 12244 7700 12284
rect 7660 12242 7700 12244
rect 7660 12202 8040 12242
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 7660 11981 8040 12021
rect 7660 11948 7700 11981
rect 4003 11908 4012 11948
rect 4052 11908 5164 11948
rect 5204 11908 7700 11948
rect 3907 11824 3916 11864
rect 3956 11824 4300 11864
rect 4340 11824 5836 11864
rect 5876 11824 5885 11864
rect 643 11740 652 11780
rect 692 11740 1228 11780
rect 1268 11740 1277 11780
rect 1795 11656 1804 11696
rect 1844 11656 2092 11696
rect 2132 11656 4972 11696
rect 5012 11656 5021 11696
rect 1123 11572 1132 11612
rect 1172 11572 1900 11612
rect 1940 11572 1949 11612
rect 3619 11572 3628 11612
rect 3668 11572 3916 11612
rect 3956 11572 3965 11612
rect 0 11528 80 11548
rect 0 11488 844 11528
rect 884 11488 893 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 1987 10984 1996 11024
rect 2036 10984 3628 11024
rect 3668 10984 3677 11024
rect 3811 10984 3820 11024
rect 3860 10984 4780 11024
rect 4820 10984 4829 11024
rect 643 10900 652 10940
rect 692 10900 1132 10940
rect 1172 10900 1181 10940
rect 835 10732 844 10772
rect 884 10732 893 10772
rect 3811 10732 3820 10772
rect 3860 10732 4108 10772
rect 4148 10732 4157 10772
rect 0 10688 80 10708
rect 844 10688 884 10732
rect 0 10648 884 10688
rect 2179 10648 2188 10688
rect 2228 10648 2476 10688
rect 2516 10648 2525 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 643 10228 652 10268
rect 692 10228 940 10268
rect 980 10228 989 10268
rect 3619 10228 3628 10268
rect 3668 10228 5836 10268
rect 5876 10228 5885 10268
rect 3427 10060 3436 10100
rect 3476 10060 4204 10100
rect 4244 10060 4253 10100
rect 3523 10016 3581 10017
rect 3438 9976 3532 10016
rect 3572 9976 3581 10016
rect 3523 9975 3581 9976
rect 0 9848 80 9868
rect 0 9808 844 9848
rect 884 9808 893 9848
rect 1891 9808 1900 9848
rect 1940 9808 2380 9848
rect 2420 9808 2429 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 0 9788 80 9808
rect 3715 9556 3724 9596
rect 3764 9556 4012 9596
rect 4052 9556 4061 9596
rect 3619 9472 3628 9512
rect 3668 9472 4396 9512
rect 4436 9472 4445 9512
rect 98760 9379 98860 9419
rect 98900 9379 98909 9419
rect 80611 9220 80620 9260
rect 80660 9251 82484 9260
rect 98731 9251 98789 9252
rect 80660 9220 82840 9251
rect 82444 9211 82840 9220
rect 98731 9211 98740 9251
rect 98780 9211 98789 9251
rect 98731 9210 98789 9211
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 82819 9083 82877 9084
rect 82819 9043 82828 9083
rect 82868 9043 82877 9083
rect 82819 9042 82877 9043
rect 98731 9045 98789 9046
rect 0 9008 80 9028
rect 0 8968 844 9008
rect 884 8968 893 9008
rect 98731 9005 98740 9045
rect 98780 9005 98789 9045
rect 98731 9004 98789 9005
rect 0 8948 80 8968
rect 98851 8877 98909 8878
rect 98760 8837 98860 8877
rect 98900 8837 98909 8877
rect 98851 8836 98909 8837
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 0 8168 80 8188
rect 0 8128 748 8168
rect 788 8128 797 8168
rect 0 8108 80 8128
rect 3427 7960 3436 8000
rect 3476 7960 5068 8000
rect 5108 7960 5117 8000
rect 4771 7708 4780 7748
rect 4820 7708 5740 7748
rect 5780 7708 5789 7748
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 0 7328 80 7348
rect 40867 7328 40925 7329
rect 0 7288 844 7328
rect 884 7288 893 7328
rect 40867 7288 40876 7328
rect 40929 7288 41011 7328
rect 0 7268 80 7288
rect 40867 7287 40925 7288
rect 34755 7204 34764 7244
rect 34804 7204 35212 7244
rect 35252 7204 35261 7244
rect 70627 7160 70685 7161
rect 4675 7120 4684 7160
rect 4724 7120 16588 7160
rect 16628 7120 16637 7160
rect 26371 7120 26380 7160
rect 26420 7120 70636 7160
rect 70676 7120 70685 7160
rect 70627 7119 70685 7120
rect 4003 7036 4012 7076
rect 4052 7036 4396 7076
rect 4436 7036 15820 7076
rect 15860 7036 15869 7076
rect 7939 6952 7948 6992
rect 7988 6952 77644 6992
rect 77684 6952 77693 6992
rect 2563 6868 2572 6908
rect 2612 6868 25708 6908
rect 25748 6868 25757 6908
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 5923 6784 5932 6824
rect 5972 6784 23788 6824
rect 23828 6784 23837 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 73315 6656 73373 6657
rect 2275 6616 2284 6656
rect 2324 6616 16396 6656
rect 16436 6616 16445 6656
rect 16579 6616 16588 6656
rect 16628 6616 17164 6656
rect 17204 6616 19948 6656
rect 19988 6616 19997 6656
rect 37123 6616 37132 6656
rect 37172 6616 73324 6656
rect 73364 6616 73373 6656
rect 73315 6615 73373 6616
rect 98947 6656 99005 6657
rect 99920 6656 100000 6676
rect 98947 6616 98956 6656
rect 98996 6616 100000 6656
rect 98947 6615 99005 6616
rect 99920 6596 100000 6616
rect 75523 6572 75581 6573
rect 6403 6532 6412 6572
rect 6452 6532 21196 6572
rect 21236 6532 21245 6572
rect 38851 6532 38860 6572
rect 38900 6532 75532 6572
rect 75572 6532 75581 6572
rect 75523 6531 75581 6532
rect 0 6488 80 6508
rect 0 6448 844 6488
rect 884 6448 893 6488
rect 2755 6448 2764 6488
rect 2804 6448 36364 6488
rect 36404 6448 36413 6488
rect 40771 6448 40780 6488
rect 40820 6448 42892 6488
rect 42932 6448 80236 6488
rect 80276 6448 80285 6488
rect 0 6428 80 6448
rect 82051 6404 82109 6405
rect 78883 6364 78892 6404
rect 78932 6364 82060 6404
rect 82100 6364 82109 6404
rect 82051 6363 82109 6364
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 19939 5944 19948 5984
rect 19988 5944 23980 5984
rect 24020 5944 24029 5984
rect 7843 5776 7852 5816
rect 7892 5776 16876 5816
rect 16916 5776 16925 5816
rect 54595 5732 54653 5733
rect 37507 5692 37516 5732
rect 37556 5692 38668 5732
rect 38708 5692 38717 5732
rect 54510 5692 54604 5732
rect 54644 5692 54653 5732
rect 54595 5691 54653 5692
rect 0 5648 80 5668
rect 0 5608 844 5648
rect 884 5608 893 5648
rect 0 5588 80 5608
rect 30595 5524 30604 5564
rect 30644 5524 33772 5564
rect 33812 5524 33821 5564
rect 547 5440 556 5480
rect 596 5440 17300 5480
rect 28579 5440 28588 5480
rect 28628 5440 34924 5480
rect 34964 5440 34973 5480
rect 17260 5396 17300 5440
rect 68995 5396 69053 5397
rect 2467 5356 2476 5396
rect 2516 5356 12364 5396
rect 12404 5356 12413 5396
rect 17260 5356 37172 5396
rect 37219 5356 37228 5396
rect 37268 5356 37612 5396
rect 37652 5356 37661 5396
rect 41251 5356 41260 5396
rect 41300 5356 69004 5396
rect 69044 5356 69053 5396
rect 8419 5312 8477 5313
rect 37132 5312 37172 5356
rect 68995 5355 69053 5356
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 8419 5272 8428 5312
rect 8468 5272 12500 5312
rect 16963 5272 16972 5312
rect 17012 5272 18412 5312
rect 18452 5272 18461 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 21763 5272 21772 5312
rect 21812 5272 23212 5312
rect 23252 5272 23980 5312
rect 24020 5272 24029 5312
rect 24355 5272 24364 5312
rect 24404 5272 26092 5312
rect 26132 5272 27244 5312
rect 27284 5272 27293 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 37132 5272 39244 5312
rect 39284 5272 39293 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 8419 5271 8477 5272
rect 12460 5228 12500 5272
rect 71491 5228 71549 5229
rect 12460 5188 30604 5228
rect 30644 5188 30653 5228
rect 32140 5188 32716 5228
rect 32756 5188 71500 5228
rect 71540 5188 71549 5228
rect 32140 5144 32180 5188
rect 71491 5187 71549 5188
rect 7075 5104 7084 5144
rect 7124 5104 12212 5144
rect 12355 5104 12364 5144
rect 12404 5104 26572 5144
rect 26612 5104 26621 5144
rect 31939 5104 31948 5144
rect 31988 5104 32140 5144
rect 32180 5104 32189 5144
rect 32323 5104 32332 5144
rect 32372 5104 35980 5144
rect 36020 5104 36940 5144
rect 36980 5104 38572 5144
rect 38612 5104 38621 5144
rect 38755 5104 38764 5144
rect 38804 5104 82732 5144
rect 82772 5104 82781 5144
rect 12172 4976 12212 5104
rect 12172 4936 45196 4976
rect 45236 4936 45245 4976
rect 47107 4936 47116 4976
rect 47156 4936 52108 4976
rect 52148 4936 53644 4976
rect 53684 4936 53693 4976
rect 643 4852 652 4892
rect 692 4852 7220 4892
rect 46819 4852 46828 4892
rect 46868 4852 54604 4892
rect 54644 4852 54653 4892
rect 0 4808 80 4828
rect 0 4768 844 4808
rect 884 4768 893 4808
rect 0 4748 80 4768
rect 7180 4640 7220 4852
rect 8515 4808 8573 4809
rect 8515 4768 8524 4808
rect 8564 4768 17260 4808
rect 17300 4768 18700 4808
rect 18740 4768 18749 4808
rect 25411 4768 25420 4808
rect 25460 4768 26956 4808
rect 26996 4768 27005 4808
rect 27052 4768 32428 4808
rect 32468 4768 32477 4808
rect 38755 4768 38764 4808
rect 38804 4768 39148 4808
rect 39188 4768 39197 4808
rect 39331 4768 39340 4808
rect 39380 4768 40300 4808
rect 40340 4768 40349 4808
rect 8515 4767 8573 4768
rect 27052 4724 27092 4768
rect 68803 4724 68861 4725
rect 10156 4684 21524 4724
rect 21571 4684 21580 4724
rect 21620 4684 22060 4724
rect 22100 4684 22109 4724
rect 23395 4684 23404 4724
rect 23444 4684 24748 4724
rect 24788 4684 24797 4724
rect 25219 4684 25228 4724
rect 25268 4684 26764 4724
rect 26804 4684 26813 4724
rect 26860 4684 27092 4724
rect 27235 4684 27244 4724
rect 27284 4684 28588 4724
rect 28628 4684 28637 4724
rect 29539 4684 29548 4724
rect 29588 4684 30988 4724
rect 31028 4684 31037 4724
rect 38659 4684 38668 4724
rect 38708 4684 38956 4724
rect 38996 4684 39005 4724
rect 43843 4684 43852 4724
rect 43892 4684 68812 4724
rect 68852 4684 68861 4724
rect 10156 4640 10196 4684
rect 21484 4640 21524 4684
rect 7180 4600 10196 4640
rect 15811 4600 15820 4640
rect 15860 4600 16588 4640
rect 16628 4600 20236 4640
rect 20276 4600 21388 4640
rect 21428 4600 21437 4640
rect 21484 4600 21620 4640
rect 22723 4600 22732 4640
rect 22772 4600 24076 4640
rect 24116 4600 25708 4640
rect 25748 4600 25757 4640
rect 21580 4556 21620 4600
rect 26860 4556 26900 4684
rect 68803 4683 68861 4684
rect 27043 4600 27052 4640
rect 27092 4600 35404 4640
rect 35444 4600 35453 4640
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 21580 4516 26900 4556
rect 26947 4516 26956 4556
rect 26996 4516 28012 4556
rect 28052 4516 28061 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 26755 4432 26764 4472
rect 26804 4432 27052 4472
rect 27092 4432 27101 4472
rect 16003 4348 16012 4388
rect 16052 4348 17260 4388
rect 17300 4348 17309 4388
rect 40675 4348 40684 4388
rect 40724 4348 41260 4388
rect 41300 4348 41309 4388
rect 53635 4348 53644 4388
rect 53684 4348 54700 4388
rect 54740 4348 54749 4388
rect 69283 4304 69341 4305
rect 7180 4264 40972 4304
rect 41012 4264 41021 4304
rect 42499 4264 42508 4304
rect 42548 4264 43852 4304
rect 43892 4264 69292 4304
rect 69332 4264 69341 4304
rect 7180 4220 7220 4264
rect 69283 4263 69341 4264
rect 69379 4220 69437 4221
rect 1219 4180 1228 4220
rect 1268 4180 7220 4220
rect 16387 4180 16396 4220
rect 16436 4180 17836 4220
rect 17876 4180 20428 4220
rect 20468 4180 20477 4220
rect 20611 4180 20620 4220
rect 20660 4180 21676 4220
rect 21716 4180 22444 4220
rect 22484 4180 22493 4220
rect 26764 4180 29644 4220
rect 29684 4180 29693 4220
rect 30499 4180 30508 4220
rect 30548 4180 30700 4220
rect 30740 4180 31948 4220
rect 31988 4180 34348 4220
rect 34388 4180 34397 4220
rect 34627 4180 34636 4220
rect 34676 4180 35156 4220
rect 47203 4180 47212 4220
rect 47252 4180 47500 4220
rect 47540 4180 50188 4220
rect 50228 4180 50380 4220
rect 50420 4180 50429 4220
rect 50476 4180 69388 4220
rect 69428 4180 69437 4220
rect 26764 4136 26804 4180
rect 35116 4136 35156 4180
rect 43363 4136 43421 4137
rect 50476 4136 50516 4180
rect 69379 4179 69437 4180
rect 59779 4136 59837 4137
rect 18691 4096 18700 4136
rect 18740 4096 21292 4136
rect 21332 4096 22828 4136
rect 22868 4096 24652 4136
rect 24692 4096 24701 4136
rect 25987 4096 25996 4136
rect 26036 4096 26764 4136
rect 26804 4096 26813 4136
rect 27340 4096 27436 4136
rect 27476 4096 28492 4136
rect 28532 4096 30796 4136
rect 30836 4096 30845 4136
rect 32227 4096 32236 4136
rect 32276 4096 34772 4136
rect 35107 4096 35116 4136
rect 35156 4096 35692 4136
rect 35732 4096 35741 4136
rect 40771 4096 40780 4136
rect 40820 4096 41260 4136
rect 41300 4096 41309 4136
rect 42787 4096 42796 4136
rect 42836 4096 42845 4136
rect 43278 4096 43372 4136
rect 43412 4096 43421 4136
rect 46147 4096 46156 4136
rect 46196 4096 46205 4136
rect 46252 4096 47404 4136
rect 47444 4096 48652 4136
rect 48692 4096 48701 4136
rect 49132 4096 50516 4136
rect 51715 4096 51724 4136
rect 51764 4096 53356 4136
rect 53396 4096 53405 4136
rect 53539 4096 53548 4136
rect 53588 4096 55468 4136
rect 55508 4096 59788 4136
rect 59828 4096 59837 4136
rect 27340 4052 27380 4096
rect 34732 4052 34772 4096
rect 42796 4052 42836 4096
rect 43363 4095 43421 4096
rect 46156 4052 46196 4096
rect 46252 4052 46292 4096
rect 8227 4012 8236 4052
rect 8276 4012 27380 4052
rect 30595 4012 30604 4052
rect 30644 4012 33484 4052
rect 33524 4012 33964 4052
rect 34004 4012 34252 4052
rect 34292 4012 34301 4052
rect 34723 4012 34732 4052
rect 34772 4012 35308 4052
rect 35348 4012 42836 4052
rect 43180 4012 46196 4052
rect 46243 4012 46252 4052
rect 46292 4012 46301 4052
rect 47299 4012 47308 4052
rect 47348 4012 49036 4052
rect 49076 4012 49085 4052
rect 0 3968 80 3988
rect 43180 3968 43220 4012
rect 44515 3968 44573 3969
rect 0 3928 844 3968
rect 884 3928 893 3968
rect 20515 3928 20524 3968
rect 20564 3928 24460 3968
rect 24500 3928 25804 3968
rect 25844 3928 25853 3968
rect 29635 3928 29644 3968
rect 29684 3928 34828 3968
rect 34868 3928 34877 3968
rect 35491 3928 35500 3968
rect 35540 3928 38572 3968
rect 38612 3928 38621 3968
rect 38668 3928 43220 3968
rect 44430 3928 44524 3968
rect 44564 3928 44573 3968
rect 0 3908 80 3928
rect 38668 3884 38708 3928
rect 44515 3927 44573 3928
rect 49132 3884 49172 4096
rect 59779 4095 59837 4096
rect 49219 4012 49228 4052
rect 49268 4012 51820 4052
rect 51860 4012 74668 4052
rect 74708 4012 74717 4052
rect 69187 3968 69245 3969
rect 49411 3928 49420 3968
rect 49460 3928 53740 3968
rect 53780 3928 56620 3968
rect 56660 3928 56669 3968
rect 57580 3928 69196 3968
rect 69236 3928 69245 3968
rect 57580 3884 57620 3928
rect 69187 3927 69245 3928
rect 25699 3844 25708 3884
rect 25748 3844 29356 3884
rect 29396 3844 30220 3884
rect 30260 3844 30269 3884
rect 34243 3844 34252 3884
rect 34292 3844 38708 3884
rect 43171 3844 43180 3884
rect 43220 3844 49172 3884
rect 53347 3844 53356 3884
rect 53396 3844 57620 3884
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49027 3760 49036 3800
rect 49076 3760 49420 3800
rect 49460 3760 49469 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 1315 3676 1324 3716
rect 1364 3676 32524 3716
rect 32564 3676 35116 3716
rect 35156 3676 35165 3716
rect 38467 3676 38476 3716
rect 38516 3676 40876 3716
rect 40916 3676 40925 3716
rect 42307 3676 42316 3716
rect 42356 3676 51724 3716
rect 51764 3676 51773 3716
rect 69475 3632 69533 3633
rect 34819 3592 34828 3632
rect 34868 3592 45140 3632
rect 45187 3592 45196 3632
rect 45236 3592 48076 3632
rect 48116 3592 69484 3632
rect 69524 3592 69533 3632
rect 45100 3548 45140 3592
rect 69475 3591 69533 3592
rect 69091 3548 69149 3549
rect 1027 3508 1036 3548
rect 1076 3508 31700 3548
rect 31747 3508 31756 3548
rect 31796 3508 35116 3548
rect 35156 3508 35165 3548
rect 35212 3508 37324 3548
rect 37364 3508 40108 3548
rect 40148 3508 41300 3548
rect 43075 3508 43084 3548
rect 43124 3508 43948 3548
rect 43988 3508 43997 3548
rect 45100 3508 45388 3548
rect 45428 3508 46060 3548
rect 46100 3508 46109 3548
rect 46156 3508 69100 3548
rect 69140 3508 69149 3548
rect 31660 3464 31700 3508
rect 35212 3464 35252 3508
rect 41260 3464 41300 3508
rect 46156 3464 46196 3508
rect 69091 3507 69149 3508
rect 20419 3424 20428 3464
rect 20468 3424 21964 3464
rect 22004 3424 22252 3464
rect 22292 3424 22301 3464
rect 23779 3424 23788 3464
rect 23828 3424 23980 3464
rect 24020 3424 25900 3464
rect 25940 3424 26572 3464
rect 26612 3424 27628 3464
rect 27668 3424 29932 3464
rect 29972 3424 31468 3464
rect 31508 3424 31517 3464
rect 31660 3424 32236 3464
rect 32276 3424 32285 3464
rect 35011 3424 35020 3464
rect 35060 3424 35212 3464
rect 35252 3424 35261 3464
rect 36931 3424 36940 3464
rect 36980 3424 41068 3464
rect 41108 3424 41117 3464
rect 41251 3424 41260 3464
rect 41300 3424 41309 3464
rect 43267 3424 43276 3464
rect 43316 3424 46196 3464
rect 46915 3424 46924 3464
rect 46964 3424 50188 3464
rect 50228 3424 52012 3464
rect 52052 3424 52972 3464
rect 53012 3424 53021 3464
rect 43276 3380 43316 3424
rect 34915 3340 34924 3380
rect 34964 3340 35308 3380
rect 35348 3340 37036 3380
rect 37076 3340 38380 3380
rect 38420 3340 38860 3380
rect 38900 3340 38909 3380
rect 40003 3340 40012 3380
rect 40052 3340 43316 3380
rect 20035 3256 20044 3296
rect 20084 3256 20908 3296
rect 20948 3256 20957 3296
rect 36739 3256 36748 3296
rect 36788 3256 39916 3296
rect 39956 3256 39965 3296
rect 41059 3256 41068 3296
rect 41108 3256 47404 3296
rect 47444 3256 47453 3296
rect 40963 3172 40972 3212
rect 41012 3172 42220 3212
rect 42260 3172 43180 3212
rect 43220 3172 43229 3212
rect 0 3128 80 3148
rect 0 3088 844 3128
rect 884 3088 893 3128
rect 38275 3088 38284 3128
rect 38324 3088 81964 3128
rect 82004 3088 82013 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 35683 3004 35692 3044
rect 35732 3004 44332 3044
rect 44372 3004 44381 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 1123 2836 1132 2876
rect 1172 2836 32428 2876
rect 32468 2836 32477 2876
rect 39043 2836 39052 2876
rect 39092 2836 40588 2876
rect 40628 2836 41068 2876
rect 41108 2836 41117 2876
rect 46339 2836 46348 2876
rect 46388 2836 47596 2876
rect 47636 2836 49228 2876
rect 49268 2836 49277 2876
rect 2371 2752 2380 2792
rect 2420 2752 34924 2792
rect 34964 2752 34973 2792
rect 35587 2752 35596 2792
rect 35636 2752 35645 2792
rect 38947 2752 38956 2792
rect 38996 2752 40204 2792
rect 40244 2752 40253 2792
rect 45475 2752 45484 2792
rect 45524 2752 46636 2792
rect 46676 2752 47020 2792
rect 47060 2752 48364 2792
rect 48404 2752 49036 2792
rect 49076 2752 50380 2792
rect 50420 2752 50956 2792
rect 50996 2752 52300 2792
rect 52340 2752 52684 2792
rect 52724 2752 52733 2792
rect 23011 2668 23020 2708
rect 23060 2668 23500 2708
rect 23540 2668 24268 2708
rect 24308 2668 24317 2708
rect 26659 2668 26668 2708
rect 26708 2668 28204 2708
rect 28244 2668 28253 2708
rect 29740 2668 31564 2708
rect 31604 2668 34348 2708
rect 34388 2668 34397 2708
rect 29740 2624 29780 2668
rect 28099 2584 28108 2624
rect 28148 2584 29740 2624
rect 29780 2584 29789 2624
rect 31747 2584 31756 2624
rect 31796 2584 32236 2624
rect 32276 2584 32524 2624
rect 32564 2584 32573 2624
rect 21475 2500 21484 2540
rect 21524 2500 26380 2540
rect 26420 2500 27820 2540
rect 27860 2500 31468 2540
rect 31508 2500 31517 2540
rect 931 2416 940 2456
rect 980 2416 31948 2456
rect 31988 2416 31997 2456
rect 32131 2416 32140 2456
rect 32180 2416 32716 2456
rect 32756 2416 32765 2456
rect 35596 2372 35636 2752
rect 47299 2708 47357 2709
rect 37507 2668 37516 2708
rect 37556 2668 42548 2708
rect 45859 2668 45868 2708
rect 45908 2668 47116 2708
rect 47156 2668 47165 2708
rect 47299 2668 47308 2708
rect 47348 2668 49516 2708
rect 49556 2668 51724 2708
rect 51764 2668 52396 2708
rect 52436 2668 52445 2708
rect 36451 2584 36460 2624
rect 36500 2584 38668 2624
rect 38708 2584 40012 2624
rect 40052 2584 40061 2624
rect 40291 2584 40300 2624
rect 40340 2584 42124 2624
rect 42164 2584 42173 2624
rect 42508 2540 42548 2668
rect 47116 2624 47156 2668
rect 47299 2667 47357 2668
rect 47116 2584 47540 2624
rect 51235 2584 51244 2624
rect 51284 2584 51820 2624
rect 51860 2584 51869 2624
rect 47299 2540 47357 2541
rect 36643 2500 36652 2540
rect 36692 2500 39052 2540
rect 39092 2500 39101 2540
rect 40387 2500 40396 2540
rect 40436 2500 42316 2540
rect 42356 2500 42365 2540
rect 42508 2500 47308 2540
rect 47348 2500 47357 2540
rect 47500 2540 47540 2584
rect 47500 2500 47788 2540
rect 47828 2500 49132 2540
rect 49172 2500 49708 2540
rect 49748 2500 51436 2540
rect 51476 2500 51485 2540
rect 47299 2499 47357 2500
rect 28195 2332 28204 2372
rect 28244 2332 30508 2372
rect 30548 2332 35636 2372
rect 0 2288 80 2308
rect 38851 2288 38909 2289
rect 0 2248 844 2288
rect 884 2248 893 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 38851 2248 38860 2288
rect 38900 2248 39340 2288
rect 39380 2248 39389 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 0 2228 80 2248
rect 38851 2247 38909 2248
rect 29635 2164 29644 2204
rect 29684 2164 32428 2204
rect 32468 2164 34156 2204
rect 34196 2164 35884 2204
rect 35924 2164 35933 2204
rect 39139 2164 39148 2204
rect 39188 2164 40300 2204
rect 40340 2164 42892 2204
rect 42932 2164 42941 2204
rect 21763 2080 21772 2120
rect 21812 2080 22732 2120
rect 22772 2080 22781 2120
rect 23107 2080 23116 2120
rect 23156 2080 23596 2120
rect 23636 2080 25996 2120
rect 26036 2080 26045 2120
rect 31651 2080 31660 2120
rect 31700 2080 57620 2120
rect 57580 2036 57620 2080
rect 22147 1996 22156 2036
rect 22196 1996 23020 2036
rect 23060 1996 23069 2036
rect 34723 1996 34732 2036
rect 34772 1996 35404 2036
rect 35444 1996 37324 2036
rect 37364 1996 37373 2036
rect 39907 1996 39916 2036
rect 39956 1996 40684 2036
rect 40724 1996 40733 2036
rect 49891 1996 49900 2036
rect 49940 1996 51244 2036
rect 51284 1996 51293 2036
rect 57580 1996 91353 2036
rect 8323 1912 8332 1952
rect 8372 1912 24844 1952
rect 24884 1912 27380 1952
rect 30787 1912 30796 1952
rect 30836 1912 33004 1952
rect 33044 1912 35596 1952
rect 35636 1912 38188 1952
rect 38228 1912 38237 1952
rect 41155 1912 41164 1952
rect 41204 1912 43756 1952
rect 43796 1912 74092 1952
rect 74132 1912 74141 1952
rect 81955 1912 81964 1952
rect 82004 1912 90932 1952
rect 27340 1868 27380 1912
rect 27340 1828 27436 1868
rect 27476 1828 29356 1868
rect 29396 1828 30412 1868
rect 30452 1828 32332 1868
rect 32372 1828 40012 1868
rect 40052 1828 40061 1868
rect 36547 1744 36556 1784
rect 36596 1744 36748 1784
rect 36788 1744 36797 1784
rect 37315 1744 37324 1784
rect 37364 1744 39148 1784
rect 39188 1744 39197 1784
rect 47299 1744 47308 1784
rect 47348 1744 48172 1784
rect 48212 1744 51052 1784
rect 51092 1744 51101 1784
rect 26083 1660 26092 1700
rect 26132 1660 28628 1700
rect 28588 1616 28628 1660
rect 28579 1576 28588 1616
rect 28628 1576 40204 1616
rect 40244 1576 40253 1616
rect 43363 1576 43372 1616
rect 43412 1576 90644 1616
rect 38851 1532 38909 1533
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 28003 1492 28012 1532
rect 28052 1492 28492 1532
rect 28532 1492 29548 1532
rect 29588 1492 32140 1532
rect 32180 1492 32189 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 35683 1492 35692 1532
rect 35732 1492 35980 1532
rect 36020 1492 36029 1532
rect 36835 1492 36844 1532
rect 36884 1492 38860 1532
rect 38900 1492 38909 1532
rect 42403 1492 42412 1532
rect 42452 1492 44428 1532
rect 44468 1492 45868 1532
rect 45908 1492 45917 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 38851 1491 38909 1492
rect 90604 1479 90644 1576
rect 90892 1479 90932 1912
rect 91313 1479 91353 1996
rect 32707 1408 32716 1448
rect 32756 1408 37460 1448
rect 90604 1439 90737 1479
rect 90777 1439 90786 1479
rect 90892 1439 91121 1479
rect 91161 1439 91170 1479
rect 91304 1439 91313 1479
rect 91353 1439 91362 1479
rect 37420 1364 37460 1408
rect 34339 1324 34348 1364
rect 34388 1324 34828 1364
rect 34868 1324 34877 1364
rect 37420 1324 67700 1364
rect 67660 1280 67700 1324
rect 34435 1240 34444 1280
rect 34484 1240 39724 1280
rect 39764 1240 44812 1280
rect 44852 1240 47500 1280
rect 47540 1240 47549 1280
rect 67660 1240 90537 1280
rect 90577 1240 90586 1280
rect 31555 1156 31564 1196
rect 31604 1156 34156 1196
rect 34196 1156 36460 1196
rect 36500 1156 36652 1196
rect 36692 1156 36701 1196
rect 39619 1156 39628 1196
rect 39668 1156 42508 1196
rect 42548 1156 51820 1196
rect 51860 1156 54412 1196
rect 54452 1156 54461 1196
rect 31843 1072 31852 1112
rect 31892 1072 34540 1112
rect 34580 1072 36556 1112
rect 36596 1072 36605 1112
rect 38755 1072 38764 1112
rect 38804 1072 39244 1112
rect 39284 1072 39293 1112
rect 40483 1072 40492 1112
rect 40532 1072 42604 1112
rect 42644 1072 44716 1112
rect 44756 1072 44908 1112
rect 44948 1072 44957 1112
rect 87820 988 90892 1028
rect 90932 988 90941 1028
rect 87820 944 87860 988
rect 35875 904 35884 944
rect 35924 904 87860 944
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 71980 36436 72020 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 70636 36016 70676 36056
rect 71980 36016 72020 36056
rect 24268 35764 24308 35804
rect 69196 35680 69236 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 69100 35512 69140 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 41164 35344 41204 35384
rect 12268 35092 12308 35132
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 8428 34084 8468 34124
rect 61036 34084 61076 34124
rect 69484 34084 69524 34124
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 68812 33832 68852 33872
rect 69388 33664 69428 33704
rect 69292 33496 69332 33536
rect 72652 33328 72692 33368
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 99820 33160 99860 33200
rect 12268 33076 12308 33116
rect 69004 32824 69044 32864
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 8524 32404 8564 32444
rect 60748 32404 60788 32444
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 83500 30052 83540 30092
rect 97324 30051 97364 30091
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 97324 29021 97364 29061
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 84940 25936 84980 25976
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 82924 23752 82964 23792
rect 99916 23752 99956 23792
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 652 15436 692 15476
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 3532 9976 3572 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 98740 9211 98780 9251
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 82828 9043 82868 9083
rect 98740 9005 98780 9045
rect 98860 8837 98900 8877
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 40876 7288 40889 7328
rect 40889 7288 40916 7328
rect 70636 7120 70676 7160
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 73324 6616 73364 6656
rect 98956 6616 98996 6656
rect 75532 6532 75572 6572
rect 82060 6364 82100 6404
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 54604 5692 54644 5732
rect 69004 5356 69044 5396
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8428 5272 8468 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 71500 5188 71540 5228
rect 8524 4768 8564 4808
rect 68812 4684 68852 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 69292 4264 69332 4304
rect 69388 4180 69428 4220
rect 43372 4096 43412 4136
rect 59788 4096 59828 4136
rect 44524 3928 44564 3968
rect 69196 3928 69236 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 69484 3592 69524 3632
rect 69100 3508 69140 3548
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 47308 2668 47348 2708
rect 47308 2500 47348 2540
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 38860 2248 38900 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 38860 1492 38900 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 71980 36476 72020 36485
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 70636 36056 70676 36065
rect 24268 35804 24308 35813
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 24268 35225 24308 35764
rect 69196 35720 69236 35729
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 69100 35552 69140 35561
rect 41164 35384 41204 35393
rect 41164 35225 41204 35344
rect 24267 35216 24309 35225
rect 24267 35176 24268 35216
rect 24308 35176 24309 35216
rect 24267 35167 24309 35176
rect 41163 35216 41205 35225
rect 41163 35176 41164 35216
rect 41204 35176 41205 35216
rect 41163 35167 41205 35176
rect 12267 35132 12309 35141
rect 12267 35092 12268 35132
rect 12308 35092 12309 35132
rect 12267 35083 12309 35092
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 8428 34124 8468 34133
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 652 15476 692 15485
rect 652 3977 692 15436
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3532 10016 3572 10025
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3532 7841 3572 9976
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 3531 7832 3573 7841
rect 3531 7792 3532 7832
rect 3572 7792 3573 7832
rect 3531 7783 3573 7792
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 8428 5312 8468 34084
rect 12268 33116 12308 35083
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 61036 34124 61076 34133
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 61036 33881 61076 34084
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 61035 33872 61077 33881
rect 61035 33832 61036 33872
rect 61076 33832 61077 33872
rect 61035 33823 61077 33832
rect 68812 33872 68852 33881
rect 12268 33067 12308 33076
rect 8428 5263 8468 5272
rect 8524 32444 8564 32453
rect 8524 4808 8564 32404
rect 60748 32444 60788 32453
rect 60748 30017 60788 32404
rect 60747 30008 60789 30017
rect 60747 29968 60748 30008
rect 60788 29968 60789 30008
rect 60747 29959 60789 29968
rect 38859 7832 38901 7841
rect 38859 7792 38860 7832
rect 38900 7792 38901 7832
rect 38859 7783 38901 7792
rect 40875 7832 40917 7841
rect 40875 7792 40876 7832
rect 40916 7792 40917 7832
rect 40875 7783 40917 7792
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 8524 4759 8564 4768
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 38860 2288 38900 7783
rect 40876 7328 40916 7783
rect 40876 7279 40916 7288
rect 54603 5732 54645 5741
rect 54603 5692 54604 5732
rect 54644 5692 54645 5732
rect 54603 5683 54645 5692
rect 54604 5598 54644 5683
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 59787 4724 59829 4733
rect 59787 4684 59788 4724
rect 59828 4684 59829 4724
rect 59787 4675 59829 4684
rect 68812 4724 68852 33832
rect 69004 32864 69044 32873
rect 69004 5396 69044 32824
rect 69004 5347 69044 5356
rect 68812 4675 68852 4684
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 43371 4136 43413 4145
rect 43371 4096 43372 4136
rect 43412 4096 43413 4136
rect 43371 4087 43413 4096
rect 59788 4136 59828 4675
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 59788 4087 59828 4096
rect 43372 4002 43412 4087
rect 44523 3968 44565 3977
rect 44523 3928 44524 3968
rect 44564 3928 44565 3968
rect 44523 3919 44565 3928
rect 44524 3834 44564 3919
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 69100 3548 69140 35512
rect 69196 3968 69236 35680
rect 69484 34124 69524 34133
rect 69388 33704 69428 33713
rect 69292 33536 69332 33545
rect 69292 4304 69332 33496
rect 69292 4255 69332 4264
rect 69388 4220 69428 33664
rect 69388 4171 69428 4180
rect 69196 3919 69236 3928
rect 69484 3632 69524 34084
rect 70636 7160 70676 36016
rect 71980 36056 72020 36436
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 71980 36007 72020 36016
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 72652 33368 72692 33377
rect 71499 7916 71541 7925
rect 71499 7876 71500 7916
rect 71540 7876 71541 7916
rect 71499 7867 71541 7876
rect 70636 7111 70676 7120
rect 71500 5228 71540 7867
rect 71500 5179 71540 5188
rect 72652 4145 72692 33328
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 99820 33200 99860 33209
rect 99860 33160 99956 33200
rect 99820 33151 99860 33160
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 83499 30344 83541 30353
rect 83499 30304 83500 30344
rect 83540 30304 83541 30344
rect 83499 30295 83541 30304
rect 97323 30344 97365 30353
rect 97323 30304 97324 30344
rect 97364 30304 97365 30344
rect 97323 30295 97365 30304
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 83500 30092 83540 30295
rect 83500 30043 83540 30052
rect 97324 30091 97364 30295
rect 97324 30042 97364 30051
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 97324 29061 97364 29070
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 97324 28421 97364 29021
rect 84939 28412 84981 28421
rect 84939 28372 84940 28412
rect 84980 28372 84981 28412
rect 84939 28363 84981 28372
rect 97323 28412 97365 28421
rect 97323 28372 97324 28412
rect 97364 28372 97365 28412
rect 97323 28363 97365 28372
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 84940 25976 84980 28363
rect 84940 25927 84980 25936
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 82924 23792 82964 23801
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 82924 17300 82964 23752
rect 99916 23792 99956 33160
rect 99916 23743 99956 23752
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 82828 17260 82964 17300
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 73323 9260 73365 9269
rect 73323 9220 73324 9260
rect 73364 9220 73365 9260
rect 73323 9211 73365 9220
rect 73324 6656 73364 9211
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 82828 9083 82868 17260
rect 98740 9269 98780 9346
rect 98739 9260 98781 9269
rect 98739 9211 98740 9260
rect 98780 9211 98781 9260
rect 98740 9202 98780 9211
rect 82828 9034 82868 9043
rect 98740 9045 98780 9054
rect 98740 8933 98780 9005
rect 75531 8924 75573 8933
rect 75531 8884 75532 8924
rect 75572 8884 75573 8924
rect 75531 8875 75573 8884
rect 98739 8924 98781 8933
rect 98739 8884 98740 8924
rect 98780 8884 98781 8924
rect 98739 8875 98781 8884
rect 98860 8877 98900 8886
rect 73324 6607 73364 6616
rect 75532 6572 75572 8875
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 98860 7925 98900 8837
rect 98859 7916 98901 7925
rect 98859 7876 98860 7916
rect 98900 7876 98901 7916
rect 98859 7867 98901 7876
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 82059 6656 82101 6665
rect 82059 6616 82060 6656
rect 82100 6616 82101 6656
rect 82059 6607 82101 6616
rect 98955 6656 98997 6665
rect 98955 6616 98956 6656
rect 98996 6616 98997 6656
rect 98955 6607 98997 6616
rect 75532 6523 75572 6532
rect 82060 6404 82100 6607
rect 98956 6522 98996 6607
rect 82060 6355 82100 6364
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 72651 4136 72693 4145
rect 72651 4096 72652 4136
rect 72692 4096 72693 4136
rect 72651 4087 72693 4096
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 69484 3583 69524 3592
rect 69100 3499 69140 3508
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 47308 2708 47348 2717
rect 47308 2540 47348 2668
rect 47308 2491 47348 2500
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 38860 1532 38900 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 38860 1483 38900 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 24268 35176 24308 35216
rect 41164 35176 41204 35216
rect 12268 35092 12308 35132
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3532 7792 3572 7832
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 61036 33832 61076 33872
rect 60748 29968 60788 30008
rect 38860 7792 38900 7832
rect 40876 7792 40916 7832
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 652 3928 692 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 54604 5692 54644 5732
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 59788 4684 59828 4724
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 43372 4096 43412 4136
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 44524 3928 44564 3968
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 71500 7876 71540 7916
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 83500 30304 83540 30344
rect 97324 30304 97364 30344
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 84940 28372 84980 28412
rect 97324 28372 97364 28412
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 73324 9220 73364 9260
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 98740 9251 98780 9260
rect 98740 9220 98780 9251
rect 75532 8884 75572 8924
rect 98740 8884 98780 8924
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 98860 7876 98900 7916
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 82060 6616 82100 6656
rect 98956 6616 98996 6656
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 72652 4096 72692 4136
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal5 >>
rect 4343 38576 4390 38618
rect 4514 38576 4558 38618
rect 4682 38576 4729 38618
rect 4343 38536 4352 38576
rect 4514 38536 4516 38576
rect 4556 38536 4558 38576
rect 4720 38536 4729 38576
rect 4343 38494 4390 38536
rect 4514 38494 4558 38536
rect 4682 38494 4729 38536
rect 19463 38576 19510 38618
rect 19634 38576 19678 38618
rect 19802 38576 19849 38618
rect 19463 38536 19472 38576
rect 19634 38536 19636 38576
rect 19676 38536 19678 38576
rect 19840 38536 19849 38576
rect 19463 38494 19510 38536
rect 19634 38494 19678 38536
rect 19802 38494 19849 38536
rect 34583 38576 34630 38618
rect 34754 38576 34798 38618
rect 34922 38576 34969 38618
rect 34583 38536 34592 38576
rect 34754 38536 34756 38576
rect 34796 38536 34798 38576
rect 34960 38536 34969 38576
rect 34583 38494 34630 38536
rect 34754 38494 34798 38536
rect 34922 38494 34969 38536
rect 49703 38576 49750 38618
rect 49874 38576 49918 38618
rect 50042 38576 50089 38618
rect 49703 38536 49712 38576
rect 49874 38536 49876 38576
rect 49916 38536 49918 38576
rect 50080 38536 50089 38576
rect 49703 38494 49750 38536
rect 49874 38494 49918 38536
rect 50042 38494 50089 38536
rect 64823 38576 64870 38618
rect 64994 38576 65038 38618
rect 65162 38576 65209 38618
rect 64823 38536 64832 38576
rect 64994 38536 64996 38576
rect 65036 38536 65038 38576
rect 65200 38536 65209 38576
rect 64823 38494 64870 38536
rect 64994 38494 65038 38536
rect 65162 38494 65209 38536
rect 79943 38576 79990 38618
rect 80114 38576 80158 38618
rect 80282 38576 80329 38618
rect 79943 38536 79952 38576
rect 80114 38536 80116 38576
rect 80156 38536 80158 38576
rect 80320 38536 80329 38576
rect 79943 38494 79990 38536
rect 80114 38494 80158 38536
rect 80282 38494 80329 38536
rect 3103 37820 3150 37862
rect 3274 37820 3318 37862
rect 3442 37820 3489 37862
rect 3103 37780 3112 37820
rect 3274 37780 3276 37820
rect 3316 37780 3318 37820
rect 3480 37780 3489 37820
rect 3103 37738 3150 37780
rect 3274 37738 3318 37780
rect 3442 37738 3489 37780
rect 18223 37820 18270 37862
rect 18394 37820 18438 37862
rect 18562 37820 18609 37862
rect 18223 37780 18232 37820
rect 18394 37780 18396 37820
rect 18436 37780 18438 37820
rect 18600 37780 18609 37820
rect 18223 37738 18270 37780
rect 18394 37738 18438 37780
rect 18562 37738 18609 37780
rect 33343 37820 33390 37862
rect 33514 37820 33558 37862
rect 33682 37820 33729 37862
rect 33343 37780 33352 37820
rect 33514 37780 33516 37820
rect 33556 37780 33558 37820
rect 33720 37780 33729 37820
rect 33343 37738 33390 37780
rect 33514 37738 33558 37780
rect 33682 37738 33729 37780
rect 48463 37820 48510 37862
rect 48634 37820 48678 37862
rect 48802 37820 48849 37862
rect 48463 37780 48472 37820
rect 48634 37780 48636 37820
rect 48676 37780 48678 37820
rect 48840 37780 48849 37820
rect 48463 37738 48510 37780
rect 48634 37738 48678 37780
rect 48802 37738 48849 37780
rect 63583 37820 63630 37862
rect 63754 37820 63798 37862
rect 63922 37820 63969 37862
rect 63583 37780 63592 37820
rect 63754 37780 63756 37820
rect 63796 37780 63798 37820
rect 63960 37780 63969 37820
rect 63583 37738 63630 37780
rect 63754 37738 63798 37780
rect 63922 37738 63969 37780
rect 78703 37820 78750 37862
rect 78874 37820 78918 37862
rect 79042 37820 79089 37862
rect 78703 37780 78712 37820
rect 78874 37780 78876 37820
rect 78916 37780 78918 37820
rect 79080 37780 79089 37820
rect 78703 37738 78750 37780
rect 78874 37738 78918 37780
rect 79042 37738 79089 37780
rect 4343 37064 4390 37106
rect 4514 37064 4558 37106
rect 4682 37064 4729 37106
rect 4343 37024 4352 37064
rect 4514 37024 4516 37064
rect 4556 37024 4558 37064
rect 4720 37024 4729 37064
rect 4343 36982 4390 37024
rect 4514 36982 4558 37024
rect 4682 36982 4729 37024
rect 19463 37064 19510 37106
rect 19634 37064 19678 37106
rect 19802 37064 19849 37106
rect 19463 37024 19472 37064
rect 19634 37024 19636 37064
rect 19676 37024 19678 37064
rect 19840 37024 19849 37064
rect 19463 36982 19510 37024
rect 19634 36982 19678 37024
rect 19802 36982 19849 37024
rect 34583 37064 34630 37106
rect 34754 37064 34798 37106
rect 34922 37064 34969 37106
rect 34583 37024 34592 37064
rect 34754 37024 34756 37064
rect 34796 37024 34798 37064
rect 34960 37024 34969 37064
rect 34583 36982 34630 37024
rect 34754 36982 34798 37024
rect 34922 36982 34969 37024
rect 49703 37064 49750 37106
rect 49874 37064 49918 37106
rect 50042 37064 50089 37106
rect 49703 37024 49712 37064
rect 49874 37024 49876 37064
rect 49916 37024 49918 37064
rect 50080 37024 50089 37064
rect 49703 36982 49750 37024
rect 49874 36982 49918 37024
rect 50042 36982 50089 37024
rect 64823 37064 64870 37106
rect 64994 37064 65038 37106
rect 65162 37064 65209 37106
rect 64823 37024 64832 37064
rect 64994 37024 64996 37064
rect 65036 37024 65038 37064
rect 65200 37024 65209 37064
rect 64823 36982 64870 37024
rect 64994 36982 65038 37024
rect 65162 36982 65209 37024
rect 79943 37064 79990 37106
rect 80114 37064 80158 37106
rect 80282 37064 80329 37106
rect 79943 37024 79952 37064
rect 80114 37024 80116 37064
rect 80156 37024 80158 37064
rect 80320 37024 80329 37064
rect 79943 36982 79990 37024
rect 80114 36982 80158 37024
rect 80282 36982 80329 37024
rect 3103 36308 3150 36350
rect 3274 36308 3318 36350
rect 3442 36308 3489 36350
rect 3103 36268 3112 36308
rect 3274 36268 3276 36308
rect 3316 36268 3318 36308
rect 3480 36268 3489 36308
rect 3103 36226 3150 36268
rect 3274 36226 3318 36268
rect 3442 36226 3489 36268
rect 18223 36308 18270 36350
rect 18394 36308 18438 36350
rect 18562 36308 18609 36350
rect 18223 36268 18232 36308
rect 18394 36268 18396 36308
rect 18436 36268 18438 36308
rect 18600 36268 18609 36308
rect 18223 36226 18270 36268
rect 18394 36226 18438 36268
rect 18562 36226 18609 36268
rect 33343 36308 33390 36350
rect 33514 36308 33558 36350
rect 33682 36308 33729 36350
rect 33343 36268 33352 36308
rect 33514 36268 33516 36308
rect 33556 36268 33558 36308
rect 33720 36268 33729 36308
rect 33343 36226 33390 36268
rect 33514 36226 33558 36268
rect 33682 36226 33729 36268
rect 48463 36308 48510 36350
rect 48634 36308 48678 36350
rect 48802 36308 48849 36350
rect 48463 36268 48472 36308
rect 48634 36268 48636 36308
rect 48676 36268 48678 36308
rect 48840 36268 48849 36308
rect 48463 36226 48510 36268
rect 48634 36226 48678 36268
rect 48802 36226 48849 36268
rect 63583 36308 63630 36350
rect 63754 36308 63798 36350
rect 63922 36308 63969 36350
rect 63583 36268 63592 36308
rect 63754 36268 63756 36308
rect 63796 36268 63798 36308
rect 63960 36268 63969 36308
rect 63583 36226 63630 36268
rect 63754 36226 63798 36268
rect 63922 36226 63969 36268
rect 78703 36308 78750 36350
rect 78874 36308 78918 36350
rect 79042 36308 79089 36350
rect 78703 36268 78712 36308
rect 78874 36268 78876 36308
rect 78916 36268 78918 36308
rect 79080 36268 79089 36308
rect 78703 36226 78750 36268
rect 78874 36226 78918 36268
rect 79042 36226 79089 36268
rect 4343 35552 4390 35594
rect 4514 35552 4558 35594
rect 4682 35552 4729 35594
rect 4343 35512 4352 35552
rect 4514 35512 4516 35552
rect 4556 35512 4558 35552
rect 4720 35512 4729 35552
rect 4343 35470 4390 35512
rect 4514 35470 4558 35512
rect 4682 35470 4729 35512
rect 19463 35552 19510 35594
rect 19634 35552 19678 35594
rect 19802 35552 19849 35594
rect 19463 35512 19472 35552
rect 19634 35512 19636 35552
rect 19676 35512 19678 35552
rect 19840 35512 19849 35552
rect 19463 35470 19510 35512
rect 19634 35470 19678 35512
rect 19802 35470 19849 35512
rect 34583 35552 34630 35594
rect 34754 35552 34798 35594
rect 34922 35552 34969 35594
rect 34583 35512 34592 35552
rect 34754 35512 34756 35552
rect 34796 35512 34798 35552
rect 34960 35512 34969 35552
rect 34583 35470 34630 35512
rect 34754 35470 34798 35512
rect 34922 35470 34969 35512
rect 49703 35552 49750 35594
rect 49874 35552 49918 35594
rect 50042 35552 50089 35594
rect 49703 35512 49712 35552
rect 49874 35512 49876 35552
rect 49916 35512 49918 35552
rect 50080 35512 50089 35552
rect 49703 35470 49750 35512
rect 49874 35470 49918 35512
rect 50042 35470 50089 35512
rect 64823 35552 64870 35594
rect 64994 35552 65038 35594
rect 65162 35552 65209 35594
rect 64823 35512 64832 35552
rect 64994 35512 64996 35552
rect 65036 35512 65038 35552
rect 65200 35512 65209 35552
rect 64823 35470 64870 35512
rect 64994 35470 65038 35512
rect 65162 35470 65209 35512
rect 79943 35552 79990 35594
rect 80114 35552 80158 35594
rect 80282 35552 80329 35594
rect 79943 35512 79952 35552
rect 80114 35512 80116 35552
rect 80156 35512 80158 35552
rect 80320 35512 80329 35552
rect 79943 35470 79990 35512
rect 80114 35470 80158 35512
rect 80282 35470 80329 35512
rect 23020 35176 24268 35216
rect 24308 35176 41164 35216
rect 41204 35176 41213 35216
rect 23020 35132 23060 35176
rect 12259 35092 12268 35132
rect 12308 35092 23060 35132
rect 3103 34796 3150 34838
rect 3274 34796 3318 34838
rect 3442 34796 3489 34838
rect 3103 34756 3112 34796
rect 3274 34756 3276 34796
rect 3316 34756 3318 34796
rect 3480 34756 3489 34796
rect 3103 34714 3150 34756
rect 3274 34714 3318 34756
rect 3442 34714 3489 34756
rect 18223 34796 18270 34838
rect 18394 34796 18438 34838
rect 18562 34796 18609 34838
rect 18223 34756 18232 34796
rect 18394 34756 18396 34796
rect 18436 34756 18438 34796
rect 18600 34756 18609 34796
rect 18223 34714 18270 34756
rect 18394 34714 18438 34756
rect 18562 34714 18609 34756
rect 33343 34796 33390 34838
rect 33514 34796 33558 34838
rect 33682 34796 33729 34838
rect 33343 34756 33352 34796
rect 33514 34756 33516 34796
rect 33556 34756 33558 34796
rect 33720 34756 33729 34796
rect 33343 34714 33390 34756
rect 33514 34714 33558 34756
rect 33682 34714 33729 34756
rect 48463 34796 48510 34838
rect 48634 34796 48678 34838
rect 48802 34796 48849 34838
rect 48463 34756 48472 34796
rect 48634 34756 48636 34796
rect 48676 34756 48678 34796
rect 48840 34756 48849 34796
rect 48463 34714 48510 34756
rect 48634 34714 48678 34756
rect 48802 34714 48849 34756
rect 63583 34796 63630 34838
rect 63754 34796 63798 34838
rect 63922 34796 63969 34838
rect 63583 34756 63592 34796
rect 63754 34756 63756 34796
rect 63796 34756 63798 34796
rect 63960 34756 63969 34796
rect 63583 34714 63630 34756
rect 63754 34714 63798 34756
rect 63922 34714 63969 34756
rect 78703 34796 78750 34838
rect 78874 34796 78918 34838
rect 79042 34796 79089 34838
rect 78703 34756 78712 34796
rect 78874 34756 78876 34796
rect 78916 34756 78918 34796
rect 79080 34756 79089 34796
rect 78703 34714 78750 34756
rect 78874 34714 78918 34756
rect 79042 34714 79089 34756
rect 93796 34222 94236 34296
rect 93796 34098 93870 34222
rect 93994 34098 94038 34222
rect 94162 34098 94236 34222
rect 4343 34040 4390 34082
rect 4514 34040 4558 34082
rect 4682 34040 4729 34082
rect 4343 34000 4352 34040
rect 4514 34000 4516 34040
rect 4556 34000 4558 34040
rect 4720 34000 4729 34040
rect 4343 33958 4390 34000
rect 4514 33958 4558 34000
rect 4682 33958 4729 34000
rect 19463 34040 19510 34082
rect 19634 34040 19678 34082
rect 19802 34040 19849 34082
rect 19463 34000 19472 34040
rect 19634 34000 19636 34040
rect 19676 34000 19678 34040
rect 19840 34000 19849 34040
rect 19463 33958 19510 34000
rect 19634 33958 19678 34000
rect 19802 33958 19849 34000
rect 34583 34040 34630 34082
rect 34754 34040 34798 34082
rect 34922 34040 34969 34082
rect 34583 34000 34592 34040
rect 34754 34000 34756 34040
rect 34796 34000 34798 34040
rect 34960 34000 34969 34040
rect 34583 33958 34630 34000
rect 34754 33958 34798 34000
rect 34922 33958 34969 34000
rect 49703 34040 49750 34082
rect 49874 34040 49918 34082
rect 50042 34040 50089 34082
rect 49703 34000 49712 34040
rect 49874 34000 49876 34040
rect 49916 34000 49918 34040
rect 50080 34000 50089 34040
rect 49703 33958 49750 34000
rect 49874 33958 49918 34000
rect 50042 33958 50089 34000
rect 64823 34040 64870 34082
rect 64994 34040 65038 34082
rect 65162 34040 65209 34082
rect 64823 34000 64832 34040
rect 64994 34000 64996 34040
rect 65036 34000 65038 34040
rect 65200 34000 65209 34040
rect 64823 33958 64870 34000
rect 64994 33958 65038 34000
rect 65162 33958 65209 34000
rect 79943 34040 79990 34082
rect 80114 34040 80158 34082
rect 80282 34040 80329 34082
rect 79943 34000 79952 34040
rect 80114 34000 80116 34040
rect 80156 34000 80158 34040
rect 80320 34000 80329 34040
rect 79943 33958 79990 34000
rect 80114 33958 80158 34000
rect 80282 33958 80329 34000
rect 93796 34054 94236 34098
rect 93796 33930 93870 34054
rect 93994 33930 94038 34054
rect 94162 33930 94236 34054
rect 61027 33832 61036 33872
rect 61076 33832 67298 33872
rect 93796 33856 94236 33930
rect 3103 33284 3150 33326
rect 3274 33284 3318 33326
rect 3442 33284 3489 33326
rect 3103 33244 3112 33284
rect 3274 33244 3276 33284
rect 3316 33244 3318 33284
rect 3480 33244 3489 33284
rect 3103 33202 3150 33244
rect 3274 33202 3318 33244
rect 3442 33202 3489 33244
rect 78703 33284 78750 33326
rect 78874 33284 78918 33326
rect 79042 33284 79089 33326
rect 78703 33244 78712 33284
rect 78874 33244 78876 33284
rect 78916 33244 78918 33284
rect 79080 33244 79089 33284
rect 78703 33202 78750 33244
rect 78874 33202 78918 33244
rect 79042 33202 79089 33244
rect 4343 32528 4390 32570
rect 4514 32528 4558 32570
rect 4682 32528 4729 32570
rect 4343 32488 4352 32528
rect 4514 32488 4516 32528
rect 4556 32488 4558 32528
rect 4720 32488 4729 32528
rect 4343 32446 4390 32488
rect 4514 32446 4558 32488
rect 4682 32446 4729 32488
rect 79943 32528 79990 32570
rect 80114 32528 80158 32570
rect 80282 32528 80329 32570
rect 79943 32488 79952 32528
rect 80114 32488 80116 32528
rect 80156 32488 80158 32528
rect 80320 32488 80329 32528
rect 79943 32446 79990 32488
rect 80114 32446 80158 32488
rect 80282 32446 80329 32488
rect 3103 31772 3150 31814
rect 3274 31772 3318 31814
rect 3442 31772 3489 31814
rect 3103 31732 3112 31772
rect 3274 31732 3276 31772
rect 3316 31732 3318 31772
rect 3480 31732 3489 31772
rect 3103 31690 3150 31732
rect 3274 31690 3318 31732
rect 3442 31690 3489 31732
rect 78703 31772 78750 31814
rect 78874 31772 78918 31814
rect 79042 31772 79089 31814
rect 78703 31732 78712 31772
rect 78874 31732 78876 31772
rect 78916 31732 78918 31772
rect 79080 31732 79089 31772
rect 78703 31690 78750 31732
rect 78874 31690 78918 31732
rect 79042 31690 79089 31732
rect 4343 31016 4390 31058
rect 4514 31016 4558 31058
rect 4682 31016 4729 31058
rect 4343 30976 4352 31016
rect 4514 30976 4516 31016
rect 4556 30976 4558 31016
rect 4720 30976 4729 31016
rect 4343 30934 4390 30976
rect 4514 30934 4558 30976
rect 4682 30934 4729 30976
rect 79943 31016 79990 31058
rect 80114 31016 80158 31058
rect 80282 31016 80329 31058
rect 79943 30976 79952 31016
rect 80114 30976 80116 31016
rect 80156 30976 80158 31016
rect 80320 30976 80329 31016
rect 79943 30934 79990 30976
rect 80114 30934 80158 30976
rect 80282 30934 80329 30976
rect 83491 30304 83500 30344
rect 83540 30304 97324 30344
rect 97364 30304 97373 30344
rect 3103 30260 3150 30302
rect 3274 30260 3318 30302
rect 3442 30260 3489 30302
rect 3103 30220 3112 30260
rect 3274 30220 3276 30260
rect 3316 30220 3318 30260
rect 3480 30220 3489 30260
rect 3103 30178 3150 30220
rect 3274 30178 3318 30220
rect 3442 30178 3489 30220
rect 78703 30260 78750 30302
rect 78874 30260 78918 30302
rect 79042 30260 79089 30302
rect 78703 30220 78712 30260
rect 78874 30220 78876 30260
rect 78916 30220 78918 30260
rect 79080 30220 79089 30260
rect 78703 30178 78750 30220
rect 78874 30178 78918 30220
rect 79042 30178 79089 30220
rect 60739 29968 60748 30008
rect 60788 29968 66386 30008
rect 4343 29504 4390 29546
rect 4514 29504 4558 29546
rect 4682 29504 4729 29546
rect 4343 29464 4352 29504
rect 4514 29464 4516 29504
rect 4556 29464 4558 29504
rect 4720 29464 4729 29504
rect 4343 29422 4390 29464
rect 4514 29422 4558 29464
rect 4682 29422 4729 29464
rect 79943 29504 79990 29546
rect 80114 29504 80158 29546
rect 80282 29504 80329 29546
rect 79943 29464 79952 29504
rect 80114 29464 80116 29504
rect 80156 29464 80158 29504
rect 80320 29464 80329 29504
rect 79943 29422 79990 29464
rect 80114 29422 80158 29464
rect 80282 29422 80329 29464
rect 95036 29462 95476 29536
rect 95036 29338 95110 29462
rect 95234 29338 95278 29462
rect 95402 29338 95476 29462
rect 95036 29294 95476 29338
rect 95036 29170 95110 29294
rect 95234 29170 95278 29294
rect 95402 29170 95476 29294
rect 95036 29096 95476 29170
rect 18196 29022 18636 29096
rect 18196 28898 18270 29022
rect 18394 28898 18438 29022
rect 18562 28898 18636 29022
rect 18196 28854 18636 28898
rect 3103 28748 3150 28790
rect 3274 28748 3318 28790
rect 3442 28748 3489 28790
rect 3103 28708 3112 28748
rect 3274 28708 3276 28748
rect 3316 28708 3318 28748
rect 3480 28708 3489 28748
rect 3103 28666 3150 28708
rect 3274 28666 3318 28708
rect 3442 28666 3489 28708
rect 18196 28730 18270 28854
rect 18394 28730 18438 28854
rect 18562 28730 18636 28854
rect 18196 28656 18636 28730
rect 33316 29022 33756 29096
rect 33316 28898 33390 29022
rect 33514 28898 33558 29022
rect 33682 28898 33756 29022
rect 33316 28854 33756 28898
rect 33316 28730 33390 28854
rect 33514 28730 33558 28854
rect 33682 28730 33756 28854
rect 33316 28656 33756 28730
rect 48436 29022 48876 29096
rect 48436 28898 48510 29022
rect 48634 28898 48678 29022
rect 48802 28898 48876 29022
rect 48436 28854 48876 28898
rect 48436 28730 48510 28854
rect 48634 28730 48678 28854
rect 48802 28730 48876 28854
rect 48436 28656 48876 28730
rect 63556 29022 63996 29096
rect 63556 28898 63630 29022
rect 63754 28898 63798 29022
rect 63922 28898 63996 29022
rect 63556 28854 63996 28898
rect 63556 28730 63630 28854
rect 63754 28730 63798 28854
rect 63922 28730 63996 28854
rect 63556 28656 63996 28730
rect 78703 28748 78750 28790
rect 78874 28748 78918 28790
rect 79042 28748 79089 28790
rect 78703 28708 78712 28748
rect 78874 28708 78876 28748
rect 78916 28708 78918 28748
rect 79080 28708 79089 28748
rect 78703 28666 78750 28708
rect 78874 28666 78918 28708
rect 79042 28666 79089 28708
rect 84931 28372 84940 28412
rect 84980 28372 97324 28412
rect 97364 28372 97373 28412
rect 93796 28222 94236 28296
rect 93796 28098 93870 28222
rect 93994 28098 94038 28222
rect 94162 28098 94236 28222
rect 93796 28054 94236 28098
rect 4343 27992 4390 28034
rect 4514 27992 4558 28034
rect 4682 27992 4729 28034
rect 4343 27952 4352 27992
rect 4514 27952 4516 27992
rect 4556 27952 4558 27992
rect 4720 27952 4729 27992
rect 4343 27910 4390 27952
rect 4514 27910 4558 27952
rect 4682 27910 4729 27952
rect 79943 27992 79990 28034
rect 80114 27992 80158 28034
rect 80282 27992 80329 28034
rect 79943 27952 79952 27992
rect 80114 27952 80116 27992
rect 80156 27952 80158 27992
rect 80320 27952 80329 27992
rect 79943 27910 79990 27952
rect 80114 27910 80158 27952
rect 80282 27910 80329 27952
rect 93796 27930 93870 28054
rect 93994 27930 94038 28054
rect 94162 27930 94236 28054
rect 93796 27856 94236 27930
rect 3103 27236 3150 27278
rect 3274 27236 3318 27278
rect 3442 27236 3489 27278
rect 3103 27196 3112 27236
rect 3274 27196 3276 27236
rect 3316 27196 3318 27236
rect 3480 27196 3489 27236
rect 3103 27154 3150 27196
rect 3274 27154 3318 27196
rect 3442 27154 3489 27196
rect 78703 27236 78750 27278
rect 78874 27236 78918 27278
rect 79042 27236 79089 27278
rect 78703 27196 78712 27236
rect 78874 27196 78876 27236
rect 78916 27196 78918 27236
rect 79080 27196 79089 27236
rect 78703 27154 78750 27196
rect 78874 27154 78918 27196
rect 79042 27154 79089 27196
rect 4343 26480 4390 26522
rect 4514 26480 4558 26522
rect 4682 26480 4729 26522
rect 4343 26440 4352 26480
rect 4514 26440 4516 26480
rect 4556 26440 4558 26480
rect 4720 26440 4729 26480
rect 4343 26398 4390 26440
rect 4514 26398 4558 26440
rect 4682 26398 4729 26440
rect 79943 26480 79990 26522
rect 80114 26480 80158 26522
rect 80282 26480 80329 26522
rect 79943 26440 79952 26480
rect 80114 26440 80116 26480
rect 80156 26440 80158 26480
rect 80320 26440 80329 26480
rect 79943 26398 79990 26440
rect 80114 26398 80158 26440
rect 80282 26398 80329 26440
rect 3103 25724 3150 25766
rect 3274 25724 3318 25766
rect 3442 25724 3489 25766
rect 3103 25684 3112 25724
rect 3274 25684 3276 25724
rect 3316 25684 3318 25724
rect 3480 25684 3489 25724
rect 3103 25642 3150 25684
rect 3274 25642 3318 25684
rect 3442 25642 3489 25684
rect 78703 25724 78750 25766
rect 78874 25724 78918 25766
rect 79042 25724 79089 25766
rect 78703 25684 78712 25724
rect 78874 25684 78876 25724
rect 78916 25684 78918 25724
rect 79080 25684 79089 25724
rect 78703 25642 78750 25684
rect 78874 25642 78918 25684
rect 79042 25642 79089 25684
rect 4343 24968 4390 25010
rect 4514 24968 4558 25010
rect 4682 24968 4729 25010
rect 4343 24928 4352 24968
rect 4514 24928 4516 24968
rect 4556 24928 4558 24968
rect 4720 24928 4729 24968
rect 4343 24886 4390 24928
rect 4514 24886 4558 24928
rect 4682 24886 4729 24928
rect 79943 24968 79990 25010
rect 80114 24968 80158 25010
rect 80282 24968 80329 25010
rect 79943 24928 79952 24968
rect 80114 24928 80116 24968
rect 80156 24928 80158 24968
rect 80320 24928 80329 24968
rect 79943 24886 79990 24928
rect 80114 24886 80158 24928
rect 80282 24886 80329 24928
rect 19436 24262 19876 24336
rect 3103 24212 3150 24254
rect 3274 24212 3318 24254
rect 3442 24212 3489 24254
rect 3103 24172 3112 24212
rect 3274 24172 3276 24212
rect 3316 24172 3318 24212
rect 3480 24172 3489 24212
rect 3103 24130 3150 24172
rect 3274 24130 3318 24172
rect 3442 24130 3489 24172
rect 19436 24138 19510 24262
rect 19634 24138 19678 24262
rect 19802 24138 19876 24262
rect 19436 24094 19876 24138
rect 19436 23970 19510 24094
rect 19634 23970 19678 24094
rect 19802 23970 19876 24094
rect 19436 23896 19876 23970
rect 34556 24262 34996 24336
rect 34556 24138 34630 24262
rect 34754 24138 34798 24262
rect 34922 24138 34996 24262
rect 34556 24094 34996 24138
rect 34556 23970 34630 24094
rect 34754 23970 34798 24094
rect 34922 23970 34996 24094
rect 34556 23896 34996 23970
rect 49676 24262 50116 24336
rect 49676 24138 49750 24262
rect 49874 24138 49918 24262
rect 50042 24138 50116 24262
rect 49676 24094 50116 24138
rect 49676 23970 49750 24094
rect 49874 23970 49918 24094
rect 50042 23970 50116 24094
rect 49676 23896 50116 23970
rect 64796 24262 65236 24336
rect 64796 24138 64870 24262
rect 64994 24138 65038 24262
rect 65162 24138 65236 24262
rect 64796 24094 65236 24138
rect 78703 24212 78750 24254
rect 78874 24212 78918 24254
rect 79042 24212 79089 24254
rect 78703 24172 78712 24212
rect 78874 24172 78876 24212
rect 78916 24172 78918 24212
rect 79080 24172 79089 24212
rect 78703 24130 78750 24172
rect 78874 24130 78918 24172
rect 79042 24130 79089 24172
rect 64796 23970 64870 24094
rect 64994 23970 65038 24094
rect 65162 23970 65236 24094
rect 64796 23896 65236 23970
rect 4343 23456 4390 23498
rect 4514 23456 4558 23498
rect 4682 23456 4729 23498
rect 4343 23416 4352 23456
rect 4514 23416 4516 23456
rect 4556 23416 4558 23456
rect 4720 23416 4729 23456
rect 4343 23374 4390 23416
rect 4514 23374 4558 23416
rect 4682 23374 4729 23416
rect 79943 23456 79990 23498
rect 80114 23456 80158 23498
rect 80282 23456 80329 23498
rect 79943 23416 79952 23456
rect 80114 23416 80116 23456
rect 80156 23416 80158 23456
rect 80320 23416 80329 23456
rect 79943 23374 79990 23416
rect 80114 23374 80158 23416
rect 80282 23374 80329 23416
rect 18196 23022 18636 23096
rect 18196 22898 18270 23022
rect 18394 22898 18438 23022
rect 18562 22898 18636 23022
rect 18196 22854 18636 22898
rect 3103 22700 3150 22742
rect 3274 22700 3318 22742
rect 3442 22700 3489 22742
rect 3103 22660 3112 22700
rect 3274 22660 3276 22700
rect 3316 22660 3318 22700
rect 3480 22660 3489 22700
rect 3103 22618 3150 22660
rect 3274 22618 3318 22660
rect 3442 22618 3489 22660
rect 18196 22730 18270 22854
rect 18394 22730 18438 22854
rect 18562 22730 18636 22854
rect 18196 22656 18636 22730
rect 33316 23022 33756 23096
rect 33316 22898 33390 23022
rect 33514 22898 33558 23022
rect 33682 22898 33756 23022
rect 33316 22854 33756 22898
rect 33316 22730 33390 22854
rect 33514 22730 33558 22854
rect 33682 22730 33756 22854
rect 33316 22656 33756 22730
rect 48436 23022 48876 23096
rect 48436 22898 48510 23022
rect 48634 22898 48678 23022
rect 48802 22898 48876 23022
rect 48436 22854 48876 22898
rect 48436 22730 48510 22854
rect 48634 22730 48678 22854
rect 48802 22730 48876 22854
rect 48436 22656 48876 22730
rect 63556 23022 63996 23096
rect 63556 22898 63630 23022
rect 63754 22898 63798 23022
rect 63922 22898 63996 23022
rect 63556 22854 63996 22898
rect 63556 22730 63630 22854
rect 63754 22730 63798 22854
rect 63922 22730 63996 22854
rect 63556 22656 63996 22730
rect 78703 22700 78750 22742
rect 78874 22700 78918 22742
rect 79042 22700 79089 22742
rect 78703 22660 78712 22700
rect 78874 22660 78876 22700
rect 78916 22660 78918 22700
rect 79080 22660 79089 22700
rect 78703 22618 78750 22660
rect 78874 22618 78918 22660
rect 79042 22618 79089 22660
rect 4343 21944 4390 21986
rect 4514 21944 4558 21986
rect 4682 21944 4729 21986
rect 4343 21904 4352 21944
rect 4514 21904 4516 21944
rect 4556 21904 4558 21944
rect 4720 21904 4729 21944
rect 4343 21862 4390 21904
rect 4514 21862 4558 21904
rect 4682 21862 4729 21904
rect 79943 21944 79990 21986
rect 80114 21944 80158 21986
rect 80282 21944 80329 21986
rect 79943 21904 79952 21944
rect 80114 21904 80116 21944
rect 80156 21904 80158 21944
rect 80320 21904 80329 21944
rect 79943 21862 79990 21904
rect 80114 21862 80158 21904
rect 80282 21862 80329 21904
rect 95063 21944 95110 21986
rect 95234 21944 95278 21986
rect 95402 21944 95449 21986
rect 95063 21904 95072 21944
rect 95234 21904 95236 21944
rect 95276 21904 95278 21944
rect 95440 21904 95449 21944
rect 95063 21862 95110 21904
rect 95234 21862 95278 21904
rect 95402 21862 95449 21904
rect 3103 21188 3150 21230
rect 3274 21188 3318 21230
rect 3442 21188 3489 21230
rect 3103 21148 3112 21188
rect 3274 21148 3276 21188
rect 3316 21148 3318 21188
rect 3480 21148 3489 21188
rect 3103 21106 3150 21148
rect 3274 21106 3318 21148
rect 3442 21106 3489 21148
rect 78703 21188 78750 21230
rect 78874 21188 78918 21230
rect 79042 21188 79089 21230
rect 78703 21148 78712 21188
rect 78874 21148 78876 21188
rect 78916 21148 78918 21188
rect 79080 21148 79089 21188
rect 78703 21106 78750 21148
rect 78874 21106 78918 21148
rect 79042 21106 79089 21148
rect 93823 21188 93870 21230
rect 93994 21188 94038 21230
rect 94162 21188 94209 21230
rect 93823 21148 93832 21188
rect 93994 21148 93996 21188
rect 94036 21148 94038 21188
rect 94200 21148 94209 21188
rect 93823 21106 93870 21148
rect 93994 21106 94038 21148
rect 94162 21106 94209 21148
rect 4343 20432 4390 20474
rect 4514 20432 4558 20474
rect 4682 20432 4729 20474
rect 4343 20392 4352 20432
rect 4514 20392 4516 20432
rect 4556 20392 4558 20432
rect 4720 20392 4729 20432
rect 4343 20350 4390 20392
rect 4514 20350 4558 20392
rect 4682 20350 4729 20392
rect 79943 20432 79990 20474
rect 80114 20432 80158 20474
rect 80282 20432 80329 20474
rect 79943 20392 79952 20432
rect 80114 20392 80116 20432
rect 80156 20392 80158 20432
rect 80320 20392 80329 20432
rect 79943 20350 79990 20392
rect 80114 20350 80158 20392
rect 80282 20350 80329 20392
rect 95063 20432 95110 20474
rect 95234 20432 95278 20474
rect 95402 20432 95449 20474
rect 95063 20392 95072 20432
rect 95234 20392 95236 20432
rect 95276 20392 95278 20432
rect 95440 20392 95449 20432
rect 95063 20350 95110 20392
rect 95234 20350 95278 20392
rect 95402 20350 95449 20392
rect 3103 19676 3150 19718
rect 3274 19676 3318 19718
rect 3442 19676 3489 19718
rect 3103 19636 3112 19676
rect 3274 19636 3276 19676
rect 3316 19636 3318 19676
rect 3480 19636 3489 19676
rect 3103 19594 3150 19636
rect 3274 19594 3318 19636
rect 3442 19594 3489 19636
rect 78703 19676 78750 19718
rect 78874 19676 78918 19718
rect 79042 19676 79089 19718
rect 78703 19636 78712 19676
rect 78874 19636 78876 19676
rect 78916 19636 78918 19676
rect 79080 19636 79089 19676
rect 78703 19594 78750 19636
rect 78874 19594 78918 19636
rect 79042 19594 79089 19636
rect 93823 19676 93870 19718
rect 93994 19676 94038 19718
rect 94162 19676 94209 19718
rect 93823 19636 93832 19676
rect 93994 19636 93996 19676
rect 94036 19636 94038 19676
rect 94200 19636 94209 19676
rect 93823 19594 93870 19636
rect 93994 19594 94038 19636
rect 94162 19594 94209 19636
rect 4343 18920 4390 18962
rect 4514 18920 4558 18962
rect 4682 18920 4729 18962
rect 4343 18880 4352 18920
rect 4514 18880 4516 18920
rect 4556 18880 4558 18920
rect 4720 18880 4729 18920
rect 4343 18838 4390 18880
rect 4514 18838 4558 18880
rect 4682 18838 4729 18880
rect 79943 18920 79990 18962
rect 80114 18920 80158 18962
rect 80282 18920 80329 18962
rect 79943 18880 79952 18920
rect 80114 18880 80116 18920
rect 80156 18880 80158 18920
rect 80320 18880 80329 18920
rect 79943 18838 79990 18880
rect 80114 18838 80158 18880
rect 80282 18838 80329 18880
rect 19436 18262 19876 18336
rect 3103 18164 3150 18206
rect 3274 18164 3318 18206
rect 3442 18164 3489 18206
rect 3103 18124 3112 18164
rect 3274 18124 3276 18164
rect 3316 18124 3318 18164
rect 3480 18124 3489 18164
rect 3103 18082 3150 18124
rect 3274 18082 3318 18124
rect 3442 18082 3489 18124
rect 19436 18138 19510 18262
rect 19634 18138 19678 18262
rect 19802 18138 19876 18262
rect 19436 18094 19876 18138
rect 19436 17970 19510 18094
rect 19634 17970 19678 18094
rect 19802 17970 19876 18094
rect 19436 17896 19876 17970
rect 34556 18262 34996 18336
rect 34556 18138 34630 18262
rect 34754 18138 34798 18262
rect 34922 18138 34996 18262
rect 34556 18094 34996 18138
rect 34556 17970 34630 18094
rect 34754 17970 34798 18094
rect 34922 17970 34996 18094
rect 34556 17896 34996 17970
rect 49676 18262 50116 18336
rect 49676 18138 49750 18262
rect 49874 18138 49918 18262
rect 50042 18138 50116 18262
rect 49676 18094 50116 18138
rect 49676 17970 49750 18094
rect 49874 17970 49918 18094
rect 50042 17970 50116 18094
rect 49676 17896 50116 17970
rect 64796 18262 65236 18336
rect 64796 18138 64870 18262
rect 64994 18138 65038 18262
rect 65162 18138 65236 18262
rect 64796 18094 65236 18138
rect 64796 17970 64870 18094
rect 64994 17970 65038 18094
rect 65162 17970 65236 18094
rect 78703 18164 78750 18206
rect 78874 18164 78918 18206
rect 79042 18164 79089 18206
rect 78703 18124 78712 18164
rect 78874 18124 78876 18164
rect 78916 18124 78918 18164
rect 79080 18124 79089 18164
rect 78703 18082 78750 18124
rect 78874 18082 78918 18124
rect 79042 18082 79089 18124
rect 64796 17896 65236 17970
rect 4343 17408 4390 17450
rect 4514 17408 4558 17450
rect 4682 17408 4729 17450
rect 4343 17368 4352 17408
rect 4514 17368 4516 17408
rect 4556 17368 4558 17408
rect 4720 17368 4729 17408
rect 4343 17326 4390 17368
rect 4514 17326 4558 17368
rect 4682 17326 4729 17368
rect 79943 17408 79990 17450
rect 80114 17408 80158 17450
rect 80282 17408 80329 17450
rect 79943 17368 79952 17408
rect 80114 17368 80116 17408
rect 80156 17368 80158 17408
rect 80320 17368 80329 17408
rect 79943 17326 79990 17368
rect 80114 17326 80158 17368
rect 80282 17326 80329 17368
rect 18196 17022 18636 17096
rect 18196 16898 18270 17022
rect 18394 16898 18438 17022
rect 18562 16898 18636 17022
rect 18196 16854 18636 16898
rect 18196 16730 18270 16854
rect 18394 16730 18438 16854
rect 18562 16730 18636 16854
rect 3103 16652 3150 16694
rect 3274 16652 3318 16694
rect 3442 16652 3489 16694
rect 18196 16656 18636 16730
rect 33316 17022 33756 17096
rect 33316 16898 33390 17022
rect 33514 16898 33558 17022
rect 33682 16898 33756 17022
rect 33316 16854 33756 16898
rect 33316 16730 33390 16854
rect 33514 16730 33558 16854
rect 33682 16730 33756 16854
rect 33316 16656 33756 16730
rect 48436 17022 48876 17096
rect 48436 16898 48510 17022
rect 48634 16898 48678 17022
rect 48802 16898 48876 17022
rect 48436 16854 48876 16898
rect 48436 16730 48510 16854
rect 48634 16730 48678 16854
rect 48802 16730 48876 16854
rect 48436 16656 48876 16730
rect 63556 17022 63996 17096
rect 63556 16898 63630 17022
rect 63754 16898 63798 17022
rect 63922 16898 63996 17022
rect 63556 16854 63996 16898
rect 63556 16730 63630 16854
rect 63754 16730 63798 16854
rect 63922 16730 63996 16854
rect 63556 16656 63996 16730
rect 3103 16612 3112 16652
rect 3274 16612 3276 16652
rect 3316 16612 3318 16652
rect 3480 16612 3489 16652
rect 3103 16570 3150 16612
rect 3274 16570 3318 16612
rect 3442 16570 3489 16612
rect 78703 16652 78750 16694
rect 78874 16652 78918 16694
rect 79042 16652 79089 16694
rect 78703 16612 78712 16652
rect 78874 16612 78876 16652
rect 78916 16612 78918 16652
rect 79080 16612 79089 16652
rect 78703 16570 78750 16612
rect 78874 16570 78918 16612
rect 79042 16570 79089 16612
rect 4343 15896 4390 15938
rect 4514 15896 4558 15938
rect 4682 15896 4729 15938
rect 4343 15856 4352 15896
rect 4514 15856 4516 15896
rect 4556 15856 4558 15896
rect 4720 15856 4729 15896
rect 4343 15814 4390 15856
rect 4514 15814 4558 15856
rect 4682 15814 4729 15856
rect 79943 15896 79990 15938
rect 80114 15896 80158 15938
rect 80282 15896 80329 15938
rect 79943 15856 79952 15896
rect 80114 15856 80116 15896
rect 80156 15856 80158 15896
rect 80320 15856 80329 15896
rect 79943 15814 79990 15856
rect 80114 15814 80158 15856
rect 80282 15814 80329 15856
rect 3103 15140 3150 15182
rect 3274 15140 3318 15182
rect 3442 15140 3489 15182
rect 3103 15100 3112 15140
rect 3274 15100 3276 15140
rect 3316 15100 3318 15140
rect 3480 15100 3489 15140
rect 3103 15058 3150 15100
rect 3274 15058 3318 15100
rect 3442 15058 3489 15100
rect 78703 15140 78750 15182
rect 78874 15140 78918 15182
rect 79042 15140 79089 15182
rect 78703 15100 78712 15140
rect 78874 15100 78876 15140
rect 78916 15100 78918 15140
rect 79080 15100 79089 15140
rect 78703 15058 78750 15100
rect 78874 15058 78918 15100
rect 79042 15058 79089 15100
rect 4343 14384 4390 14426
rect 4514 14384 4558 14426
rect 4682 14384 4729 14426
rect 4343 14344 4352 14384
rect 4514 14344 4516 14384
rect 4556 14344 4558 14384
rect 4720 14344 4729 14384
rect 4343 14302 4390 14344
rect 4514 14302 4558 14344
rect 4682 14302 4729 14344
rect 79943 14384 79990 14426
rect 80114 14384 80158 14426
rect 80282 14384 80329 14426
rect 79943 14344 79952 14384
rect 80114 14344 80116 14384
rect 80156 14344 80158 14384
rect 80320 14344 80329 14384
rect 79943 14302 79990 14344
rect 80114 14302 80158 14344
rect 80282 14302 80329 14344
rect 3103 13628 3150 13670
rect 3274 13628 3318 13670
rect 3442 13628 3489 13670
rect 3103 13588 3112 13628
rect 3274 13588 3276 13628
rect 3316 13588 3318 13628
rect 3480 13588 3489 13628
rect 3103 13546 3150 13588
rect 3274 13546 3318 13588
rect 3442 13546 3489 13588
rect 78703 13628 78750 13670
rect 78874 13628 78918 13670
rect 79042 13628 79089 13670
rect 78703 13588 78712 13628
rect 78874 13588 78876 13628
rect 78916 13588 78918 13628
rect 79080 13588 79089 13628
rect 78703 13546 78750 13588
rect 78874 13546 78918 13588
rect 79042 13546 79089 13588
rect 4343 12872 4390 12914
rect 4514 12872 4558 12914
rect 4682 12872 4729 12914
rect 4343 12832 4352 12872
rect 4514 12832 4516 12872
rect 4556 12832 4558 12872
rect 4720 12832 4729 12872
rect 4343 12790 4390 12832
rect 4514 12790 4558 12832
rect 4682 12790 4729 12832
rect 79943 12872 79990 12914
rect 80114 12872 80158 12914
rect 80282 12872 80329 12914
rect 79943 12832 79952 12872
rect 80114 12832 80116 12872
rect 80156 12832 80158 12872
rect 80320 12832 80329 12872
rect 79943 12790 79990 12832
rect 80114 12790 80158 12832
rect 80282 12790 80329 12832
rect 19436 12262 19876 12336
rect 3103 12116 3150 12158
rect 3274 12116 3318 12158
rect 3442 12116 3489 12158
rect 3103 12076 3112 12116
rect 3274 12076 3276 12116
rect 3316 12076 3318 12116
rect 3480 12076 3489 12116
rect 3103 12034 3150 12076
rect 3274 12034 3318 12076
rect 3442 12034 3489 12076
rect 19436 12138 19510 12262
rect 19634 12138 19678 12262
rect 19802 12138 19876 12262
rect 19436 12094 19876 12138
rect 19436 11970 19510 12094
rect 19634 11970 19678 12094
rect 19802 11970 19876 12094
rect 19436 11896 19876 11970
rect 34556 12262 34996 12336
rect 34556 12138 34630 12262
rect 34754 12138 34798 12262
rect 34922 12138 34996 12262
rect 34556 12094 34996 12138
rect 34556 11970 34630 12094
rect 34754 11970 34798 12094
rect 34922 11970 34996 12094
rect 34556 11896 34996 11970
rect 49676 12262 50116 12336
rect 49676 12138 49750 12262
rect 49874 12138 49918 12262
rect 50042 12138 50116 12262
rect 49676 12094 50116 12138
rect 49676 11970 49750 12094
rect 49874 11970 49918 12094
rect 50042 11970 50116 12094
rect 49676 11896 50116 11970
rect 64796 12262 65236 12336
rect 64796 12138 64870 12262
rect 64994 12138 65038 12262
rect 65162 12138 65236 12262
rect 95036 12262 95476 12336
rect 64796 12094 65236 12138
rect 64796 11970 64870 12094
rect 64994 11970 65038 12094
rect 65162 11970 65236 12094
rect 78703 12116 78750 12158
rect 78874 12116 78918 12158
rect 79042 12116 79089 12158
rect 78703 12076 78712 12116
rect 78874 12076 78876 12116
rect 78916 12076 78918 12116
rect 79080 12076 79089 12116
rect 78703 12034 78750 12076
rect 78874 12034 78918 12076
rect 79042 12034 79089 12076
rect 95036 12138 95110 12262
rect 95234 12138 95278 12262
rect 95402 12138 95476 12262
rect 95036 12094 95476 12138
rect 64796 11896 65236 11970
rect 95036 11970 95110 12094
rect 95234 11970 95278 12094
rect 95402 11970 95476 12094
rect 95036 11896 95476 11970
rect 4343 11360 4390 11402
rect 4514 11360 4558 11402
rect 4682 11360 4729 11402
rect 4343 11320 4352 11360
rect 4514 11320 4516 11360
rect 4556 11320 4558 11360
rect 4720 11320 4729 11360
rect 4343 11278 4390 11320
rect 4514 11278 4558 11320
rect 4682 11278 4729 11320
rect 79943 11360 79990 11402
rect 80114 11360 80158 11402
rect 80282 11360 80329 11402
rect 79943 11320 79952 11360
rect 80114 11320 80116 11360
rect 80156 11320 80158 11360
rect 80320 11320 80329 11360
rect 79943 11278 79990 11320
rect 80114 11278 80158 11320
rect 80282 11278 80329 11320
rect 18196 11022 18636 11096
rect 18196 10898 18270 11022
rect 18394 10898 18438 11022
rect 18562 10898 18636 11022
rect 18196 10854 18636 10898
rect 18196 10730 18270 10854
rect 18394 10730 18438 10854
rect 18562 10730 18636 10854
rect 18196 10656 18636 10730
rect 33316 11022 33756 11096
rect 33316 10898 33390 11022
rect 33514 10898 33558 11022
rect 33682 10898 33756 11022
rect 33316 10854 33756 10898
rect 33316 10730 33390 10854
rect 33514 10730 33558 10854
rect 33682 10730 33756 10854
rect 33316 10656 33756 10730
rect 48436 11022 48876 11096
rect 48436 10898 48510 11022
rect 48634 10898 48678 11022
rect 48802 10898 48876 11022
rect 48436 10854 48876 10898
rect 48436 10730 48510 10854
rect 48634 10730 48678 10854
rect 48802 10730 48876 10854
rect 48436 10656 48876 10730
rect 63556 11022 63996 11096
rect 63556 10898 63630 11022
rect 63754 10898 63798 11022
rect 63922 10898 63996 11022
rect 63556 10854 63996 10898
rect 63556 10730 63630 10854
rect 63754 10730 63798 10854
rect 63922 10730 63996 10854
rect 63556 10656 63996 10730
rect 93796 11022 94236 11096
rect 93796 10898 93870 11022
rect 93994 10898 94038 11022
rect 94162 10898 94236 11022
rect 93796 10854 94236 10898
rect 93796 10730 93870 10854
rect 93994 10730 94038 10854
rect 94162 10730 94236 10854
rect 93796 10656 94236 10730
rect 3103 10604 3150 10646
rect 3274 10604 3318 10646
rect 3442 10604 3489 10646
rect 3103 10564 3112 10604
rect 3274 10564 3276 10604
rect 3316 10564 3318 10604
rect 3480 10564 3489 10604
rect 3103 10522 3150 10564
rect 3274 10522 3318 10564
rect 3442 10522 3489 10564
rect 78703 10604 78750 10646
rect 78874 10604 78918 10646
rect 79042 10604 79089 10646
rect 78703 10564 78712 10604
rect 78874 10564 78876 10604
rect 78916 10564 78918 10604
rect 79080 10564 79089 10604
rect 78703 10522 78750 10564
rect 78874 10522 78918 10564
rect 79042 10522 79089 10564
rect 4343 9848 4390 9890
rect 4514 9848 4558 9890
rect 4682 9848 4729 9890
rect 4343 9808 4352 9848
rect 4514 9808 4516 9848
rect 4556 9808 4558 9848
rect 4720 9808 4729 9848
rect 4343 9766 4390 9808
rect 4514 9766 4558 9808
rect 4682 9766 4729 9808
rect 79943 9848 79990 9890
rect 80114 9848 80158 9890
rect 80282 9848 80329 9890
rect 79943 9808 79952 9848
rect 80114 9808 80116 9848
rect 80156 9808 80158 9848
rect 80320 9808 80329 9848
rect 79943 9766 79990 9808
rect 80114 9766 80158 9808
rect 80282 9766 80329 9808
rect 73315 9220 73324 9260
rect 73364 9220 98740 9260
rect 98780 9220 98789 9260
rect 3103 9092 3150 9134
rect 3274 9092 3318 9134
rect 3442 9092 3489 9134
rect 3103 9052 3112 9092
rect 3274 9052 3276 9092
rect 3316 9052 3318 9092
rect 3480 9052 3489 9092
rect 3103 9010 3150 9052
rect 3274 9010 3318 9052
rect 3442 9010 3489 9052
rect 78703 9092 78750 9134
rect 78874 9092 78918 9134
rect 79042 9092 79089 9134
rect 78703 9052 78712 9092
rect 78874 9052 78876 9092
rect 78916 9052 78918 9092
rect 79080 9052 79089 9092
rect 78703 9010 78750 9052
rect 78874 9010 78918 9052
rect 79042 9010 79089 9052
rect 75523 8884 75532 8924
rect 75572 8884 98740 8924
rect 98780 8884 98789 8924
rect 4343 8336 4390 8378
rect 4514 8336 4558 8378
rect 4682 8336 4729 8378
rect 4343 8296 4352 8336
rect 4514 8296 4516 8336
rect 4556 8296 4558 8336
rect 4720 8296 4729 8336
rect 4343 8254 4390 8296
rect 4514 8254 4558 8296
rect 4682 8254 4729 8296
rect 79943 8336 79990 8378
rect 80114 8336 80158 8378
rect 80282 8336 80329 8378
rect 79943 8296 79952 8336
rect 80114 8296 80116 8336
rect 80156 8296 80158 8336
rect 80320 8296 80329 8336
rect 79943 8254 79990 8296
rect 80114 8254 80158 8296
rect 80282 8254 80329 8296
rect 71491 7876 71500 7916
rect 71540 7876 98860 7916
rect 98900 7876 98909 7916
rect 3523 7792 3532 7832
rect 3572 7792 38860 7832
rect 38900 7792 40876 7832
rect 40916 7792 40925 7832
rect 3103 7580 3150 7622
rect 3274 7580 3318 7622
rect 3442 7580 3489 7622
rect 3103 7540 3112 7580
rect 3274 7540 3276 7580
rect 3316 7540 3318 7580
rect 3480 7540 3489 7580
rect 3103 7498 3150 7540
rect 3274 7498 3318 7540
rect 3442 7498 3489 7540
rect 78703 7580 78750 7622
rect 78874 7580 78918 7622
rect 79042 7580 79089 7622
rect 78703 7540 78712 7580
rect 78874 7540 78876 7580
rect 78916 7540 78918 7580
rect 79080 7540 79089 7580
rect 78703 7498 78750 7540
rect 78874 7498 78918 7540
rect 79042 7498 79089 7540
rect 4343 6824 4390 6866
rect 4514 6824 4558 6866
rect 4682 6824 4729 6866
rect 4343 6784 4352 6824
rect 4514 6784 4516 6824
rect 4556 6784 4558 6824
rect 4720 6784 4729 6824
rect 4343 6742 4390 6784
rect 4514 6742 4558 6784
rect 4682 6742 4729 6784
rect 79943 6824 79990 6866
rect 80114 6824 80158 6866
rect 80282 6824 80329 6866
rect 79943 6784 79952 6824
rect 80114 6784 80116 6824
rect 80156 6784 80158 6824
rect 80320 6784 80329 6824
rect 79943 6742 79990 6784
rect 80114 6742 80158 6784
rect 80282 6742 80329 6784
rect 82051 6616 82060 6656
rect 82100 6616 98956 6656
rect 98996 6616 99005 6656
rect 95036 6262 95476 6336
rect 95036 6138 95110 6262
rect 95234 6138 95278 6262
rect 95402 6138 95476 6262
rect 3103 6068 3150 6110
rect 3274 6068 3318 6110
rect 3442 6068 3489 6110
rect 3103 6028 3112 6068
rect 3274 6028 3276 6068
rect 3316 6028 3318 6068
rect 3480 6028 3489 6068
rect 3103 5986 3150 6028
rect 3274 5986 3318 6028
rect 3442 5986 3489 6028
rect 78703 6068 78750 6110
rect 78874 6068 78918 6110
rect 79042 6068 79089 6110
rect 78703 6028 78712 6068
rect 78874 6028 78876 6068
rect 78916 6028 78918 6068
rect 79080 6028 79089 6068
rect 78703 5986 78750 6028
rect 78874 5986 78918 6028
rect 79042 5986 79089 6028
rect 95036 6094 95476 6138
rect 95036 5970 95110 6094
rect 95234 5970 95278 6094
rect 95402 5970 95476 6094
rect 95036 5896 95476 5970
rect 54595 5692 54604 5732
rect 54644 5692 67298 5732
rect 4343 5312 4390 5354
rect 4514 5312 4558 5354
rect 4682 5312 4729 5354
rect 4343 5272 4352 5312
rect 4514 5272 4516 5312
rect 4556 5272 4558 5312
rect 4720 5272 4729 5312
rect 4343 5230 4390 5272
rect 4514 5230 4558 5272
rect 4682 5230 4729 5272
rect 19463 5312 19510 5354
rect 19634 5312 19678 5354
rect 19802 5312 19849 5354
rect 19463 5272 19472 5312
rect 19634 5272 19636 5312
rect 19676 5272 19678 5312
rect 19840 5272 19849 5312
rect 19463 5230 19510 5272
rect 19634 5230 19678 5272
rect 19802 5230 19849 5272
rect 34583 5312 34630 5354
rect 34754 5312 34798 5354
rect 34922 5312 34969 5354
rect 34583 5272 34592 5312
rect 34754 5272 34756 5312
rect 34796 5272 34798 5312
rect 34960 5272 34969 5312
rect 34583 5230 34630 5272
rect 34754 5230 34798 5272
rect 34922 5230 34969 5272
rect 49703 5312 49750 5354
rect 49874 5312 49918 5354
rect 50042 5312 50089 5354
rect 49703 5272 49712 5312
rect 49874 5272 49876 5312
rect 49916 5272 49918 5312
rect 50080 5272 50089 5312
rect 49703 5230 49750 5272
rect 49874 5230 49918 5272
rect 50042 5230 50089 5272
rect 64823 5312 64870 5354
rect 64994 5312 65038 5354
rect 65162 5312 65209 5354
rect 64823 5272 64832 5312
rect 64994 5272 64996 5312
rect 65036 5272 65038 5312
rect 65200 5272 65209 5312
rect 64823 5230 64870 5272
rect 64994 5230 65038 5272
rect 65162 5230 65209 5272
rect 79943 5312 79990 5354
rect 80114 5312 80158 5354
rect 80282 5312 80329 5354
rect 79943 5272 79952 5312
rect 80114 5272 80116 5312
rect 80156 5272 80158 5312
rect 80320 5272 80329 5312
rect 79943 5230 79990 5272
rect 80114 5230 80158 5272
rect 80282 5230 80329 5272
rect 93796 5022 94236 5096
rect 93796 4898 93870 5022
rect 93994 4898 94038 5022
rect 94162 4898 94236 5022
rect 93796 4854 94236 4898
rect 59779 4684 59788 4724
rect 59828 4684 66386 4724
rect 93796 4730 93870 4854
rect 93994 4730 94038 4854
rect 94162 4730 94236 4854
rect 93796 4656 94236 4730
rect 3103 4556 3150 4598
rect 3274 4556 3318 4598
rect 3442 4556 3489 4598
rect 3103 4516 3112 4556
rect 3274 4516 3276 4556
rect 3316 4516 3318 4556
rect 3480 4516 3489 4556
rect 3103 4474 3150 4516
rect 3274 4474 3318 4516
rect 3442 4474 3489 4516
rect 18223 4556 18270 4598
rect 18394 4556 18438 4598
rect 18562 4556 18609 4598
rect 18223 4516 18232 4556
rect 18394 4516 18396 4556
rect 18436 4516 18438 4556
rect 18600 4516 18609 4556
rect 18223 4474 18270 4516
rect 18394 4474 18438 4516
rect 18562 4474 18609 4516
rect 33343 4556 33390 4598
rect 33514 4556 33558 4598
rect 33682 4556 33729 4598
rect 33343 4516 33352 4556
rect 33514 4516 33516 4556
rect 33556 4516 33558 4556
rect 33720 4516 33729 4556
rect 33343 4474 33390 4516
rect 33514 4474 33558 4516
rect 33682 4474 33729 4516
rect 48463 4556 48510 4598
rect 48634 4556 48678 4598
rect 48802 4556 48849 4598
rect 48463 4516 48472 4556
rect 48634 4516 48636 4556
rect 48676 4516 48678 4556
rect 48840 4516 48849 4556
rect 48463 4474 48510 4516
rect 48634 4474 48678 4516
rect 48802 4474 48849 4516
rect 63583 4556 63630 4598
rect 63754 4556 63798 4598
rect 63922 4556 63969 4598
rect 63583 4516 63592 4556
rect 63754 4516 63756 4556
rect 63796 4516 63798 4556
rect 63960 4516 63969 4556
rect 63583 4474 63630 4516
rect 63754 4474 63798 4516
rect 63922 4474 63969 4516
rect 78703 4556 78750 4598
rect 78874 4556 78918 4598
rect 79042 4556 79089 4598
rect 78703 4516 78712 4556
rect 78874 4516 78876 4556
rect 78916 4516 78918 4556
rect 79080 4516 79089 4556
rect 78703 4474 78750 4516
rect 78874 4474 78918 4516
rect 79042 4474 79089 4516
rect 43363 4096 43372 4136
rect 43412 4096 72652 4136
rect 72692 4096 72701 4136
rect 643 3928 652 3968
rect 692 3928 44524 3968
rect 44564 3928 44573 3968
rect 4343 3800 4390 3842
rect 4514 3800 4558 3842
rect 4682 3800 4729 3842
rect 4343 3760 4352 3800
rect 4514 3760 4516 3800
rect 4556 3760 4558 3800
rect 4720 3760 4729 3800
rect 4343 3718 4390 3760
rect 4514 3718 4558 3760
rect 4682 3718 4729 3760
rect 19463 3800 19510 3842
rect 19634 3800 19678 3842
rect 19802 3800 19849 3842
rect 19463 3760 19472 3800
rect 19634 3760 19636 3800
rect 19676 3760 19678 3800
rect 19840 3760 19849 3800
rect 19463 3718 19510 3760
rect 19634 3718 19678 3760
rect 19802 3718 19849 3760
rect 34583 3800 34630 3842
rect 34754 3800 34798 3842
rect 34922 3800 34969 3842
rect 34583 3760 34592 3800
rect 34754 3760 34756 3800
rect 34796 3760 34798 3800
rect 34960 3760 34969 3800
rect 34583 3718 34630 3760
rect 34754 3718 34798 3760
rect 34922 3718 34969 3760
rect 49703 3800 49750 3842
rect 49874 3800 49918 3842
rect 50042 3800 50089 3842
rect 49703 3760 49712 3800
rect 49874 3760 49876 3800
rect 49916 3760 49918 3800
rect 50080 3760 50089 3800
rect 49703 3718 49750 3760
rect 49874 3718 49918 3760
rect 50042 3718 50089 3760
rect 64823 3800 64870 3842
rect 64994 3800 65038 3842
rect 65162 3800 65209 3842
rect 64823 3760 64832 3800
rect 64994 3760 64996 3800
rect 65036 3760 65038 3800
rect 65200 3760 65209 3800
rect 64823 3718 64870 3760
rect 64994 3718 65038 3760
rect 65162 3718 65209 3760
rect 79943 3800 79990 3842
rect 80114 3800 80158 3842
rect 80282 3800 80329 3842
rect 79943 3760 79952 3800
rect 80114 3760 80116 3800
rect 80156 3760 80158 3800
rect 80320 3760 80329 3800
rect 79943 3718 79990 3760
rect 80114 3718 80158 3760
rect 80282 3718 80329 3760
rect 3103 3044 3150 3086
rect 3274 3044 3318 3086
rect 3442 3044 3489 3086
rect 3103 3004 3112 3044
rect 3274 3004 3276 3044
rect 3316 3004 3318 3044
rect 3480 3004 3489 3044
rect 3103 2962 3150 3004
rect 3274 2962 3318 3004
rect 3442 2962 3489 3004
rect 18223 3044 18270 3086
rect 18394 3044 18438 3086
rect 18562 3044 18609 3086
rect 18223 3004 18232 3044
rect 18394 3004 18396 3044
rect 18436 3004 18438 3044
rect 18600 3004 18609 3044
rect 18223 2962 18270 3004
rect 18394 2962 18438 3004
rect 18562 2962 18609 3004
rect 33343 3044 33390 3086
rect 33514 3044 33558 3086
rect 33682 3044 33729 3086
rect 33343 3004 33352 3044
rect 33514 3004 33516 3044
rect 33556 3004 33558 3044
rect 33720 3004 33729 3044
rect 33343 2962 33390 3004
rect 33514 2962 33558 3004
rect 33682 2962 33729 3004
rect 48463 3044 48510 3086
rect 48634 3044 48678 3086
rect 48802 3044 48849 3086
rect 48463 3004 48472 3044
rect 48634 3004 48636 3044
rect 48676 3004 48678 3044
rect 48840 3004 48849 3044
rect 48463 2962 48510 3004
rect 48634 2962 48678 3004
rect 48802 2962 48849 3004
rect 63583 3044 63630 3086
rect 63754 3044 63798 3086
rect 63922 3044 63969 3086
rect 63583 3004 63592 3044
rect 63754 3004 63756 3044
rect 63796 3004 63798 3044
rect 63960 3004 63969 3044
rect 63583 2962 63630 3004
rect 63754 2962 63798 3004
rect 63922 2962 63969 3004
rect 78703 3044 78750 3086
rect 78874 3044 78918 3086
rect 79042 3044 79089 3086
rect 78703 3004 78712 3044
rect 78874 3004 78876 3044
rect 78916 3004 78918 3044
rect 79080 3004 79089 3044
rect 78703 2962 78750 3004
rect 78874 2962 78918 3004
rect 79042 2962 79089 3004
rect 4343 2288 4390 2330
rect 4514 2288 4558 2330
rect 4682 2288 4729 2330
rect 4343 2248 4352 2288
rect 4514 2248 4516 2288
rect 4556 2248 4558 2288
rect 4720 2248 4729 2288
rect 4343 2206 4390 2248
rect 4514 2206 4558 2248
rect 4682 2206 4729 2248
rect 19463 2288 19510 2330
rect 19634 2288 19678 2330
rect 19802 2288 19849 2330
rect 19463 2248 19472 2288
rect 19634 2248 19636 2288
rect 19676 2248 19678 2288
rect 19840 2248 19849 2288
rect 19463 2206 19510 2248
rect 19634 2206 19678 2248
rect 19802 2206 19849 2248
rect 34583 2288 34630 2330
rect 34754 2288 34798 2330
rect 34922 2288 34969 2330
rect 34583 2248 34592 2288
rect 34754 2248 34756 2288
rect 34796 2248 34798 2288
rect 34960 2248 34969 2288
rect 34583 2206 34630 2248
rect 34754 2206 34798 2248
rect 34922 2206 34969 2248
rect 49703 2288 49750 2330
rect 49874 2288 49918 2330
rect 50042 2288 50089 2330
rect 49703 2248 49712 2288
rect 49874 2248 49876 2288
rect 49916 2248 49918 2288
rect 50080 2248 50089 2288
rect 49703 2206 49750 2248
rect 49874 2206 49918 2248
rect 50042 2206 50089 2248
rect 64823 2288 64870 2330
rect 64994 2288 65038 2330
rect 65162 2288 65209 2330
rect 64823 2248 64832 2288
rect 64994 2248 64996 2288
rect 65036 2248 65038 2288
rect 65200 2248 65209 2288
rect 64823 2206 64870 2248
rect 64994 2206 65038 2248
rect 65162 2206 65209 2248
rect 79943 2288 79990 2330
rect 80114 2288 80158 2330
rect 80282 2288 80329 2330
rect 79943 2248 79952 2288
rect 80114 2248 80116 2288
rect 80156 2248 80158 2288
rect 80320 2248 80329 2288
rect 79943 2206 79990 2248
rect 80114 2206 80158 2248
rect 80282 2206 80329 2248
rect 3103 1532 3150 1574
rect 3274 1532 3318 1574
rect 3442 1532 3489 1574
rect 3103 1492 3112 1532
rect 3274 1492 3276 1532
rect 3316 1492 3318 1532
rect 3480 1492 3489 1532
rect 3103 1450 3150 1492
rect 3274 1450 3318 1492
rect 3442 1450 3489 1492
rect 18223 1532 18270 1574
rect 18394 1532 18438 1574
rect 18562 1532 18609 1574
rect 18223 1492 18232 1532
rect 18394 1492 18396 1532
rect 18436 1492 18438 1532
rect 18600 1492 18609 1532
rect 18223 1450 18270 1492
rect 18394 1450 18438 1492
rect 18562 1450 18609 1492
rect 33343 1532 33390 1574
rect 33514 1532 33558 1574
rect 33682 1532 33729 1574
rect 33343 1492 33352 1532
rect 33514 1492 33516 1532
rect 33556 1492 33558 1532
rect 33720 1492 33729 1532
rect 33343 1450 33390 1492
rect 33514 1450 33558 1492
rect 33682 1450 33729 1492
rect 48463 1532 48510 1574
rect 48634 1532 48678 1574
rect 48802 1532 48849 1574
rect 48463 1492 48472 1532
rect 48634 1492 48636 1532
rect 48676 1492 48678 1532
rect 48840 1492 48849 1532
rect 48463 1450 48510 1492
rect 48634 1450 48678 1492
rect 48802 1450 48849 1492
rect 63583 1532 63630 1574
rect 63754 1532 63798 1574
rect 63922 1532 63969 1574
rect 63583 1492 63592 1532
rect 63754 1492 63756 1532
rect 63796 1492 63798 1532
rect 63960 1492 63969 1532
rect 63583 1450 63630 1492
rect 63754 1450 63798 1492
rect 63922 1450 63969 1492
rect 78703 1532 78750 1574
rect 78874 1532 78918 1574
rect 79042 1532 79089 1574
rect 78703 1492 78712 1532
rect 78874 1492 78876 1532
rect 78916 1492 78918 1532
rect 79080 1492 79089 1532
rect 78703 1450 78750 1492
rect 78874 1450 78918 1492
rect 79042 1450 79089 1492
rect 4343 776 4390 818
rect 4514 776 4558 818
rect 4682 776 4729 818
rect 4343 736 4352 776
rect 4514 736 4516 776
rect 4556 736 4558 776
rect 4720 736 4729 776
rect 4343 694 4390 736
rect 4514 694 4558 736
rect 4682 694 4729 736
rect 19463 776 19510 818
rect 19634 776 19678 818
rect 19802 776 19849 818
rect 19463 736 19472 776
rect 19634 736 19636 776
rect 19676 736 19678 776
rect 19840 736 19849 776
rect 19463 694 19510 736
rect 19634 694 19678 736
rect 19802 694 19849 736
rect 34583 776 34630 818
rect 34754 776 34798 818
rect 34922 776 34969 818
rect 34583 736 34592 776
rect 34754 736 34756 776
rect 34796 736 34798 776
rect 34960 736 34969 776
rect 34583 694 34630 736
rect 34754 694 34798 736
rect 34922 694 34969 736
rect 49703 776 49750 818
rect 49874 776 49918 818
rect 50042 776 50089 818
rect 49703 736 49712 776
rect 49874 736 49876 776
rect 49916 736 49918 776
rect 50080 736 50089 776
rect 49703 694 49750 736
rect 49874 694 49918 736
rect 50042 694 50089 736
rect 64823 776 64870 818
rect 64994 776 65038 818
rect 65162 776 65209 818
rect 64823 736 64832 776
rect 64994 736 64996 776
rect 65036 736 65038 776
rect 65200 736 65209 776
rect 64823 694 64870 736
rect 64994 694 65038 736
rect 65162 694 65209 736
rect 79943 776 79990 818
rect 80114 776 80158 818
rect 80282 776 80329 818
rect 79943 736 79952 776
rect 80114 736 80116 776
rect 80156 736 80158 776
rect 80320 736 80329 776
rect 79943 694 79990 736
rect 80114 694 80158 736
rect 80282 694 80329 736
<< via5 >>
rect 4390 38576 4514 38618
rect 4558 38576 4682 38618
rect 4390 38536 4392 38576
rect 4392 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4514 38576
rect 4558 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4680 38576
rect 4680 38536 4682 38576
rect 4390 38494 4514 38536
rect 4558 38494 4682 38536
rect 19510 38576 19634 38618
rect 19678 38576 19802 38618
rect 19510 38536 19512 38576
rect 19512 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19634 38576
rect 19678 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19800 38576
rect 19800 38536 19802 38576
rect 19510 38494 19634 38536
rect 19678 38494 19802 38536
rect 34630 38576 34754 38618
rect 34798 38576 34922 38618
rect 34630 38536 34632 38576
rect 34632 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34754 38576
rect 34798 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34920 38576
rect 34920 38536 34922 38576
rect 34630 38494 34754 38536
rect 34798 38494 34922 38536
rect 49750 38576 49874 38618
rect 49918 38576 50042 38618
rect 49750 38536 49752 38576
rect 49752 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49874 38576
rect 49918 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50040 38576
rect 50040 38536 50042 38576
rect 49750 38494 49874 38536
rect 49918 38494 50042 38536
rect 64870 38576 64994 38618
rect 65038 38576 65162 38618
rect 64870 38536 64872 38576
rect 64872 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64994 38576
rect 65038 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65160 38576
rect 65160 38536 65162 38576
rect 64870 38494 64994 38536
rect 65038 38494 65162 38536
rect 79990 38576 80114 38618
rect 80158 38576 80282 38618
rect 79990 38536 79992 38576
rect 79992 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80114 38576
rect 80158 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80280 38576
rect 80280 38536 80282 38576
rect 79990 38494 80114 38536
rect 80158 38494 80282 38536
rect 3150 37820 3274 37862
rect 3318 37820 3442 37862
rect 3150 37780 3152 37820
rect 3152 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3274 37820
rect 3318 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3440 37820
rect 3440 37780 3442 37820
rect 3150 37738 3274 37780
rect 3318 37738 3442 37780
rect 18270 37820 18394 37862
rect 18438 37820 18562 37862
rect 18270 37780 18272 37820
rect 18272 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18394 37820
rect 18438 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18560 37820
rect 18560 37780 18562 37820
rect 18270 37738 18394 37780
rect 18438 37738 18562 37780
rect 33390 37820 33514 37862
rect 33558 37820 33682 37862
rect 33390 37780 33392 37820
rect 33392 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33514 37820
rect 33558 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33680 37820
rect 33680 37780 33682 37820
rect 33390 37738 33514 37780
rect 33558 37738 33682 37780
rect 48510 37820 48634 37862
rect 48678 37820 48802 37862
rect 48510 37780 48512 37820
rect 48512 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48634 37820
rect 48678 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48800 37820
rect 48800 37780 48802 37820
rect 48510 37738 48634 37780
rect 48678 37738 48802 37780
rect 63630 37820 63754 37862
rect 63798 37820 63922 37862
rect 63630 37780 63632 37820
rect 63632 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63754 37820
rect 63798 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63920 37820
rect 63920 37780 63922 37820
rect 63630 37738 63754 37780
rect 63798 37738 63922 37780
rect 78750 37820 78874 37862
rect 78918 37820 79042 37862
rect 78750 37780 78752 37820
rect 78752 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78874 37820
rect 78918 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79040 37820
rect 79040 37780 79042 37820
rect 78750 37738 78874 37780
rect 78918 37738 79042 37780
rect 4390 37064 4514 37106
rect 4558 37064 4682 37106
rect 4390 37024 4392 37064
rect 4392 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4514 37064
rect 4558 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4680 37064
rect 4680 37024 4682 37064
rect 4390 36982 4514 37024
rect 4558 36982 4682 37024
rect 19510 37064 19634 37106
rect 19678 37064 19802 37106
rect 19510 37024 19512 37064
rect 19512 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19634 37064
rect 19678 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19800 37064
rect 19800 37024 19802 37064
rect 19510 36982 19634 37024
rect 19678 36982 19802 37024
rect 34630 37064 34754 37106
rect 34798 37064 34922 37106
rect 34630 37024 34632 37064
rect 34632 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34754 37064
rect 34798 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34920 37064
rect 34920 37024 34922 37064
rect 34630 36982 34754 37024
rect 34798 36982 34922 37024
rect 49750 37064 49874 37106
rect 49918 37064 50042 37106
rect 49750 37024 49752 37064
rect 49752 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49874 37064
rect 49918 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50040 37064
rect 50040 37024 50042 37064
rect 49750 36982 49874 37024
rect 49918 36982 50042 37024
rect 64870 37064 64994 37106
rect 65038 37064 65162 37106
rect 64870 37024 64872 37064
rect 64872 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64994 37064
rect 65038 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65160 37064
rect 65160 37024 65162 37064
rect 64870 36982 64994 37024
rect 65038 36982 65162 37024
rect 79990 37064 80114 37106
rect 80158 37064 80282 37106
rect 79990 37024 79992 37064
rect 79992 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80114 37064
rect 80158 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80280 37064
rect 80280 37024 80282 37064
rect 79990 36982 80114 37024
rect 80158 36982 80282 37024
rect 3150 36308 3274 36350
rect 3318 36308 3442 36350
rect 3150 36268 3152 36308
rect 3152 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3274 36308
rect 3318 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3440 36308
rect 3440 36268 3442 36308
rect 3150 36226 3274 36268
rect 3318 36226 3442 36268
rect 18270 36308 18394 36350
rect 18438 36308 18562 36350
rect 18270 36268 18272 36308
rect 18272 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18394 36308
rect 18438 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18560 36308
rect 18560 36268 18562 36308
rect 18270 36226 18394 36268
rect 18438 36226 18562 36268
rect 33390 36308 33514 36350
rect 33558 36308 33682 36350
rect 33390 36268 33392 36308
rect 33392 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33514 36308
rect 33558 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33680 36308
rect 33680 36268 33682 36308
rect 33390 36226 33514 36268
rect 33558 36226 33682 36268
rect 48510 36308 48634 36350
rect 48678 36308 48802 36350
rect 48510 36268 48512 36308
rect 48512 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48634 36308
rect 48678 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48800 36308
rect 48800 36268 48802 36308
rect 48510 36226 48634 36268
rect 48678 36226 48802 36268
rect 63630 36308 63754 36350
rect 63798 36308 63922 36350
rect 63630 36268 63632 36308
rect 63632 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63754 36308
rect 63798 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63920 36308
rect 63920 36268 63922 36308
rect 63630 36226 63754 36268
rect 63798 36226 63922 36268
rect 78750 36308 78874 36350
rect 78918 36308 79042 36350
rect 78750 36268 78752 36308
rect 78752 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78874 36308
rect 78918 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79040 36308
rect 79040 36268 79042 36308
rect 78750 36226 78874 36268
rect 78918 36226 79042 36268
rect 4390 35552 4514 35594
rect 4558 35552 4682 35594
rect 4390 35512 4392 35552
rect 4392 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4514 35552
rect 4558 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4680 35552
rect 4680 35512 4682 35552
rect 4390 35470 4514 35512
rect 4558 35470 4682 35512
rect 19510 35552 19634 35594
rect 19678 35552 19802 35594
rect 19510 35512 19512 35552
rect 19512 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19634 35552
rect 19678 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19800 35552
rect 19800 35512 19802 35552
rect 19510 35470 19634 35512
rect 19678 35470 19802 35512
rect 34630 35552 34754 35594
rect 34798 35552 34922 35594
rect 34630 35512 34632 35552
rect 34632 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34754 35552
rect 34798 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34920 35552
rect 34920 35512 34922 35552
rect 34630 35470 34754 35512
rect 34798 35470 34922 35512
rect 49750 35552 49874 35594
rect 49918 35552 50042 35594
rect 49750 35512 49752 35552
rect 49752 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49874 35552
rect 49918 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50040 35552
rect 50040 35512 50042 35552
rect 49750 35470 49874 35512
rect 49918 35470 50042 35512
rect 64870 35552 64994 35594
rect 65038 35552 65162 35594
rect 64870 35512 64872 35552
rect 64872 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64994 35552
rect 65038 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65160 35552
rect 65160 35512 65162 35552
rect 64870 35470 64994 35512
rect 65038 35470 65162 35512
rect 79990 35552 80114 35594
rect 80158 35552 80282 35594
rect 79990 35512 79992 35552
rect 79992 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80114 35552
rect 80158 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80280 35552
rect 80280 35512 80282 35552
rect 79990 35470 80114 35512
rect 80158 35470 80282 35512
rect 3150 34796 3274 34838
rect 3318 34796 3442 34838
rect 3150 34756 3152 34796
rect 3152 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3274 34796
rect 3318 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3440 34796
rect 3440 34756 3442 34796
rect 3150 34714 3274 34756
rect 3318 34714 3442 34756
rect 18270 34796 18394 34838
rect 18438 34796 18562 34838
rect 18270 34756 18272 34796
rect 18272 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18394 34796
rect 18438 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18560 34796
rect 18560 34756 18562 34796
rect 18270 34714 18394 34756
rect 18438 34714 18562 34756
rect 33390 34796 33514 34838
rect 33558 34796 33682 34838
rect 33390 34756 33392 34796
rect 33392 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33514 34796
rect 33558 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33680 34796
rect 33680 34756 33682 34796
rect 33390 34714 33514 34756
rect 33558 34714 33682 34756
rect 48510 34796 48634 34838
rect 48678 34796 48802 34838
rect 48510 34756 48512 34796
rect 48512 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48634 34796
rect 48678 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48800 34796
rect 48800 34756 48802 34796
rect 48510 34714 48634 34756
rect 48678 34714 48802 34756
rect 63630 34796 63754 34838
rect 63798 34796 63922 34838
rect 63630 34756 63632 34796
rect 63632 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63754 34796
rect 63798 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63920 34796
rect 63920 34756 63922 34796
rect 63630 34714 63754 34756
rect 63798 34714 63922 34756
rect 78750 34796 78874 34838
rect 78918 34796 79042 34838
rect 78750 34756 78752 34796
rect 78752 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78874 34796
rect 78918 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79040 34796
rect 79040 34756 79042 34796
rect 78750 34714 78874 34756
rect 78918 34714 79042 34756
rect 93870 34098 93994 34222
rect 94038 34098 94162 34222
rect 4390 34040 4514 34082
rect 4558 34040 4682 34082
rect 4390 34000 4392 34040
rect 4392 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4514 34040
rect 4558 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4680 34040
rect 4680 34000 4682 34040
rect 4390 33958 4514 34000
rect 4558 33958 4682 34000
rect 19510 34040 19634 34082
rect 19678 34040 19802 34082
rect 19510 34000 19512 34040
rect 19512 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19634 34040
rect 19678 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19800 34040
rect 19800 34000 19802 34040
rect 19510 33958 19634 34000
rect 19678 33958 19802 34000
rect 34630 34040 34754 34082
rect 34798 34040 34922 34082
rect 34630 34000 34632 34040
rect 34632 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34754 34040
rect 34798 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34920 34040
rect 34920 34000 34922 34040
rect 34630 33958 34754 34000
rect 34798 33958 34922 34000
rect 49750 34040 49874 34082
rect 49918 34040 50042 34082
rect 49750 34000 49752 34040
rect 49752 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49874 34040
rect 49918 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50040 34040
rect 50040 34000 50042 34040
rect 49750 33958 49874 34000
rect 49918 33958 50042 34000
rect 64870 34040 64994 34082
rect 65038 34040 65162 34082
rect 64870 34000 64872 34040
rect 64872 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64994 34040
rect 65038 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65160 34040
rect 65160 34000 65162 34040
rect 64870 33958 64994 34000
rect 65038 33958 65162 34000
rect 79990 34040 80114 34082
rect 80158 34040 80282 34082
rect 79990 34000 79992 34040
rect 79992 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80114 34040
rect 80158 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80280 34040
rect 80280 34000 80282 34040
rect 79990 33958 80114 34000
rect 80158 33958 80282 34000
rect 93870 33930 93994 34054
rect 94038 33930 94162 34054
rect 67298 33790 67422 33914
rect 3150 33284 3274 33326
rect 3318 33284 3442 33326
rect 3150 33244 3152 33284
rect 3152 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3274 33284
rect 3318 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3440 33284
rect 3440 33244 3442 33284
rect 3150 33202 3274 33244
rect 3318 33202 3442 33244
rect 78750 33284 78874 33326
rect 78918 33284 79042 33326
rect 78750 33244 78752 33284
rect 78752 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78874 33284
rect 78918 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79040 33284
rect 79040 33244 79042 33284
rect 78750 33202 78874 33244
rect 78918 33202 79042 33244
rect 4390 32528 4514 32570
rect 4558 32528 4682 32570
rect 4390 32488 4392 32528
rect 4392 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4514 32528
rect 4558 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4680 32528
rect 4680 32488 4682 32528
rect 4390 32446 4514 32488
rect 4558 32446 4682 32488
rect 79990 32528 80114 32570
rect 80158 32528 80282 32570
rect 79990 32488 79992 32528
rect 79992 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80114 32528
rect 80158 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80280 32528
rect 80280 32488 80282 32528
rect 79990 32446 80114 32488
rect 80158 32446 80282 32488
rect 3150 31772 3274 31814
rect 3318 31772 3442 31814
rect 3150 31732 3152 31772
rect 3152 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3274 31772
rect 3318 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3440 31772
rect 3440 31732 3442 31772
rect 3150 31690 3274 31732
rect 3318 31690 3442 31732
rect 78750 31772 78874 31814
rect 78918 31772 79042 31814
rect 78750 31732 78752 31772
rect 78752 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78874 31772
rect 78918 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79040 31772
rect 79040 31732 79042 31772
rect 78750 31690 78874 31732
rect 78918 31690 79042 31732
rect 4390 31016 4514 31058
rect 4558 31016 4682 31058
rect 4390 30976 4392 31016
rect 4392 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4514 31016
rect 4558 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4680 31016
rect 4680 30976 4682 31016
rect 4390 30934 4514 30976
rect 4558 30934 4682 30976
rect 79990 31016 80114 31058
rect 80158 31016 80282 31058
rect 79990 30976 79992 31016
rect 79992 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80114 31016
rect 80158 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80280 31016
rect 80280 30976 80282 31016
rect 79990 30934 80114 30976
rect 80158 30934 80282 30976
rect 3150 30260 3274 30302
rect 3318 30260 3442 30302
rect 3150 30220 3152 30260
rect 3152 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3274 30260
rect 3318 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3440 30260
rect 3440 30220 3442 30260
rect 3150 30178 3274 30220
rect 3318 30178 3442 30220
rect 78750 30260 78874 30302
rect 78918 30260 79042 30302
rect 78750 30220 78752 30260
rect 78752 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78874 30260
rect 78918 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79040 30260
rect 79040 30220 79042 30260
rect 78750 30178 78874 30220
rect 78918 30178 79042 30220
rect 66386 29926 66510 30050
rect 4390 29504 4514 29546
rect 4558 29504 4682 29546
rect 4390 29464 4392 29504
rect 4392 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4514 29504
rect 4558 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4680 29504
rect 4680 29464 4682 29504
rect 4390 29422 4514 29464
rect 4558 29422 4682 29464
rect 79990 29504 80114 29546
rect 80158 29504 80282 29546
rect 79990 29464 79992 29504
rect 79992 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80114 29504
rect 80158 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80280 29504
rect 80280 29464 80282 29504
rect 79990 29422 80114 29464
rect 80158 29422 80282 29464
rect 95110 29338 95234 29462
rect 95278 29338 95402 29462
rect 95110 29170 95234 29294
rect 95278 29170 95402 29294
rect 18270 28898 18394 29022
rect 18438 28898 18562 29022
rect 3150 28748 3274 28790
rect 3318 28748 3442 28790
rect 3150 28708 3152 28748
rect 3152 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3274 28748
rect 3318 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3440 28748
rect 3440 28708 3442 28748
rect 3150 28666 3274 28708
rect 3318 28666 3442 28708
rect 18270 28730 18394 28854
rect 18438 28730 18562 28854
rect 33390 28898 33514 29022
rect 33558 28898 33682 29022
rect 33390 28730 33514 28854
rect 33558 28730 33682 28854
rect 48510 28898 48634 29022
rect 48678 28898 48802 29022
rect 48510 28730 48634 28854
rect 48678 28730 48802 28854
rect 63630 28898 63754 29022
rect 63798 28898 63922 29022
rect 63630 28730 63754 28854
rect 63798 28730 63922 28854
rect 78750 28748 78874 28790
rect 78918 28748 79042 28790
rect 78750 28708 78752 28748
rect 78752 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78874 28748
rect 78918 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79040 28748
rect 79040 28708 79042 28748
rect 78750 28666 78874 28708
rect 78918 28666 79042 28708
rect 93870 28098 93994 28222
rect 94038 28098 94162 28222
rect 4390 27992 4514 28034
rect 4558 27992 4682 28034
rect 4390 27952 4392 27992
rect 4392 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4514 27992
rect 4558 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4680 27992
rect 4680 27952 4682 27992
rect 4390 27910 4514 27952
rect 4558 27910 4682 27952
rect 79990 27992 80114 28034
rect 80158 27992 80282 28034
rect 79990 27952 79992 27992
rect 79992 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80114 27992
rect 80158 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80280 27992
rect 80280 27952 80282 27992
rect 79990 27910 80114 27952
rect 80158 27910 80282 27952
rect 93870 27930 93994 28054
rect 94038 27930 94162 28054
rect 3150 27236 3274 27278
rect 3318 27236 3442 27278
rect 3150 27196 3152 27236
rect 3152 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3274 27236
rect 3318 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3440 27236
rect 3440 27196 3442 27236
rect 3150 27154 3274 27196
rect 3318 27154 3442 27196
rect 78750 27236 78874 27278
rect 78918 27236 79042 27278
rect 78750 27196 78752 27236
rect 78752 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78874 27236
rect 78918 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79040 27236
rect 79040 27196 79042 27236
rect 78750 27154 78874 27196
rect 78918 27154 79042 27196
rect 4390 26480 4514 26522
rect 4558 26480 4682 26522
rect 4390 26440 4392 26480
rect 4392 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4514 26480
rect 4558 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4680 26480
rect 4680 26440 4682 26480
rect 4390 26398 4514 26440
rect 4558 26398 4682 26440
rect 79990 26480 80114 26522
rect 80158 26480 80282 26522
rect 79990 26440 79992 26480
rect 79992 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80114 26480
rect 80158 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80280 26480
rect 80280 26440 80282 26480
rect 79990 26398 80114 26440
rect 80158 26398 80282 26440
rect 3150 25724 3274 25766
rect 3318 25724 3442 25766
rect 3150 25684 3152 25724
rect 3152 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3274 25724
rect 3318 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3440 25724
rect 3440 25684 3442 25724
rect 3150 25642 3274 25684
rect 3318 25642 3442 25684
rect 78750 25724 78874 25766
rect 78918 25724 79042 25766
rect 78750 25684 78752 25724
rect 78752 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78874 25724
rect 78918 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79040 25724
rect 79040 25684 79042 25724
rect 78750 25642 78874 25684
rect 78918 25642 79042 25684
rect 4390 24968 4514 25010
rect 4558 24968 4682 25010
rect 4390 24928 4392 24968
rect 4392 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4514 24968
rect 4558 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4680 24968
rect 4680 24928 4682 24968
rect 4390 24886 4514 24928
rect 4558 24886 4682 24928
rect 79990 24968 80114 25010
rect 80158 24968 80282 25010
rect 79990 24928 79992 24968
rect 79992 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80114 24968
rect 80158 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80280 24968
rect 80280 24928 80282 24968
rect 79990 24886 80114 24928
rect 80158 24886 80282 24928
rect 3150 24212 3274 24254
rect 3318 24212 3442 24254
rect 3150 24172 3152 24212
rect 3152 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3274 24212
rect 3318 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3440 24212
rect 3440 24172 3442 24212
rect 3150 24130 3274 24172
rect 3318 24130 3442 24172
rect 19510 24138 19634 24262
rect 19678 24138 19802 24262
rect 19510 23970 19634 24094
rect 19678 23970 19802 24094
rect 34630 24138 34754 24262
rect 34798 24138 34922 24262
rect 34630 23970 34754 24094
rect 34798 23970 34922 24094
rect 49750 24138 49874 24262
rect 49918 24138 50042 24262
rect 49750 23970 49874 24094
rect 49918 23970 50042 24094
rect 64870 24138 64994 24262
rect 65038 24138 65162 24262
rect 78750 24212 78874 24254
rect 78918 24212 79042 24254
rect 78750 24172 78752 24212
rect 78752 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78874 24212
rect 78918 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79040 24212
rect 79040 24172 79042 24212
rect 78750 24130 78874 24172
rect 78918 24130 79042 24172
rect 64870 23970 64994 24094
rect 65038 23970 65162 24094
rect 4390 23456 4514 23498
rect 4558 23456 4682 23498
rect 4390 23416 4392 23456
rect 4392 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4514 23456
rect 4558 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4680 23456
rect 4680 23416 4682 23456
rect 4390 23374 4514 23416
rect 4558 23374 4682 23416
rect 79990 23456 80114 23498
rect 80158 23456 80282 23498
rect 79990 23416 79992 23456
rect 79992 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80114 23456
rect 80158 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80280 23456
rect 80280 23416 80282 23456
rect 79990 23374 80114 23416
rect 80158 23374 80282 23416
rect 18270 22898 18394 23022
rect 18438 22898 18562 23022
rect 3150 22700 3274 22742
rect 3318 22700 3442 22742
rect 3150 22660 3152 22700
rect 3152 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3274 22700
rect 3318 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3440 22700
rect 3440 22660 3442 22700
rect 3150 22618 3274 22660
rect 3318 22618 3442 22660
rect 18270 22730 18394 22854
rect 18438 22730 18562 22854
rect 33390 22898 33514 23022
rect 33558 22898 33682 23022
rect 33390 22730 33514 22854
rect 33558 22730 33682 22854
rect 48510 22898 48634 23022
rect 48678 22898 48802 23022
rect 48510 22730 48634 22854
rect 48678 22730 48802 22854
rect 63630 22898 63754 23022
rect 63798 22898 63922 23022
rect 63630 22730 63754 22854
rect 63798 22730 63922 22854
rect 78750 22700 78874 22742
rect 78918 22700 79042 22742
rect 78750 22660 78752 22700
rect 78752 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78874 22700
rect 78918 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79040 22700
rect 79040 22660 79042 22700
rect 78750 22618 78874 22660
rect 78918 22618 79042 22660
rect 4390 21944 4514 21986
rect 4558 21944 4682 21986
rect 4390 21904 4392 21944
rect 4392 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4514 21944
rect 4558 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4680 21944
rect 4680 21904 4682 21944
rect 4390 21862 4514 21904
rect 4558 21862 4682 21904
rect 79990 21944 80114 21986
rect 80158 21944 80282 21986
rect 79990 21904 79992 21944
rect 79992 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80114 21944
rect 80158 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80280 21944
rect 80280 21904 80282 21944
rect 79990 21862 80114 21904
rect 80158 21862 80282 21904
rect 95110 21944 95234 21986
rect 95278 21944 95402 21986
rect 95110 21904 95112 21944
rect 95112 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95234 21944
rect 95278 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95400 21944
rect 95400 21904 95402 21944
rect 95110 21862 95234 21904
rect 95278 21862 95402 21904
rect 3150 21188 3274 21230
rect 3318 21188 3442 21230
rect 3150 21148 3152 21188
rect 3152 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3274 21188
rect 3318 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3440 21188
rect 3440 21148 3442 21188
rect 3150 21106 3274 21148
rect 3318 21106 3442 21148
rect 78750 21188 78874 21230
rect 78918 21188 79042 21230
rect 78750 21148 78752 21188
rect 78752 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78874 21188
rect 78918 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79040 21188
rect 79040 21148 79042 21188
rect 78750 21106 78874 21148
rect 78918 21106 79042 21148
rect 93870 21188 93994 21230
rect 94038 21188 94162 21230
rect 93870 21148 93872 21188
rect 93872 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93994 21188
rect 94038 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94160 21188
rect 94160 21148 94162 21188
rect 93870 21106 93994 21148
rect 94038 21106 94162 21148
rect 4390 20432 4514 20474
rect 4558 20432 4682 20474
rect 4390 20392 4392 20432
rect 4392 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4514 20432
rect 4558 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4680 20432
rect 4680 20392 4682 20432
rect 4390 20350 4514 20392
rect 4558 20350 4682 20392
rect 79990 20432 80114 20474
rect 80158 20432 80282 20474
rect 79990 20392 79992 20432
rect 79992 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80114 20432
rect 80158 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80280 20432
rect 80280 20392 80282 20432
rect 79990 20350 80114 20392
rect 80158 20350 80282 20392
rect 95110 20432 95234 20474
rect 95278 20432 95402 20474
rect 95110 20392 95112 20432
rect 95112 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95234 20432
rect 95278 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95400 20432
rect 95400 20392 95402 20432
rect 95110 20350 95234 20392
rect 95278 20350 95402 20392
rect 3150 19676 3274 19718
rect 3318 19676 3442 19718
rect 3150 19636 3152 19676
rect 3152 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3274 19676
rect 3318 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3440 19676
rect 3440 19636 3442 19676
rect 3150 19594 3274 19636
rect 3318 19594 3442 19636
rect 78750 19676 78874 19718
rect 78918 19676 79042 19718
rect 78750 19636 78752 19676
rect 78752 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78874 19676
rect 78918 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79040 19676
rect 79040 19636 79042 19676
rect 78750 19594 78874 19636
rect 78918 19594 79042 19636
rect 93870 19676 93994 19718
rect 94038 19676 94162 19718
rect 93870 19636 93872 19676
rect 93872 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93994 19676
rect 94038 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94160 19676
rect 94160 19636 94162 19676
rect 93870 19594 93994 19636
rect 94038 19594 94162 19636
rect 4390 18920 4514 18962
rect 4558 18920 4682 18962
rect 4390 18880 4392 18920
rect 4392 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4514 18920
rect 4558 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4680 18920
rect 4680 18880 4682 18920
rect 4390 18838 4514 18880
rect 4558 18838 4682 18880
rect 79990 18920 80114 18962
rect 80158 18920 80282 18962
rect 79990 18880 79992 18920
rect 79992 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80114 18920
rect 80158 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80280 18920
rect 80280 18880 80282 18920
rect 79990 18838 80114 18880
rect 80158 18838 80282 18880
rect 3150 18164 3274 18206
rect 3318 18164 3442 18206
rect 3150 18124 3152 18164
rect 3152 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3274 18164
rect 3318 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3440 18164
rect 3440 18124 3442 18164
rect 3150 18082 3274 18124
rect 3318 18082 3442 18124
rect 19510 18138 19634 18262
rect 19678 18138 19802 18262
rect 19510 17970 19634 18094
rect 19678 17970 19802 18094
rect 34630 18138 34754 18262
rect 34798 18138 34922 18262
rect 34630 17970 34754 18094
rect 34798 17970 34922 18094
rect 49750 18138 49874 18262
rect 49918 18138 50042 18262
rect 49750 17970 49874 18094
rect 49918 17970 50042 18094
rect 64870 18138 64994 18262
rect 65038 18138 65162 18262
rect 64870 17970 64994 18094
rect 65038 17970 65162 18094
rect 78750 18164 78874 18206
rect 78918 18164 79042 18206
rect 78750 18124 78752 18164
rect 78752 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78874 18164
rect 78918 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79040 18164
rect 79040 18124 79042 18164
rect 78750 18082 78874 18124
rect 78918 18082 79042 18124
rect 4390 17408 4514 17450
rect 4558 17408 4682 17450
rect 4390 17368 4392 17408
rect 4392 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4514 17408
rect 4558 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4680 17408
rect 4680 17368 4682 17408
rect 4390 17326 4514 17368
rect 4558 17326 4682 17368
rect 79990 17408 80114 17450
rect 80158 17408 80282 17450
rect 79990 17368 79992 17408
rect 79992 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80114 17408
rect 80158 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80280 17408
rect 80280 17368 80282 17408
rect 79990 17326 80114 17368
rect 80158 17326 80282 17368
rect 18270 16898 18394 17022
rect 18438 16898 18562 17022
rect 18270 16730 18394 16854
rect 18438 16730 18562 16854
rect 3150 16652 3274 16694
rect 3318 16652 3442 16694
rect 33390 16898 33514 17022
rect 33558 16898 33682 17022
rect 33390 16730 33514 16854
rect 33558 16730 33682 16854
rect 48510 16898 48634 17022
rect 48678 16898 48802 17022
rect 48510 16730 48634 16854
rect 48678 16730 48802 16854
rect 63630 16898 63754 17022
rect 63798 16898 63922 17022
rect 63630 16730 63754 16854
rect 63798 16730 63922 16854
rect 3150 16612 3152 16652
rect 3152 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3274 16652
rect 3318 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3440 16652
rect 3440 16612 3442 16652
rect 3150 16570 3274 16612
rect 3318 16570 3442 16612
rect 78750 16652 78874 16694
rect 78918 16652 79042 16694
rect 78750 16612 78752 16652
rect 78752 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78874 16652
rect 78918 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79040 16652
rect 79040 16612 79042 16652
rect 78750 16570 78874 16612
rect 78918 16570 79042 16612
rect 4390 15896 4514 15938
rect 4558 15896 4682 15938
rect 4390 15856 4392 15896
rect 4392 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4514 15896
rect 4558 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4680 15896
rect 4680 15856 4682 15896
rect 4390 15814 4514 15856
rect 4558 15814 4682 15856
rect 79990 15896 80114 15938
rect 80158 15896 80282 15938
rect 79990 15856 79992 15896
rect 79992 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80114 15896
rect 80158 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80280 15896
rect 80280 15856 80282 15896
rect 79990 15814 80114 15856
rect 80158 15814 80282 15856
rect 3150 15140 3274 15182
rect 3318 15140 3442 15182
rect 3150 15100 3152 15140
rect 3152 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3274 15140
rect 3318 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3440 15140
rect 3440 15100 3442 15140
rect 3150 15058 3274 15100
rect 3318 15058 3442 15100
rect 78750 15140 78874 15182
rect 78918 15140 79042 15182
rect 78750 15100 78752 15140
rect 78752 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78874 15140
rect 78918 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79040 15140
rect 79040 15100 79042 15140
rect 78750 15058 78874 15100
rect 78918 15058 79042 15100
rect 4390 14384 4514 14426
rect 4558 14384 4682 14426
rect 4390 14344 4392 14384
rect 4392 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4514 14384
rect 4558 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4680 14384
rect 4680 14344 4682 14384
rect 4390 14302 4514 14344
rect 4558 14302 4682 14344
rect 79990 14384 80114 14426
rect 80158 14384 80282 14426
rect 79990 14344 79992 14384
rect 79992 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80114 14384
rect 80158 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80280 14384
rect 80280 14344 80282 14384
rect 79990 14302 80114 14344
rect 80158 14302 80282 14344
rect 3150 13628 3274 13670
rect 3318 13628 3442 13670
rect 3150 13588 3152 13628
rect 3152 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3274 13628
rect 3318 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3440 13628
rect 3440 13588 3442 13628
rect 3150 13546 3274 13588
rect 3318 13546 3442 13588
rect 78750 13628 78874 13670
rect 78918 13628 79042 13670
rect 78750 13588 78752 13628
rect 78752 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78874 13628
rect 78918 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79040 13628
rect 79040 13588 79042 13628
rect 78750 13546 78874 13588
rect 78918 13546 79042 13588
rect 4390 12872 4514 12914
rect 4558 12872 4682 12914
rect 4390 12832 4392 12872
rect 4392 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4514 12872
rect 4558 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4680 12872
rect 4680 12832 4682 12872
rect 4390 12790 4514 12832
rect 4558 12790 4682 12832
rect 79990 12872 80114 12914
rect 80158 12872 80282 12914
rect 79990 12832 79992 12872
rect 79992 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80114 12872
rect 80158 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80280 12872
rect 80280 12832 80282 12872
rect 79990 12790 80114 12832
rect 80158 12790 80282 12832
rect 3150 12116 3274 12158
rect 3318 12116 3442 12158
rect 3150 12076 3152 12116
rect 3152 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3274 12116
rect 3318 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3440 12116
rect 3440 12076 3442 12116
rect 3150 12034 3274 12076
rect 3318 12034 3442 12076
rect 19510 12138 19634 12262
rect 19678 12138 19802 12262
rect 19510 11970 19634 12094
rect 19678 11970 19802 12094
rect 34630 12138 34754 12262
rect 34798 12138 34922 12262
rect 34630 11970 34754 12094
rect 34798 11970 34922 12094
rect 49750 12138 49874 12262
rect 49918 12138 50042 12262
rect 49750 11970 49874 12094
rect 49918 11970 50042 12094
rect 64870 12138 64994 12262
rect 65038 12138 65162 12262
rect 64870 11970 64994 12094
rect 65038 11970 65162 12094
rect 78750 12116 78874 12158
rect 78918 12116 79042 12158
rect 78750 12076 78752 12116
rect 78752 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78874 12116
rect 78918 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79040 12116
rect 79040 12076 79042 12116
rect 78750 12034 78874 12076
rect 78918 12034 79042 12076
rect 95110 12138 95234 12262
rect 95278 12138 95402 12262
rect 95110 11970 95234 12094
rect 95278 11970 95402 12094
rect 4390 11360 4514 11402
rect 4558 11360 4682 11402
rect 4390 11320 4392 11360
rect 4392 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4514 11360
rect 4558 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4680 11360
rect 4680 11320 4682 11360
rect 4390 11278 4514 11320
rect 4558 11278 4682 11320
rect 79990 11360 80114 11402
rect 80158 11360 80282 11402
rect 79990 11320 79992 11360
rect 79992 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80114 11360
rect 80158 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80280 11360
rect 80280 11320 80282 11360
rect 79990 11278 80114 11320
rect 80158 11278 80282 11320
rect 18270 10898 18394 11022
rect 18438 10898 18562 11022
rect 18270 10730 18394 10854
rect 18438 10730 18562 10854
rect 33390 10898 33514 11022
rect 33558 10898 33682 11022
rect 33390 10730 33514 10854
rect 33558 10730 33682 10854
rect 48510 10898 48634 11022
rect 48678 10898 48802 11022
rect 48510 10730 48634 10854
rect 48678 10730 48802 10854
rect 63630 10898 63754 11022
rect 63798 10898 63922 11022
rect 63630 10730 63754 10854
rect 63798 10730 63922 10854
rect 93870 10898 93994 11022
rect 94038 10898 94162 11022
rect 93870 10730 93994 10854
rect 94038 10730 94162 10854
rect 3150 10604 3274 10646
rect 3318 10604 3442 10646
rect 3150 10564 3152 10604
rect 3152 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3274 10604
rect 3318 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3440 10604
rect 3440 10564 3442 10604
rect 3150 10522 3274 10564
rect 3318 10522 3442 10564
rect 78750 10604 78874 10646
rect 78918 10604 79042 10646
rect 78750 10564 78752 10604
rect 78752 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78874 10604
rect 78918 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79040 10604
rect 79040 10564 79042 10604
rect 78750 10522 78874 10564
rect 78918 10522 79042 10564
rect 4390 9848 4514 9890
rect 4558 9848 4682 9890
rect 4390 9808 4392 9848
rect 4392 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4514 9848
rect 4558 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4680 9848
rect 4680 9808 4682 9848
rect 4390 9766 4514 9808
rect 4558 9766 4682 9808
rect 79990 9848 80114 9890
rect 80158 9848 80282 9890
rect 79990 9808 79992 9848
rect 79992 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80114 9848
rect 80158 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80280 9848
rect 80280 9808 80282 9848
rect 79990 9766 80114 9808
rect 80158 9766 80282 9808
rect 3150 9092 3274 9134
rect 3318 9092 3442 9134
rect 3150 9052 3152 9092
rect 3152 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3274 9092
rect 3318 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3440 9092
rect 3440 9052 3442 9092
rect 3150 9010 3274 9052
rect 3318 9010 3442 9052
rect 78750 9092 78874 9134
rect 78918 9092 79042 9134
rect 78750 9052 78752 9092
rect 78752 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78874 9092
rect 78918 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79040 9092
rect 79040 9052 79042 9092
rect 78750 9010 78874 9052
rect 78918 9010 79042 9052
rect 4390 8336 4514 8378
rect 4558 8336 4682 8378
rect 4390 8296 4392 8336
rect 4392 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4514 8336
rect 4558 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4680 8336
rect 4680 8296 4682 8336
rect 4390 8254 4514 8296
rect 4558 8254 4682 8296
rect 79990 8336 80114 8378
rect 80158 8336 80282 8378
rect 79990 8296 79992 8336
rect 79992 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80114 8336
rect 80158 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80280 8336
rect 80280 8296 80282 8336
rect 79990 8254 80114 8296
rect 80158 8254 80282 8296
rect 3150 7580 3274 7622
rect 3318 7580 3442 7622
rect 3150 7540 3152 7580
rect 3152 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3274 7580
rect 3318 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3440 7580
rect 3440 7540 3442 7580
rect 3150 7498 3274 7540
rect 3318 7498 3442 7540
rect 78750 7580 78874 7622
rect 78918 7580 79042 7622
rect 78750 7540 78752 7580
rect 78752 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78874 7580
rect 78918 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79040 7580
rect 79040 7540 79042 7580
rect 78750 7498 78874 7540
rect 78918 7498 79042 7540
rect 4390 6824 4514 6866
rect 4558 6824 4682 6866
rect 4390 6784 4392 6824
rect 4392 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4514 6824
rect 4558 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4680 6824
rect 4680 6784 4682 6824
rect 4390 6742 4514 6784
rect 4558 6742 4682 6784
rect 79990 6824 80114 6866
rect 80158 6824 80282 6866
rect 79990 6784 79992 6824
rect 79992 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80114 6824
rect 80158 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80280 6824
rect 80280 6784 80282 6824
rect 79990 6742 80114 6784
rect 80158 6742 80282 6784
rect 95110 6138 95234 6262
rect 95278 6138 95402 6262
rect 3150 6068 3274 6110
rect 3318 6068 3442 6110
rect 3150 6028 3152 6068
rect 3152 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3274 6068
rect 3318 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3440 6068
rect 3440 6028 3442 6068
rect 3150 5986 3274 6028
rect 3318 5986 3442 6028
rect 78750 6068 78874 6110
rect 78918 6068 79042 6110
rect 78750 6028 78752 6068
rect 78752 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78874 6068
rect 78918 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79040 6068
rect 79040 6028 79042 6068
rect 78750 5986 78874 6028
rect 78918 5986 79042 6028
rect 95110 5970 95234 6094
rect 95278 5970 95402 6094
rect 67298 5650 67422 5774
rect 4390 5312 4514 5354
rect 4558 5312 4682 5354
rect 4390 5272 4392 5312
rect 4392 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4514 5312
rect 4558 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4680 5312
rect 4680 5272 4682 5312
rect 4390 5230 4514 5272
rect 4558 5230 4682 5272
rect 19510 5312 19634 5354
rect 19678 5312 19802 5354
rect 19510 5272 19512 5312
rect 19512 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19634 5312
rect 19678 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19800 5312
rect 19800 5272 19802 5312
rect 19510 5230 19634 5272
rect 19678 5230 19802 5272
rect 34630 5312 34754 5354
rect 34798 5312 34922 5354
rect 34630 5272 34632 5312
rect 34632 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34754 5312
rect 34798 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34920 5312
rect 34920 5272 34922 5312
rect 34630 5230 34754 5272
rect 34798 5230 34922 5272
rect 49750 5312 49874 5354
rect 49918 5312 50042 5354
rect 49750 5272 49752 5312
rect 49752 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49874 5312
rect 49918 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50040 5312
rect 50040 5272 50042 5312
rect 49750 5230 49874 5272
rect 49918 5230 50042 5272
rect 64870 5312 64994 5354
rect 65038 5312 65162 5354
rect 64870 5272 64872 5312
rect 64872 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64994 5312
rect 65038 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65160 5312
rect 65160 5272 65162 5312
rect 64870 5230 64994 5272
rect 65038 5230 65162 5272
rect 79990 5312 80114 5354
rect 80158 5312 80282 5354
rect 79990 5272 79992 5312
rect 79992 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80114 5312
rect 80158 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80280 5312
rect 80280 5272 80282 5312
rect 79990 5230 80114 5272
rect 80158 5230 80282 5272
rect 93870 4898 93994 5022
rect 94038 4898 94162 5022
rect 66386 4642 66510 4766
rect 93870 4730 93994 4854
rect 94038 4730 94162 4854
rect 3150 4556 3274 4598
rect 3318 4556 3442 4598
rect 3150 4516 3152 4556
rect 3152 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3274 4556
rect 3318 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3440 4556
rect 3440 4516 3442 4556
rect 3150 4474 3274 4516
rect 3318 4474 3442 4516
rect 18270 4556 18394 4598
rect 18438 4556 18562 4598
rect 18270 4516 18272 4556
rect 18272 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18394 4556
rect 18438 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18560 4556
rect 18560 4516 18562 4556
rect 18270 4474 18394 4516
rect 18438 4474 18562 4516
rect 33390 4556 33514 4598
rect 33558 4556 33682 4598
rect 33390 4516 33392 4556
rect 33392 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33514 4556
rect 33558 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33680 4556
rect 33680 4516 33682 4556
rect 33390 4474 33514 4516
rect 33558 4474 33682 4516
rect 48510 4556 48634 4598
rect 48678 4556 48802 4598
rect 48510 4516 48512 4556
rect 48512 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48634 4556
rect 48678 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48800 4556
rect 48800 4516 48802 4556
rect 48510 4474 48634 4516
rect 48678 4474 48802 4516
rect 63630 4556 63754 4598
rect 63798 4556 63922 4598
rect 63630 4516 63632 4556
rect 63632 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63754 4556
rect 63798 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63920 4556
rect 63920 4516 63922 4556
rect 63630 4474 63754 4516
rect 63798 4474 63922 4516
rect 78750 4556 78874 4598
rect 78918 4556 79042 4598
rect 78750 4516 78752 4556
rect 78752 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78874 4556
rect 78918 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79040 4556
rect 79040 4516 79042 4556
rect 78750 4474 78874 4516
rect 78918 4474 79042 4516
rect 4390 3800 4514 3842
rect 4558 3800 4682 3842
rect 4390 3760 4392 3800
rect 4392 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4514 3800
rect 4558 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4680 3800
rect 4680 3760 4682 3800
rect 4390 3718 4514 3760
rect 4558 3718 4682 3760
rect 19510 3800 19634 3842
rect 19678 3800 19802 3842
rect 19510 3760 19512 3800
rect 19512 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19634 3800
rect 19678 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19800 3800
rect 19800 3760 19802 3800
rect 19510 3718 19634 3760
rect 19678 3718 19802 3760
rect 34630 3800 34754 3842
rect 34798 3800 34922 3842
rect 34630 3760 34632 3800
rect 34632 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34754 3800
rect 34798 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34920 3800
rect 34920 3760 34922 3800
rect 34630 3718 34754 3760
rect 34798 3718 34922 3760
rect 49750 3800 49874 3842
rect 49918 3800 50042 3842
rect 49750 3760 49752 3800
rect 49752 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49874 3800
rect 49918 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50040 3800
rect 50040 3760 50042 3800
rect 49750 3718 49874 3760
rect 49918 3718 50042 3760
rect 64870 3800 64994 3842
rect 65038 3800 65162 3842
rect 64870 3760 64872 3800
rect 64872 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64994 3800
rect 65038 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65160 3800
rect 65160 3760 65162 3800
rect 64870 3718 64994 3760
rect 65038 3718 65162 3760
rect 79990 3800 80114 3842
rect 80158 3800 80282 3842
rect 79990 3760 79992 3800
rect 79992 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80114 3800
rect 80158 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80280 3800
rect 80280 3760 80282 3800
rect 79990 3718 80114 3760
rect 80158 3718 80282 3760
rect 3150 3044 3274 3086
rect 3318 3044 3442 3086
rect 3150 3004 3152 3044
rect 3152 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3274 3044
rect 3318 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3440 3044
rect 3440 3004 3442 3044
rect 3150 2962 3274 3004
rect 3318 2962 3442 3004
rect 18270 3044 18394 3086
rect 18438 3044 18562 3086
rect 18270 3004 18272 3044
rect 18272 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18394 3044
rect 18438 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18560 3044
rect 18560 3004 18562 3044
rect 18270 2962 18394 3004
rect 18438 2962 18562 3004
rect 33390 3044 33514 3086
rect 33558 3044 33682 3086
rect 33390 3004 33392 3044
rect 33392 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33514 3044
rect 33558 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33680 3044
rect 33680 3004 33682 3044
rect 33390 2962 33514 3004
rect 33558 2962 33682 3004
rect 48510 3044 48634 3086
rect 48678 3044 48802 3086
rect 48510 3004 48512 3044
rect 48512 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48634 3044
rect 48678 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48800 3044
rect 48800 3004 48802 3044
rect 48510 2962 48634 3004
rect 48678 2962 48802 3004
rect 63630 3044 63754 3086
rect 63798 3044 63922 3086
rect 63630 3004 63632 3044
rect 63632 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63754 3044
rect 63798 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63920 3044
rect 63920 3004 63922 3044
rect 63630 2962 63754 3004
rect 63798 2962 63922 3004
rect 78750 3044 78874 3086
rect 78918 3044 79042 3086
rect 78750 3004 78752 3044
rect 78752 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78874 3044
rect 78918 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79040 3044
rect 79040 3004 79042 3044
rect 78750 2962 78874 3004
rect 78918 2962 79042 3004
rect 4390 2288 4514 2330
rect 4558 2288 4682 2330
rect 4390 2248 4392 2288
rect 4392 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4514 2288
rect 4558 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4680 2288
rect 4680 2248 4682 2288
rect 4390 2206 4514 2248
rect 4558 2206 4682 2248
rect 19510 2288 19634 2330
rect 19678 2288 19802 2330
rect 19510 2248 19512 2288
rect 19512 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19634 2288
rect 19678 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19800 2288
rect 19800 2248 19802 2288
rect 19510 2206 19634 2248
rect 19678 2206 19802 2248
rect 34630 2288 34754 2330
rect 34798 2288 34922 2330
rect 34630 2248 34632 2288
rect 34632 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34754 2288
rect 34798 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34920 2288
rect 34920 2248 34922 2288
rect 34630 2206 34754 2248
rect 34798 2206 34922 2248
rect 49750 2288 49874 2330
rect 49918 2288 50042 2330
rect 49750 2248 49752 2288
rect 49752 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49874 2288
rect 49918 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50040 2288
rect 50040 2248 50042 2288
rect 49750 2206 49874 2248
rect 49918 2206 50042 2248
rect 64870 2288 64994 2330
rect 65038 2288 65162 2330
rect 64870 2248 64872 2288
rect 64872 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64994 2288
rect 65038 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65160 2288
rect 65160 2248 65162 2288
rect 64870 2206 64994 2248
rect 65038 2206 65162 2248
rect 79990 2288 80114 2330
rect 80158 2288 80282 2330
rect 79990 2248 79992 2288
rect 79992 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80114 2288
rect 80158 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80280 2288
rect 80280 2248 80282 2288
rect 79990 2206 80114 2248
rect 80158 2206 80282 2248
rect 3150 1532 3274 1574
rect 3318 1532 3442 1574
rect 3150 1492 3152 1532
rect 3152 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3274 1532
rect 3318 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3440 1532
rect 3440 1492 3442 1532
rect 3150 1450 3274 1492
rect 3318 1450 3442 1492
rect 18270 1532 18394 1574
rect 18438 1532 18562 1574
rect 18270 1492 18272 1532
rect 18272 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18394 1532
rect 18438 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18560 1532
rect 18560 1492 18562 1532
rect 18270 1450 18394 1492
rect 18438 1450 18562 1492
rect 33390 1532 33514 1574
rect 33558 1532 33682 1574
rect 33390 1492 33392 1532
rect 33392 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33514 1532
rect 33558 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33680 1532
rect 33680 1492 33682 1532
rect 33390 1450 33514 1492
rect 33558 1450 33682 1492
rect 48510 1532 48634 1574
rect 48678 1532 48802 1574
rect 48510 1492 48512 1532
rect 48512 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48634 1532
rect 48678 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48800 1532
rect 48800 1492 48802 1532
rect 48510 1450 48634 1492
rect 48678 1450 48802 1492
rect 63630 1532 63754 1574
rect 63798 1532 63922 1574
rect 63630 1492 63632 1532
rect 63632 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63754 1532
rect 63798 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63920 1532
rect 63920 1492 63922 1532
rect 63630 1450 63754 1492
rect 63798 1450 63922 1492
rect 78750 1532 78874 1574
rect 78918 1532 79042 1574
rect 78750 1492 78752 1532
rect 78752 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78874 1532
rect 78918 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79040 1532
rect 79040 1492 79042 1532
rect 78750 1450 78874 1492
rect 78918 1450 79042 1492
rect 4390 776 4514 818
rect 4558 776 4682 818
rect 4390 736 4392 776
rect 4392 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4514 776
rect 4558 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4680 776
rect 4680 736 4682 776
rect 4390 694 4514 736
rect 4558 694 4682 736
rect 19510 776 19634 818
rect 19678 776 19802 818
rect 19510 736 19512 776
rect 19512 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19634 776
rect 19678 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19800 776
rect 19800 736 19802 776
rect 19510 694 19634 736
rect 19678 694 19802 736
rect 34630 776 34754 818
rect 34798 776 34922 818
rect 34630 736 34632 776
rect 34632 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34754 776
rect 34798 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34920 776
rect 34920 736 34922 776
rect 34630 694 34754 736
rect 34798 694 34922 736
rect 49750 776 49874 818
rect 49918 776 50042 818
rect 49750 736 49752 776
rect 49752 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49874 776
rect 49918 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50040 776
rect 50040 736 50042 776
rect 49750 694 49874 736
rect 49918 694 50042 736
rect 64870 776 64994 818
rect 65038 776 65162 818
rect 64870 736 64872 776
rect 64872 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64994 776
rect 65038 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65160 776
rect 65160 736 65162 776
rect 64870 694 64994 736
rect 65038 694 65162 736
rect 79990 776 80114 818
rect 80158 776 80282 818
rect 79990 736 79992 776
rect 79992 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80114 776
rect 80158 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80280 776
rect 80280 736 80282 776
rect 79990 694 80114 736
rect 80158 694 80282 736
<< metal6 >>
rect 4316 38618 4756 38682
rect 3076 37862 3516 38600
rect 3076 37738 3150 37862
rect 3274 37738 3318 37862
rect 3442 37738 3516 37862
rect 3076 36350 3516 37738
rect 3076 36226 3150 36350
rect 3274 36226 3318 36350
rect 3442 36226 3516 36350
rect 3076 34838 3516 36226
rect 3076 34714 3150 34838
rect 3274 34714 3318 34838
rect 3442 34714 3516 34838
rect 3076 33326 3516 34714
rect 3076 33202 3150 33326
rect 3274 33202 3318 33326
rect 3442 33202 3516 33326
rect 3076 31814 3516 33202
rect 3076 31690 3150 31814
rect 3274 31690 3318 31814
rect 3442 31690 3516 31814
rect 3076 30302 3516 31690
rect 3076 30178 3150 30302
rect 3274 30178 3318 30302
rect 3442 30178 3516 30302
rect 3076 28790 3516 30178
rect 3076 28666 3150 28790
rect 3274 28666 3318 28790
rect 3442 28666 3516 28790
rect 3076 27278 3516 28666
rect 3076 27154 3150 27278
rect 3274 27154 3318 27278
rect 3442 27154 3516 27278
rect 3076 25766 3516 27154
rect 3076 25642 3150 25766
rect 3274 25642 3318 25766
rect 3442 25642 3516 25766
rect 3076 24254 3516 25642
rect 3076 24130 3150 24254
rect 3274 24130 3318 24254
rect 3442 24130 3516 24254
rect 3076 22742 3516 24130
rect 3076 22618 3150 22742
rect 3274 22618 3318 22742
rect 3442 22618 3516 22742
rect 3076 21230 3516 22618
rect 3076 21106 3150 21230
rect 3274 21106 3318 21230
rect 3442 21106 3516 21230
rect 3076 19718 3516 21106
rect 3076 19594 3150 19718
rect 3274 19594 3318 19718
rect 3442 19594 3516 19718
rect 3076 18206 3516 19594
rect 3076 18082 3150 18206
rect 3274 18082 3318 18206
rect 3442 18082 3516 18206
rect 3076 16694 3516 18082
rect 3076 16570 3150 16694
rect 3274 16570 3318 16694
rect 3442 16570 3516 16694
rect 3076 15182 3516 16570
rect 3076 15058 3150 15182
rect 3274 15058 3318 15182
rect 3442 15058 3516 15182
rect 3076 13670 3516 15058
rect 3076 13546 3150 13670
rect 3274 13546 3318 13670
rect 3442 13546 3516 13670
rect 3076 12158 3516 13546
rect 3076 12034 3150 12158
rect 3274 12034 3318 12158
rect 3442 12034 3516 12158
rect 3076 10646 3516 12034
rect 3076 10522 3150 10646
rect 3274 10522 3318 10646
rect 3442 10522 3516 10646
rect 3076 9134 3516 10522
rect 3076 9010 3150 9134
rect 3274 9010 3318 9134
rect 3442 9010 3516 9134
rect 3076 7622 3516 9010
rect 3076 7498 3150 7622
rect 3274 7498 3318 7622
rect 3442 7498 3516 7622
rect 3076 6110 3516 7498
rect 3076 5986 3150 6110
rect 3274 5986 3318 6110
rect 3442 5986 3516 6110
rect 3076 4598 3516 5986
rect 3076 4474 3150 4598
rect 3274 4474 3318 4598
rect 3442 4474 3516 4598
rect 3076 3086 3516 4474
rect 3076 2962 3150 3086
rect 3274 2962 3318 3086
rect 3442 2962 3516 3086
rect 3076 1574 3516 2962
rect 3076 1450 3150 1574
rect 3274 1450 3318 1574
rect 3442 1450 3516 1574
rect 3076 712 3516 1450
rect 4316 38494 4390 38618
rect 4514 38494 4558 38618
rect 4682 38494 4756 38618
rect 19436 38618 19876 38682
rect 4316 37106 4756 38494
rect 4316 36982 4390 37106
rect 4514 36982 4558 37106
rect 4682 36982 4756 37106
rect 4316 35594 4756 36982
rect 4316 35470 4390 35594
rect 4514 35470 4558 35594
rect 4682 35470 4756 35594
rect 4316 34082 4756 35470
rect 4316 33958 4390 34082
rect 4514 33958 4558 34082
rect 4682 33958 4756 34082
rect 4316 32570 4756 33958
rect 4316 32446 4390 32570
rect 4514 32446 4558 32570
rect 4682 32446 4756 32570
rect 4316 31058 4756 32446
rect 4316 30934 4390 31058
rect 4514 30934 4558 31058
rect 4682 30934 4756 31058
rect 4316 29546 4756 30934
rect 4316 29422 4390 29546
rect 4514 29422 4558 29546
rect 4682 29422 4756 29546
rect 4316 28034 4756 29422
rect 4316 27910 4390 28034
rect 4514 27910 4558 28034
rect 4682 27910 4756 28034
rect 4316 26522 4756 27910
rect 4316 26398 4390 26522
rect 4514 26398 4558 26522
rect 4682 26398 4756 26522
rect 4316 25010 4756 26398
rect 4316 24886 4390 25010
rect 4514 24886 4558 25010
rect 4682 24886 4756 25010
rect 4316 23498 4756 24886
rect 4316 23374 4390 23498
rect 4514 23374 4558 23498
rect 4682 23374 4756 23498
rect 4316 21986 4756 23374
rect 4316 21862 4390 21986
rect 4514 21862 4558 21986
rect 4682 21862 4756 21986
rect 4316 20474 4756 21862
rect 4316 20350 4390 20474
rect 4514 20350 4558 20474
rect 4682 20350 4756 20474
rect 4316 18962 4756 20350
rect 4316 18838 4390 18962
rect 4514 18838 4558 18962
rect 4682 18838 4756 18962
rect 4316 17450 4756 18838
rect 4316 17326 4390 17450
rect 4514 17326 4558 17450
rect 4682 17326 4756 17450
rect 4316 15938 4756 17326
rect 4316 15814 4390 15938
rect 4514 15814 4558 15938
rect 4682 15814 4756 15938
rect 4316 14426 4756 15814
rect 4316 14302 4390 14426
rect 4514 14302 4558 14426
rect 4682 14302 4756 14426
rect 4316 12914 4756 14302
rect 4316 12790 4390 12914
rect 4514 12790 4558 12914
rect 4682 12790 4756 12914
rect 4316 11402 4756 12790
rect 4316 11278 4390 11402
rect 4514 11278 4558 11402
rect 4682 11278 4756 11402
rect 4316 9890 4756 11278
rect 4316 9766 4390 9890
rect 4514 9766 4558 9890
rect 4682 9766 4756 9890
rect 4316 8378 4756 9766
rect 4316 8254 4390 8378
rect 4514 8254 4558 8378
rect 4682 8254 4756 8378
rect 4316 6866 4756 8254
rect 4316 6742 4390 6866
rect 4514 6742 4558 6866
rect 4682 6742 4756 6866
rect 4316 5354 4756 6742
rect 4316 5230 4390 5354
rect 4514 5230 4558 5354
rect 4682 5230 4756 5354
rect 4316 3842 4756 5230
rect 4316 3718 4390 3842
rect 4514 3718 4558 3842
rect 4682 3718 4756 3842
rect 4316 2330 4756 3718
rect 4316 2206 4390 2330
rect 4514 2206 4558 2330
rect 4682 2206 4756 2330
rect 4316 818 4756 2206
rect 4316 694 4390 818
rect 4514 694 4558 818
rect 4682 694 4756 818
rect 18196 37862 18636 38600
rect 18196 37738 18270 37862
rect 18394 37738 18438 37862
rect 18562 37738 18636 37862
rect 18196 36350 18636 37738
rect 18196 36226 18270 36350
rect 18394 36226 18438 36350
rect 18562 36226 18636 36350
rect 18196 34838 18636 36226
rect 18196 34714 18270 34838
rect 18394 34714 18438 34838
rect 18562 34714 18636 34838
rect 18196 29022 18636 34714
rect 18196 28898 18270 29022
rect 18394 28898 18438 29022
rect 18562 28898 18636 29022
rect 18196 28854 18636 28898
rect 18196 28730 18270 28854
rect 18394 28730 18438 28854
rect 18562 28730 18636 28854
rect 18196 23022 18636 28730
rect 18196 22898 18270 23022
rect 18394 22898 18438 23022
rect 18562 22898 18636 23022
rect 18196 22854 18636 22898
rect 18196 22730 18270 22854
rect 18394 22730 18438 22854
rect 18562 22730 18636 22854
rect 18196 17022 18636 22730
rect 18196 16898 18270 17022
rect 18394 16898 18438 17022
rect 18562 16898 18636 17022
rect 18196 16854 18636 16898
rect 18196 16730 18270 16854
rect 18394 16730 18438 16854
rect 18562 16730 18636 16854
rect 18196 11022 18636 16730
rect 18196 10898 18270 11022
rect 18394 10898 18438 11022
rect 18562 10898 18636 11022
rect 18196 10854 18636 10898
rect 18196 10730 18270 10854
rect 18394 10730 18438 10854
rect 18562 10730 18636 10854
rect 18196 4598 18636 10730
rect 18196 4474 18270 4598
rect 18394 4474 18438 4598
rect 18562 4474 18636 4598
rect 18196 3086 18636 4474
rect 18196 2962 18270 3086
rect 18394 2962 18438 3086
rect 18562 2962 18636 3086
rect 18196 1574 18636 2962
rect 18196 1450 18270 1574
rect 18394 1450 18438 1574
rect 18562 1450 18636 1574
rect 18196 712 18636 1450
rect 19436 38494 19510 38618
rect 19634 38494 19678 38618
rect 19802 38494 19876 38618
rect 34556 38618 34996 38682
rect 19436 37106 19876 38494
rect 19436 36982 19510 37106
rect 19634 36982 19678 37106
rect 19802 36982 19876 37106
rect 19436 35594 19876 36982
rect 19436 35470 19510 35594
rect 19634 35470 19678 35594
rect 19802 35470 19876 35594
rect 19436 34082 19876 35470
rect 19436 33958 19510 34082
rect 19634 33958 19678 34082
rect 19802 33958 19876 34082
rect 19436 24262 19876 33958
rect 19436 24138 19510 24262
rect 19634 24138 19678 24262
rect 19802 24138 19876 24262
rect 19436 24094 19876 24138
rect 19436 23970 19510 24094
rect 19634 23970 19678 24094
rect 19802 23970 19876 24094
rect 19436 18262 19876 23970
rect 19436 18138 19510 18262
rect 19634 18138 19678 18262
rect 19802 18138 19876 18262
rect 19436 18094 19876 18138
rect 19436 17970 19510 18094
rect 19634 17970 19678 18094
rect 19802 17970 19876 18094
rect 19436 12262 19876 17970
rect 19436 12138 19510 12262
rect 19634 12138 19678 12262
rect 19802 12138 19876 12262
rect 19436 12094 19876 12138
rect 19436 11970 19510 12094
rect 19634 11970 19678 12094
rect 19802 11970 19876 12094
rect 19436 5354 19876 11970
rect 19436 5230 19510 5354
rect 19634 5230 19678 5354
rect 19802 5230 19876 5354
rect 19436 3842 19876 5230
rect 19436 3718 19510 3842
rect 19634 3718 19678 3842
rect 19802 3718 19876 3842
rect 19436 2330 19876 3718
rect 19436 2206 19510 2330
rect 19634 2206 19678 2330
rect 19802 2206 19876 2330
rect 19436 818 19876 2206
rect 4316 630 4756 694
rect 19436 694 19510 818
rect 19634 694 19678 818
rect 19802 694 19876 818
rect 33316 37862 33756 38600
rect 33316 37738 33390 37862
rect 33514 37738 33558 37862
rect 33682 37738 33756 37862
rect 33316 36350 33756 37738
rect 33316 36226 33390 36350
rect 33514 36226 33558 36350
rect 33682 36226 33756 36350
rect 33316 34838 33756 36226
rect 33316 34714 33390 34838
rect 33514 34714 33558 34838
rect 33682 34714 33756 34838
rect 33316 29022 33756 34714
rect 33316 28898 33390 29022
rect 33514 28898 33558 29022
rect 33682 28898 33756 29022
rect 33316 28854 33756 28898
rect 33316 28730 33390 28854
rect 33514 28730 33558 28854
rect 33682 28730 33756 28854
rect 33316 23022 33756 28730
rect 33316 22898 33390 23022
rect 33514 22898 33558 23022
rect 33682 22898 33756 23022
rect 33316 22854 33756 22898
rect 33316 22730 33390 22854
rect 33514 22730 33558 22854
rect 33682 22730 33756 22854
rect 33316 17022 33756 22730
rect 33316 16898 33390 17022
rect 33514 16898 33558 17022
rect 33682 16898 33756 17022
rect 33316 16854 33756 16898
rect 33316 16730 33390 16854
rect 33514 16730 33558 16854
rect 33682 16730 33756 16854
rect 33316 11022 33756 16730
rect 33316 10898 33390 11022
rect 33514 10898 33558 11022
rect 33682 10898 33756 11022
rect 33316 10854 33756 10898
rect 33316 10730 33390 10854
rect 33514 10730 33558 10854
rect 33682 10730 33756 10854
rect 33316 4598 33756 10730
rect 33316 4474 33390 4598
rect 33514 4474 33558 4598
rect 33682 4474 33756 4598
rect 33316 3086 33756 4474
rect 33316 2962 33390 3086
rect 33514 2962 33558 3086
rect 33682 2962 33756 3086
rect 33316 1574 33756 2962
rect 33316 1450 33390 1574
rect 33514 1450 33558 1574
rect 33682 1450 33756 1574
rect 33316 712 33756 1450
rect 34556 38494 34630 38618
rect 34754 38494 34798 38618
rect 34922 38494 34996 38618
rect 49676 38618 50116 38682
rect 34556 37106 34996 38494
rect 34556 36982 34630 37106
rect 34754 36982 34798 37106
rect 34922 36982 34996 37106
rect 34556 35594 34996 36982
rect 34556 35470 34630 35594
rect 34754 35470 34798 35594
rect 34922 35470 34996 35594
rect 34556 34082 34996 35470
rect 34556 33958 34630 34082
rect 34754 33958 34798 34082
rect 34922 33958 34996 34082
rect 34556 24262 34996 33958
rect 34556 24138 34630 24262
rect 34754 24138 34798 24262
rect 34922 24138 34996 24262
rect 34556 24094 34996 24138
rect 34556 23970 34630 24094
rect 34754 23970 34798 24094
rect 34922 23970 34996 24094
rect 34556 18262 34996 23970
rect 34556 18138 34630 18262
rect 34754 18138 34798 18262
rect 34922 18138 34996 18262
rect 34556 18094 34996 18138
rect 34556 17970 34630 18094
rect 34754 17970 34798 18094
rect 34922 17970 34996 18094
rect 34556 12262 34996 17970
rect 34556 12138 34630 12262
rect 34754 12138 34798 12262
rect 34922 12138 34996 12262
rect 34556 12094 34996 12138
rect 34556 11970 34630 12094
rect 34754 11970 34798 12094
rect 34922 11970 34996 12094
rect 34556 5354 34996 11970
rect 34556 5230 34630 5354
rect 34754 5230 34798 5354
rect 34922 5230 34996 5354
rect 34556 3842 34996 5230
rect 34556 3718 34630 3842
rect 34754 3718 34798 3842
rect 34922 3718 34996 3842
rect 34556 2330 34996 3718
rect 34556 2206 34630 2330
rect 34754 2206 34798 2330
rect 34922 2206 34996 2330
rect 34556 818 34996 2206
rect 19436 630 19876 694
rect 34556 694 34630 818
rect 34754 694 34798 818
rect 34922 694 34996 818
rect 48436 37862 48876 38600
rect 48436 37738 48510 37862
rect 48634 37738 48678 37862
rect 48802 37738 48876 37862
rect 48436 36350 48876 37738
rect 48436 36226 48510 36350
rect 48634 36226 48678 36350
rect 48802 36226 48876 36350
rect 48436 34838 48876 36226
rect 48436 34714 48510 34838
rect 48634 34714 48678 34838
rect 48802 34714 48876 34838
rect 48436 29022 48876 34714
rect 48436 28898 48510 29022
rect 48634 28898 48678 29022
rect 48802 28898 48876 29022
rect 48436 28854 48876 28898
rect 48436 28730 48510 28854
rect 48634 28730 48678 28854
rect 48802 28730 48876 28854
rect 48436 23022 48876 28730
rect 48436 22898 48510 23022
rect 48634 22898 48678 23022
rect 48802 22898 48876 23022
rect 48436 22854 48876 22898
rect 48436 22730 48510 22854
rect 48634 22730 48678 22854
rect 48802 22730 48876 22854
rect 48436 17022 48876 22730
rect 48436 16898 48510 17022
rect 48634 16898 48678 17022
rect 48802 16898 48876 17022
rect 48436 16854 48876 16898
rect 48436 16730 48510 16854
rect 48634 16730 48678 16854
rect 48802 16730 48876 16854
rect 48436 11022 48876 16730
rect 48436 10898 48510 11022
rect 48634 10898 48678 11022
rect 48802 10898 48876 11022
rect 48436 10854 48876 10898
rect 48436 10730 48510 10854
rect 48634 10730 48678 10854
rect 48802 10730 48876 10854
rect 48436 4598 48876 10730
rect 48436 4474 48510 4598
rect 48634 4474 48678 4598
rect 48802 4474 48876 4598
rect 48436 3086 48876 4474
rect 48436 2962 48510 3086
rect 48634 2962 48678 3086
rect 48802 2962 48876 3086
rect 48436 1574 48876 2962
rect 48436 1450 48510 1574
rect 48634 1450 48678 1574
rect 48802 1450 48876 1574
rect 48436 712 48876 1450
rect 49676 38494 49750 38618
rect 49874 38494 49918 38618
rect 50042 38494 50116 38618
rect 64796 38618 65236 38682
rect 49676 37106 50116 38494
rect 49676 36982 49750 37106
rect 49874 36982 49918 37106
rect 50042 36982 50116 37106
rect 49676 35594 50116 36982
rect 49676 35470 49750 35594
rect 49874 35470 49918 35594
rect 50042 35470 50116 35594
rect 49676 34082 50116 35470
rect 49676 33958 49750 34082
rect 49874 33958 49918 34082
rect 50042 33958 50116 34082
rect 49676 24262 50116 33958
rect 49676 24138 49750 24262
rect 49874 24138 49918 24262
rect 50042 24138 50116 24262
rect 49676 24094 50116 24138
rect 49676 23970 49750 24094
rect 49874 23970 49918 24094
rect 50042 23970 50116 24094
rect 49676 18262 50116 23970
rect 49676 18138 49750 18262
rect 49874 18138 49918 18262
rect 50042 18138 50116 18262
rect 49676 18094 50116 18138
rect 49676 17970 49750 18094
rect 49874 17970 49918 18094
rect 50042 17970 50116 18094
rect 49676 12262 50116 17970
rect 49676 12138 49750 12262
rect 49874 12138 49918 12262
rect 50042 12138 50116 12262
rect 49676 12094 50116 12138
rect 49676 11970 49750 12094
rect 49874 11970 49918 12094
rect 50042 11970 50116 12094
rect 49676 5354 50116 11970
rect 49676 5230 49750 5354
rect 49874 5230 49918 5354
rect 50042 5230 50116 5354
rect 49676 3842 50116 5230
rect 49676 3718 49750 3842
rect 49874 3718 49918 3842
rect 50042 3718 50116 3842
rect 49676 2330 50116 3718
rect 49676 2206 49750 2330
rect 49874 2206 49918 2330
rect 50042 2206 50116 2330
rect 49676 818 50116 2206
rect 34556 630 34996 694
rect 49676 694 49750 818
rect 49874 694 49918 818
rect 50042 694 50116 818
rect 63556 37862 63996 38600
rect 63556 37738 63630 37862
rect 63754 37738 63798 37862
rect 63922 37738 63996 37862
rect 63556 36350 63996 37738
rect 63556 36226 63630 36350
rect 63754 36226 63798 36350
rect 63922 36226 63996 36350
rect 63556 34838 63996 36226
rect 63556 34714 63630 34838
rect 63754 34714 63798 34838
rect 63922 34714 63996 34838
rect 63556 29022 63996 34714
rect 63556 28898 63630 29022
rect 63754 28898 63798 29022
rect 63922 28898 63996 29022
rect 63556 28854 63996 28898
rect 63556 28730 63630 28854
rect 63754 28730 63798 28854
rect 63922 28730 63996 28854
rect 63556 23022 63996 28730
rect 63556 22898 63630 23022
rect 63754 22898 63798 23022
rect 63922 22898 63996 23022
rect 63556 22854 63996 22898
rect 63556 22730 63630 22854
rect 63754 22730 63798 22854
rect 63922 22730 63996 22854
rect 63556 17022 63996 22730
rect 63556 16898 63630 17022
rect 63754 16898 63798 17022
rect 63922 16898 63996 17022
rect 63556 16854 63996 16898
rect 63556 16730 63630 16854
rect 63754 16730 63798 16854
rect 63922 16730 63996 16854
rect 63556 11022 63996 16730
rect 63556 10898 63630 11022
rect 63754 10898 63798 11022
rect 63922 10898 63996 11022
rect 63556 10854 63996 10898
rect 63556 10730 63630 10854
rect 63754 10730 63798 10854
rect 63922 10730 63996 10854
rect 63556 4598 63996 10730
rect 63556 4474 63630 4598
rect 63754 4474 63798 4598
rect 63922 4474 63996 4598
rect 63556 3086 63996 4474
rect 63556 2962 63630 3086
rect 63754 2962 63798 3086
rect 63922 2962 63996 3086
rect 63556 1574 63996 2962
rect 63556 1450 63630 1574
rect 63754 1450 63798 1574
rect 63922 1450 63996 1574
rect 63556 712 63996 1450
rect 64796 38494 64870 38618
rect 64994 38494 65038 38618
rect 65162 38494 65236 38618
rect 79916 38618 80356 38682
rect 64796 37106 65236 38494
rect 64796 36982 64870 37106
rect 64994 36982 65038 37106
rect 65162 36982 65236 37106
rect 64796 35594 65236 36982
rect 64796 35470 64870 35594
rect 64994 35470 65038 35594
rect 65162 35470 65236 35594
rect 64796 34082 65236 35470
rect 64796 33958 64870 34082
rect 64994 33958 65038 34082
rect 65162 33958 65236 34082
rect 78676 37862 79116 38600
rect 78676 37738 78750 37862
rect 78874 37738 78918 37862
rect 79042 37738 79116 37862
rect 78676 36350 79116 37738
rect 78676 36226 78750 36350
rect 78874 36226 78918 36350
rect 79042 36226 79116 36350
rect 78676 34838 79116 36226
rect 78676 34714 78750 34838
rect 78874 34714 78918 34838
rect 79042 34714 79116 34838
rect 64796 24262 65236 33958
rect 67196 33914 67524 34016
rect 67196 33790 67298 33914
rect 67422 33790 67524 33914
rect 64796 24138 64870 24262
rect 64994 24138 65038 24262
rect 65162 24138 65236 24262
rect 64796 24094 65236 24138
rect 64796 23970 64870 24094
rect 64994 23970 65038 24094
rect 65162 23970 65236 24094
rect 64796 18262 65236 23970
rect 64796 18138 64870 18262
rect 64994 18138 65038 18262
rect 65162 18138 65236 18262
rect 64796 18094 65236 18138
rect 64796 17970 64870 18094
rect 64994 17970 65038 18094
rect 65162 17970 65236 18094
rect 64796 12262 65236 17970
rect 64796 12138 64870 12262
rect 64994 12138 65038 12262
rect 65162 12138 65236 12262
rect 64796 12094 65236 12138
rect 64796 11970 64870 12094
rect 64994 11970 65038 12094
rect 65162 11970 65236 12094
rect 64796 5354 65236 11970
rect 64796 5230 64870 5354
rect 64994 5230 65038 5354
rect 65162 5230 65236 5354
rect 64796 3842 65236 5230
rect 66284 30050 66612 30152
rect 66284 29926 66386 30050
rect 66510 29926 66612 30050
rect 66284 4766 66612 29926
rect 67196 5774 67524 33790
rect 67196 5650 67298 5774
rect 67422 5650 67524 5774
rect 67196 5548 67524 5650
rect 78676 33326 79116 34714
rect 78676 33202 78750 33326
rect 78874 33202 78918 33326
rect 79042 33202 79116 33326
rect 78676 31814 79116 33202
rect 78676 31690 78750 31814
rect 78874 31690 78918 31814
rect 79042 31690 79116 31814
rect 78676 30302 79116 31690
rect 78676 30178 78750 30302
rect 78874 30178 78918 30302
rect 79042 30178 79116 30302
rect 78676 28790 79116 30178
rect 78676 28666 78750 28790
rect 78874 28666 78918 28790
rect 79042 28666 79116 28790
rect 78676 27278 79116 28666
rect 78676 27154 78750 27278
rect 78874 27154 78918 27278
rect 79042 27154 79116 27278
rect 78676 25766 79116 27154
rect 78676 25642 78750 25766
rect 78874 25642 78918 25766
rect 79042 25642 79116 25766
rect 78676 24254 79116 25642
rect 78676 24130 78750 24254
rect 78874 24130 78918 24254
rect 79042 24130 79116 24254
rect 78676 22742 79116 24130
rect 78676 22618 78750 22742
rect 78874 22618 78918 22742
rect 79042 22618 79116 22742
rect 78676 21230 79116 22618
rect 78676 21106 78750 21230
rect 78874 21106 78918 21230
rect 79042 21106 79116 21230
rect 78676 19718 79116 21106
rect 78676 19594 78750 19718
rect 78874 19594 78918 19718
rect 79042 19594 79116 19718
rect 78676 18206 79116 19594
rect 78676 18082 78750 18206
rect 78874 18082 78918 18206
rect 79042 18082 79116 18206
rect 78676 16694 79116 18082
rect 78676 16570 78750 16694
rect 78874 16570 78918 16694
rect 79042 16570 79116 16694
rect 78676 15182 79116 16570
rect 78676 15058 78750 15182
rect 78874 15058 78918 15182
rect 79042 15058 79116 15182
rect 78676 13670 79116 15058
rect 78676 13546 78750 13670
rect 78874 13546 78918 13670
rect 79042 13546 79116 13670
rect 78676 12158 79116 13546
rect 78676 12034 78750 12158
rect 78874 12034 78918 12158
rect 79042 12034 79116 12158
rect 78676 10646 79116 12034
rect 78676 10522 78750 10646
rect 78874 10522 78918 10646
rect 79042 10522 79116 10646
rect 78676 9134 79116 10522
rect 78676 9010 78750 9134
rect 78874 9010 78918 9134
rect 79042 9010 79116 9134
rect 78676 7622 79116 9010
rect 78676 7498 78750 7622
rect 78874 7498 78918 7622
rect 79042 7498 79116 7622
rect 78676 6110 79116 7498
rect 78676 5986 78750 6110
rect 78874 5986 78918 6110
rect 79042 5986 79116 6110
rect 66284 4642 66386 4766
rect 66510 4642 66612 4766
rect 66284 4540 66612 4642
rect 78676 4598 79116 5986
rect 64796 3718 64870 3842
rect 64994 3718 65038 3842
rect 65162 3718 65236 3842
rect 64796 2330 65236 3718
rect 64796 2206 64870 2330
rect 64994 2206 65038 2330
rect 65162 2206 65236 2330
rect 64796 818 65236 2206
rect 49676 630 50116 694
rect 64796 694 64870 818
rect 64994 694 65038 818
rect 65162 694 65236 818
rect 78676 4474 78750 4598
rect 78874 4474 78918 4598
rect 79042 4474 79116 4598
rect 78676 3086 79116 4474
rect 78676 2962 78750 3086
rect 78874 2962 78918 3086
rect 79042 2962 79116 3086
rect 78676 1574 79116 2962
rect 78676 1450 78750 1574
rect 78874 1450 78918 1574
rect 79042 1450 79116 1574
rect 78676 712 79116 1450
rect 79916 38494 79990 38618
rect 80114 38494 80158 38618
rect 80282 38494 80356 38618
rect 79916 37106 80356 38494
rect 79916 36982 79990 37106
rect 80114 36982 80158 37106
rect 80282 36982 80356 37106
rect 79916 35594 80356 36982
rect 79916 35470 79990 35594
rect 80114 35470 80158 35594
rect 80282 35470 80356 35594
rect 79916 34082 80356 35470
rect 79916 33958 79990 34082
rect 80114 33958 80158 34082
rect 80282 33958 80356 34082
rect 79916 32570 80356 33958
rect 79916 32446 79990 32570
rect 80114 32446 80158 32570
rect 80282 32446 80356 32570
rect 79916 31058 80356 32446
rect 79916 30934 79990 31058
rect 80114 30934 80158 31058
rect 80282 30934 80356 31058
rect 79916 29546 80356 30934
rect 79916 29422 79990 29546
rect 80114 29422 80158 29546
rect 80282 29422 80356 29546
rect 79916 28034 80356 29422
rect 79916 27910 79990 28034
rect 80114 27910 80158 28034
rect 80282 27910 80356 28034
rect 79916 26522 80356 27910
rect 79916 26398 79990 26522
rect 80114 26398 80158 26522
rect 80282 26398 80356 26522
rect 79916 25010 80356 26398
rect 79916 24886 79990 25010
rect 80114 24886 80158 25010
rect 80282 24886 80356 25010
rect 79916 23498 80356 24886
rect 79916 23374 79990 23498
rect 80114 23374 80158 23498
rect 80282 23374 80356 23498
rect 79916 21986 80356 23374
rect 79916 21862 79990 21986
rect 80114 21862 80158 21986
rect 80282 21862 80356 21986
rect 79916 20474 80356 21862
rect 79916 20350 79990 20474
rect 80114 20350 80158 20474
rect 80282 20350 80356 20474
rect 79916 18962 80356 20350
rect 79916 18838 79990 18962
rect 80114 18838 80158 18962
rect 80282 18838 80356 18962
rect 79916 17450 80356 18838
rect 79916 17326 79990 17450
rect 80114 17326 80158 17450
rect 80282 17326 80356 17450
rect 79916 15938 80356 17326
rect 79916 15814 79990 15938
rect 80114 15814 80158 15938
rect 80282 15814 80356 15938
rect 79916 14426 80356 15814
rect 79916 14302 79990 14426
rect 80114 14302 80158 14426
rect 80282 14302 80356 14426
rect 79916 12914 80356 14302
rect 79916 12790 79990 12914
rect 80114 12790 80158 12914
rect 80282 12790 80356 12914
rect 79916 11402 80356 12790
rect 79916 11278 79990 11402
rect 80114 11278 80158 11402
rect 80282 11278 80356 11402
rect 79916 9890 80356 11278
rect 79916 9766 79990 9890
rect 80114 9766 80158 9890
rect 80282 9766 80356 9890
rect 79916 8378 80356 9766
rect 79916 8254 79990 8378
rect 80114 8254 80158 8378
rect 80282 8254 80356 8378
rect 79916 6866 80356 8254
rect 79916 6742 79990 6866
rect 80114 6742 80158 6866
rect 80282 6742 80356 6866
rect 79916 5354 80356 6742
rect 79916 5230 79990 5354
rect 80114 5230 80158 5354
rect 80282 5230 80356 5354
rect 79916 3842 80356 5230
rect 79916 3718 79990 3842
rect 80114 3718 80158 3842
rect 80282 3718 80356 3842
rect 79916 2330 80356 3718
rect 79916 2206 79990 2330
rect 80114 2206 80158 2330
rect 80282 2206 80356 2330
rect 79916 818 80356 2206
rect 64796 630 65236 694
rect 79916 694 79990 818
rect 80114 694 80158 818
rect 80282 694 80356 818
rect 93796 34222 94236 38600
rect 93796 34098 93870 34222
rect 93994 34098 94038 34222
rect 94162 34098 94236 34222
rect 93796 34054 94236 34098
rect 93796 33930 93870 34054
rect 93994 33930 94038 34054
rect 94162 33930 94236 34054
rect 93796 28222 94236 33930
rect 93796 28098 93870 28222
rect 93994 28098 94038 28222
rect 94162 28098 94236 28222
rect 93796 28054 94236 28098
rect 93796 27930 93870 28054
rect 93994 27930 94038 28054
rect 94162 27930 94236 28054
rect 93796 21230 94236 27930
rect 93796 21106 93870 21230
rect 93994 21106 94038 21230
rect 94162 21106 94236 21230
rect 93796 19718 94236 21106
rect 93796 19594 93870 19718
rect 93994 19594 94038 19718
rect 94162 19594 94236 19718
rect 93796 11022 94236 19594
rect 93796 10898 93870 11022
rect 93994 10898 94038 11022
rect 94162 10898 94236 11022
rect 93796 10854 94236 10898
rect 93796 10730 93870 10854
rect 93994 10730 94038 10854
rect 94162 10730 94236 10854
rect 93796 5022 94236 10730
rect 93796 4898 93870 5022
rect 93994 4898 94038 5022
rect 94162 4898 94236 5022
rect 93796 4854 94236 4898
rect 93796 4730 93870 4854
rect 93994 4730 94038 4854
rect 94162 4730 94236 4854
rect 93796 712 94236 4730
rect 95036 29462 95476 38600
rect 95036 29338 95110 29462
rect 95234 29338 95278 29462
rect 95402 29338 95476 29462
rect 95036 29294 95476 29338
rect 95036 29170 95110 29294
rect 95234 29170 95278 29294
rect 95402 29170 95476 29294
rect 95036 21986 95476 29170
rect 95036 21862 95110 21986
rect 95234 21862 95278 21986
rect 95402 21862 95476 21986
rect 95036 20474 95476 21862
rect 95036 20350 95110 20474
rect 95234 20350 95278 20474
rect 95402 20350 95476 20474
rect 95036 12262 95476 20350
rect 95036 12138 95110 12262
rect 95234 12138 95278 12262
rect 95402 12138 95476 12262
rect 95036 12094 95476 12138
rect 95036 11970 95110 12094
rect 95234 11970 95278 12094
rect 95402 11970 95476 12094
rect 95036 6262 95476 11970
rect 95036 6138 95110 6262
rect 95234 6138 95278 6262
rect 95402 6138 95476 6262
rect 95036 6094 95476 6138
rect 95036 5970 95110 6094
rect 95234 5970 95278 6094
rect 95402 5970 95476 6094
rect 95036 712 95476 5970
rect 79916 630 80356 694
use sg13g2_inv_1  _128_
timestamp 1676382929
transform 1 0 22848 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  _129_
timestamp 1676382929
transform 1 0 42144 0 1 34020
box -48 -56 336 834
use sg13g2_mux2_1  _130_
timestamp 1677247768
transform 1 0 39360 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _131_
timestamp 1677247768
transform 1 0 41664 0 1 35532
box -48 -56 1008 834
use sg13g2_nor2_1  _132_
timestamp 1676627187
transform 1 0 42240 0 1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _133_
timestamp 1683973020
transform 1 0 42912 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2b_1  _134_
timestamp 1685181386
transform 1 0 32160 0 -1 3780
box -54 -56 528 834
use sg13g2_and2_1  _135_
timestamp 1676901763
transform 1 0 32064 0 -1 5292
box -48 -56 528 834
use sg13g2_and2_1  _136_
timestamp 1676901763
transform 1 0 31584 0 1 2268
box -48 -56 528 834
use sg13g2_and2_1  _137_
timestamp 1676901763
transform 1 0 32064 0 1 2268
box -48 -56 528 834
use sg13g2_nor2_1  _138_
timestamp 1676627187
transform 1 0 41568 0 1 34020
box -48 -56 432 834
use sg13g2_and2_1  _139_
timestamp 1676901763
transform 1 0 34560 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _140_
timestamp 1685175443
transform 1 0 40896 0 -1 3780
box -48 -56 538 834
use sg13g2_nor2_1  _141_
timestamp 1676627187
transform 1 0 35040 0 1 3780
box -48 -56 432 834
use sg13g2_a22oi_1  _142_
timestamp 1685173987
transform 1 0 38208 0 -1 3780
box -48 -56 624 834
use sg13g2_o21ai_1  _143_
timestamp 1685175443
transform 1 0 40608 0 1 3780
box -48 -56 538 834
use sg13g2_nand2_1  _144_
timestamp 1676557249
transform 1 0 35616 0 1 756
box -48 -56 432 834
use sg13g2_a22oi_1  _145_
timestamp 1685173987
transform 1 0 34752 0 -1 3780
box -48 -56 624 834
use sg13g2_nand2_1  _146_
timestamp 1676557249
transform 1 0 34752 0 1 2268
box -48 -56 432 834
use sg13g2_nand2_1  _147_
timestamp 1676557249
transform 1 0 36864 0 -1 5292
box -48 -56 432 834
use sg13g2_a22oi_1  _148_
timestamp 1685173987
transform 1 0 36864 0 -1 3780
box -48 -56 624 834
use sg13g2_nand2_1  _149_
timestamp 1676557249
transform 1 0 36192 0 1 3780
box -48 -56 432 834
use sg13g2_nand2b_1  _150_
timestamp 1676567195
transform 1 0 39936 0 1 3780
box -48 -56 528 834
use sg13g2_a22oi_1  _151_
timestamp 1685173987
transform -1 0 39072 0 -1 5292
box -48 -56 624 834
use sg13g2_nand2_1  _152_
timestamp 1676557249
transform 1 0 39072 0 -1 5292
box -48 -56 432 834
use sg13g2_mux4_1  _153_
timestamp 1677257233
transform 1 0 42624 0 1 3780
box -48 -56 2064 834
use sg13g2_nor2b_1  _154_
timestamp 1685181386
transform 1 0 20352 0 -1 37044
box -54 -56 528 834
use sg13g2_nand2b_1  _155_
timestamp 1676567195
transform 1 0 19200 0 1 37044
box -48 -56 528 834
use sg13g2_and2_1  _156_
timestamp 1676901763
transform 1 0 24288 0 -1 37044
box -48 -56 528 834
use sg13g2_nor3_1  _157_
timestamp 1676639442
transform 1 0 27072 0 -1 37044
box -48 -56 528 834
use sg13g2_nand4_1  _158_
timestamp 1685201930
transform 1 0 26784 0 -1 38556
box -48 -56 624 834
use sg13g2_inv_1  _159_
timestamp 1676382929
transform 1 0 20832 0 -1 37044
box -48 -56 336 834
use sg13g2_nand3_1  _160_
timestamp 1683988354
transform 1 0 21504 0 1 35532
box -48 -56 528 834
use sg13g2_a21o_1  _161_
timestamp 1677175127
transform 1 0 21216 0 -1 37044
box -48 -56 720 834
use sg13g2_and2_1  _162_
timestamp 1676901763
transform 1 0 20928 0 -1 38556
box -48 -56 528 834
use sg13g2_nand3_1  _163_
timestamp 1683988354
transform 1 0 23136 0 -1 37044
box -48 -56 528 834
use sg13g2_xnor2_1  _164_
timestamp 1677516600
transform 1 0 21984 0 -1 37044
box -48 -56 816 834
use sg13g2_and3_1  _165_
timestamp 1676971669
transform 1 0 24960 0 -1 37044
box -48 -56 720 834
use sg13g2_a21oi_1  _166_
timestamp 1683973020
transform 1 0 23616 0 -1 37044
box -48 -56 528 834
use sg13g2_xor2_1  _167_
timestamp 1677577977
transform 1 0 26688 0 -1 35532
box -48 -56 816 834
use sg13g2_and2_1  _168_
timestamp 1676901763
transform 1 0 27552 0 -1 37044
box -48 -56 528 834
use sg13g2_and4_1  _169_
timestamp 1676985977
transform 1 0 26304 0 -1 37044
box -48 -56 816 834
use sg13g2_a21oi_1  _170_
timestamp 1683973020
transform 1 0 25824 0 -1 37044
box -48 -56 528 834
use sg13g2_nor2_1  _171_
timestamp 1676627187
transform 1 0 25824 0 1 37044
box -48 -56 432 834
use sg13g2_nand2_1  _172_
timestamp 1676557249
transform 1 0 29184 0 -1 38556
box -48 -56 432 834
use sg13g2_xor2_1  _173_
timestamp 1677577977
transform 1 0 28416 0 -1 38556
box -48 -56 816 834
use sg13g2_xnor2_1  _174_
timestamp 1677516600
transform 1 0 29088 0 1 37044
box -48 -56 816 834
use sg13g2_mux2_1  _175_
timestamp 1677247768
transform 1 0 23616 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _176_
timestamp 1677247768
transform 1 0 27840 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _177_
timestamp 1677247768
transform 1 0 28800 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _178_
timestamp 1677247768
transform 1 0 31392 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _179_
timestamp 1677247768
transform 1 0 34944 0 -1 37044
box -48 -56 1008 834
use sg13g2_mux2_1  _180_
timestamp 1677247768
transform 1 0 46560 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _181_
timestamp 1677247768
transform 1 0 49920 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _182_
timestamp 1677247768
transform 1 0 52128 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _183_
timestamp 1677247768
transform 1 0 53088 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _184_
timestamp 1677247768
transform 1 0 46368 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _185_
timestamp 1677247768
transform 1 0 38592 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _186_
timestamp 1677247768
transform 1 0 34656 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _187_
timestamp 1677247768
transform 1 0 31104 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _188_
timestamp 1677247768
transform 1 0 30144 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _189_
timestamp 1677247768
transform 1 0 30048 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _190_
timestamp 1677247768
transform 1 0 45696 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _191_
timestamp 1677247768
transform 1 0 46944 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _192_
timestamp 1677247768
transform 1 0 49632 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _193_
timestamp 1677247768
transform 1 0 51552 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _194_
timestamp 1677247768
transform 1 0 53184 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _195_
timestamp 1677247768
transform 1 0 48960 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _196_
timestamp 1677247768
transform 1 0 51264 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _197_
timestamp 1677247768
transform 1 0 42048 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _198_
timestamp 1677247768
transform 1 0 44256 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _199_
timestamp 1677247768
transform 1 0 33984 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _200_
timestamp 1677247768
transform 1 0 31392 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _201_
timestamp 1677247768
transform 1 0 29184 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _202_
timestamp 1677247768
transform 1 0 27648 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _203_
timestamp 1677247768
transform 1 0 26208 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _204_
timestamp 1677247768
transform 1 0 25536 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _205_
timestamp 1677247768
transform 1 0 23904 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _206_
timestamp 1677247768
transform 1 0 20064 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _207_
timestamp 1677247768
transform 1 0 21216 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _208_
timestamp 1677247768
transform 1 0 21600 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _209_
timestamp 1677247768
transform 1 0 22560 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _210_
timestamp 1677247768
transform 1 0 25632 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _211_
timestamp 1677247768
transform 1 0 39840 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _212_
timestamp 1677247768
transform 1 0 38496 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _213_
timestamp 1677247768
transform 1 0 36480 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _214_
timestamp 1677247768
transform 1 0 3840 0 1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  _215_
timestamp 1677247768
transform 1 0 1920 0 1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  _216_
timestamp 1677247768
transform 1 0 3552 0 1 21924
box -48 -56 1008 834
use sg13g2_mux2_1  _217_
timestamp 1677247768
transform 1 0 4224 0 -1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  _218_
timestamp 1677247768
transform 1 0 10752 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _219_
timestamp 1677247768
transform 1 0 13248 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _220_
timestamp 1677247768
transform 1 0 14016 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _221_
timestamp 1677247768
transform 1 0 4320 0 1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  _222_
timestamp 1677247768
transform 1 0 3840 0 -1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  _223_
timestamp 1677247768
transform 1 0 1536 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  _224_
timestamp 1677247768
transform 1 0 1344 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _225_
timestamp 1677247768
transform 1 0 1344 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _226_
timestamp 1677247768
transform 1 0 1344 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _227_
timestamp 1677247768
transform 1 0 672 0 1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  _228_
timestamp 1677247768
transform 1 0 1440 0 1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  _229_
timestamp 1677247768
transform 1 0 3744 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  _230_
timestamp 1677247768
transform 1 0 4320 0 -1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  _231_
timestamp 1677247768
transform 1 0 15456 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _232_
timestamp 1677247768
transform 1 0 19584 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _233_
timestamp 1677247768
transform 1 0 18144 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _234_
timestamp 1677247768
transform 1 0 16416 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _235_
timestamp 1677247768
transform 1 0 16800 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _236_
timestamp 1677247768
transform 1 0 4224 0 1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _237_
timestamp 1677247768
transform 1 0 3744 0 1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  _238_
timestamp 1677247768
transform 1 0 3456 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _239_
timestamp 1677247768
transform 1 0 4128 0 1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _240_
timestamp 1677247768
transform 1 0 4128 0 1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _241_
timestamp 1677247768
transform 1 0 77184 0 -1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  _242_
timestamp 1677247768
transform 1 0 81504 0 1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  _243_
timestamp 1677247768
transform 1 0 81120 0 -1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  _244_
timestamp 1677247768
transform 1 0 79776 0 1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  _245_
timestamp 1677247768
transform 1 0 80064 0 -1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  _246_
timestamp 1677247768
transform 1 0 79872 0 -1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  _247_
timestamp 1677247768
transform 1 0 79008 0 1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  _248_
timestamp 1677247768
transform 1 0 79200 0 1 27972
box -48 -56 1008 834
use sg13g2_mux2_1  _249_
timestamp 1677247768
transform 1 0 80832 0 -1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  _250_
timestamp 1677247768
transform 1 0 80544 0 1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  _251_
timestamp 1677247768
transform 1 0 80544 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _252_
timestamp 1677247768
transform 1 0 79584 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _253_
timestamp 1677247768
transform 1 0 43392 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _254_
timestamp 1677247768
transform 1 0 41088 0 1 37044
box -48 -56 1008 834
use sg13g2_mux2_1  _255_
timestamp 1677247768
transform 1 0 40896 0 -1 38556
box -48 -56 1008 834
use sg13g2_mux2_1  _256_
timestamp 1677247768
transform 1 0 38304 0 -1 38556
box -48 -56 1008 834
use sg13g2_mux2_1  _257_
timestamp 1677247768
transform 1 0 38304 0 1 35532
box -48 -56 1008 834
use sg13g2_nor2_1  _258_
timestamp 1676627187
transform 1 0 40320 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _259_
timestamp 1683973020
transform 1 0 40992 0 1 34020
box -48 -56 528 834
use sg13g2_nor2_1  _260_
timestamp 1676627187
transform 1 0 42624 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _261_
timestamp 1683973020
transform 1 0 43392 0 -1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _262_
timestamp 1677247768
transform 1 0 47616 0 -1 2268
box -48 -56 1008 834
use sg13g2_a21o_1  _263_
timestamp 1677175127
transform 1 0 18816 0 1 35532
box -48 -56 720 834
use sg13g2_dfrbpq_1  _264_
timestamp 1746535128
transform 1 0 20064 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _265_
timestamp 1746535128
transform 1 0 22656 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _266_
timestamp 1746535128
transform 1 0 22368 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _267_
timestamp 1746535128
transform 1 0 25536 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _268_
timestamp 1746535128
transform 1 0 26208 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _269_
timestamp 1746535128
transform 1 0 28992 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _270_
timestamp 1746535128
transform 1 0 29856 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _271_
timestamp 1746535128
transform 1 0 24576 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _272_
timestamp 1746535128
transform 1 0 27936 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _273_
timestamp 1746535128
transform 1 0 29760 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _274_
timestamp 1746535128
transform 1 0 32352 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _275_
timestamp 1746535128
transform 1 0 35328 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _276_
timestamp 1746535128
transform 1 0 47328 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _277_
timestamp 1746535128
transform 1 0 50496 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _278_
timestamp 1746535128
transform 1 0 53088 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _279_
timestamp 1746535128
transform 1 0 54048 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _280_
timestamp 1746535128
transform 1 0 47904 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _281_
timestamp 1746535128
transform 1 0 37248 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _282_
timestamp 1746535128
transform 1 0 34560 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _283_
timestamp 1746535128
transform 1 0 32064 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _284_
timestamp 1746535128
transform 1 0 29472 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _285_
timestamp 1746535128
transform 1 0 31008 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _286_
timestamp 1746535128
transform 1 0 46176 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _287_
timestamp 1746535128
transform 1 0 47904 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _288_
timestamp 1746535128
transform 1 0 50496 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _289_
timestamp 1746535128
transform 1 0 52224 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _290_
timestamp 1746535128
transform 1 0 54144 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _291_
timestamp 1746535128
transform 1 0 49920 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _292_
timestamp 1746535128
transform 1 0 51936 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _293_
timestamp 1746535128
transform 1 0 42432 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _294_
timestamp 1746535128
transform 1 0 45024 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _295_
timestamp 1746535128
transform 1 0 34272 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _296_
timestamp 1746535128
transform 1 0 31680 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _297_
timestamp 1746535128
transform 1 0 29088 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _298_
timestamp 1746535128
transform 1 0 28032 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _299_
timestamp 1746535128
transform 1 0 27168 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _300_
timestamp 1746535128
transform 1 0 26112 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _301_
timestamp 1746535128
transform 1 0 23328 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _302_
timestamp 1746535128
transform 1 0 19968 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _303_
timestamp 1746535128
transform 1 0 21504 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _304_
timestamp 1746535128
transform 1 0 21792 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _305_
timestamp 1746535128
transform 1 0 23520 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _306_
timestamp 1746535128
transform 1 0 26112 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _307_
timestamp 1746535128
transform 1 0 39840 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _308_
timestamp 1746535128
transform 1 0 38688 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _309_
timestamp 1746535128
transform 1 0 36864 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _310_
timestamp 1746535128
transform 1 0 3360 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _311_
timestamp 1746535128
transform 1 0 2880 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _312_
timestamp 1746535128
transform 1 0 3360 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _313_
timestamp 1746535128
transform 1 0 3360 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _314_
timestamp 1746535128
transform 1 0 11712 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _315_
timestamp 1746535128
transform 1 0 14208 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _316_
timestamp 1746535128
transform 1 0 15168 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _317_
timestamp 1746535128
transform 1 0 3360 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _318_
timestamp 1746535128
transform 1 0 3360 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _319_
timestamp 1746535128
transform 1 0 2496 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _320_
timestamp 1746535128
transform 1 0 768 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _321_
timestamp 1746535128
transform 1 0 1536 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _322_
timestamp 1746535128
transform 1 0 1536 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _323_
timestamp 1746535128
transform 1 0 1632 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _324_
timestamp 1746535128
transform 1 0 1152 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _325_
timestamp 1746535128
transform 1 0 3360 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _326_
timestamp 1746535128
transform 1 0 3360 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _327_
timestamp 1746535128
transform 1 0 16416 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _328_
timestamp 1746535128
transform 1 0 20928 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _329_
timestamp 1746535128
transform 1 0 19104 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _330_
timestamp 1746535128
transform 1 0 15936 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _331_
timestamp 1746535128
transform 1 0 17376 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _332_
timestamp 1746535128
transform 1 0 3360 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _333_
timestamp 1746535128
transform 1 0 3360 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _334_
timestamp 1746535128
transform 1 0 3360 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _335_
timestamp 1746535128
transform 1 0 3360 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _336_
timestamp 1746535128
transform 1 0 3360 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _337_
timestamp 1746535128
transform 1 0 78144 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _338_
timestamp 1746535128
transform 1 0 82656 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _339_
timestamp 1746535128
transform 1 0 80736 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _340_
timestamp 1746535128
transform 1 0 80448 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _341_
timestamp 1746535128
transform 1 0 80352 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _342_
timestamp 1746535128
transform 1 0 80736 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _343_
timestamp 1746535128
transform 1 0 79968 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _344_
timestamp 1746535128
transform 1 0 80160 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _345_
timestamp 1746535128
transform 1 0 80736 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _346_
timestamp 1746535128
transform 1 0 80736 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _347_
timestamp 1746535128
transform 1 0 80736 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _348_
timestamp 1746535128
transform 1 0 80736 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _349_
timestamp 1746535128
transform 1 0 44352 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _350_
timestamp 1746535128
transform 1 0 42048 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _351_
timestamp 1746535128
transform 1 0 40992 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _352_
timestamp 1746535128
transform 1 0 37728 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _353_
timestamp 1746535128
transform 1 0 38400 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _354_
timestamp 1746535128
transform 1 0 40704 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _355_
timestamp 1746535128
transform 1 0 43968 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _356_
timestamp 1746535128
transform 1 0 48576 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _357_
timestamp 1746535128
transform 1 0 17760 0 -1 37044
box -48 -56 2640 834
use sg13g2_dlhq_1  _358_
timestamp 1678805552
transform 1 0 43872 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _359_
timestamp 1678805552
transform 1 0 45984 0 1 2268
box -50 -56 1692 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 38496 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 41088 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 31776 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 32544 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 32544 0 1 2268
box -48 -56 336 834
use sg13g2_buf_16  clkbuf_0_clk
timestamp 1676553496
transform 1 0 62592 0 1 34020
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_0_clk_regs
timestamp 1676553496
transform 1 0 43008 0 1 34020
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_0__f_clk
timestamp 1676553496
transform 1 0 47424 0 1 35532
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_1__f_clk
timestamp 1676553496
transform 1 0 74016 0 1 27972
box -48 -56 2448 834
use sg13g2_buf_8  clkbuf_4_0_0_clk_regs
timestamp 1676451365
transform 1 0 33312 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_1_0_clk_regs
timestamp 1676451365
transform 1 0 37344 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_2_0_clk_regs
timestamp 1676451365
transform 1 0 24192 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_3_0_clk_regs
timestamp 1676451365
transform 1 0 25440 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_4_0_clk_regs
timestamp 1676451365
transform 1 0 7104 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_5_0_clk_regs
timestamp 1676451365
transform 1 0 4704 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_6_0_clk_regs
timestamp 1676451365
transform 1 0 19680 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_7_0_clk_regs
timestamp 1676451365
transform 1 0 16800 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_8_0_clk_regs
timestamp 1676451365
transform 1 0 52512 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_9_0_clk_regs
timestamp 1676451365
transform 1 0 51264 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_10_0_clk_regs
timestamp 1676451365
transform 1 0 61344 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_11_0_clk_regs
timestamp 1676451365
transform 1 0 65760 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_12_0_clk_regs
timestamp 1676451365
transform 1 0 72000 0 1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_13_0_clk_regs
timestamp 1676451365
transform 1 0 70080 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_14_0_clk_regs
timestamp 1676451365
transform 1 0 74016 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_15_0_clk_regs
timestamp 1676451365
transform 1 0 74016 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_16  clkbuf_regs_0_clk
timestamp 1676553496
transform 1 0 43104 0 -1 5292
box -48 -56 2448 834
use sg13g2_inv_1  clkload0
timestamp 1676382929
transform 1 0 15168 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1676382929
transform 1 0 74016 0 -1 24948
box -48 -56 336 834
use sg13g2_buf_16  delaybuf_0_clk
timestamp 1676553496
transform 1 0 32352 0 1 35532
box -48 -56 2448 834
use sg13g2_buf_1  fanout14
timestamp 1676381911
transform 1 0 4224 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout15
timestamp 1676381911
transform 1 0 3456 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout16
timestamp 1676381911
transform 1 0 4800 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout17
timestamp 1676381911
transform 1 0 13632 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout18
timestamp 1676381911
transform 1 0 20928 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout19
timestamp 1676381911
transform 1 0 21408 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  fanout20
timestamp 1676381911
transform 1 0 21120 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout21
timestamp 1676381911
transform 1 0 31008 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout22
timestamp 1676381911
transform 1 0 27456 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout23
timestamp 1676381911
transform 1 0 20544 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform 1 0 42240 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform 1 0 47520 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform 1 0 79872 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform 1 0 80352 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform 1 0 41280 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform 1 0 21696 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout30
timestamp 1676381911
transform 1 0 1824 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform 1 0 2208 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout32
timestamp 1676381911
transform 1 0 2400 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform 1 0 4320 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform 1 0 12192 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform 1 0 26880 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform 1 0 25152 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform 1 0 26496 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform 1 0 23136 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform 1 0 23520 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform 1 0 23904 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform 1 0 5376 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform 1 0 46752 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout43
timestamp 1676381911
transform 1 0 44832 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform 1 0 81600 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform 1 0 81696 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout46
timestamp 1676381911
transform 1 0 45216 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_259
timestamp 1677580104
transform 1 0 25440 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_271
timestamp 1679581782
transform 1 0 26592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_278
timestamp 1679581782
transform 1 0 27264 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_285
timestamp 1677579658
transform 1 0 27936 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_313
timestamp 1679581782
transform 1 0 30624 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_320
timestamp 1677579658
transform 1 0 31296 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_331
timestamp 1679581782
transform 1 0 32352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_338
timestamp 1679581782
transform 1 0 33024 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_345
timestamp 1677580104
transform 1 0 33696 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_347
timestamp 1677579658
transform 1 0 33888 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_358
timestamp 1679581782
transform 1 0 34944 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_369
timestamp 1679577901
transform 1 0 36000 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_373
timestamp 1677579658
transform 1 0 36384 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_384
timestamp 1679581782
transform 1 0 37440 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_391
timestamp 1679577901
transform 1 0 38112 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_395
timestamp 1677580104
transform 1 0 38496 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_424
timestamp 1679581782
transform 1 0 41280 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_431
timestamp 1677579658
transform 1 0 41952 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_442
timestamp 1679581782
transform 1 0 43008 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_449
timestamp 1679577901
transform 1 0 43680 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_453
timestamp 1677580104
transform 1 0 44064 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_465
timestamp 1679581782
transform 1 0 45216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_472
timestamp 1679581782
transform 1 0 45888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_479
timestamp 1679581782
transform 1 0 46560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_486
timestamp 1679581782
transform 1 0 47232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_493
timestamp 1679581782
transform 1 0 47904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_500
timestamp 1679581782
transform 1 0 48576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_507
timestamp 1679581782
transform 1 0 49248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_514
timestamp 1679581782
transform 1 0 49920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_521
timestamp 1679581782
transform 1 0 50592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_538
timestamp 1679581782
transform 1 0 52224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_545
timestamp 1679581782
transform 1 0 52896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_552
timestamp 1679581782
transform 1 0 53568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_559
timestamp 1679581782
transform 1 0 54240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_566
timestamp 1679581782
transform 1 0 54912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_573
timestamp 1679581782
transform 1 0 55584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_580
timestamp 1679581782
transform 1 0 56256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_587
timestamp 1679581782
transform 1 0 56928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_594
timestamp 1679581782
transform 1 0 57600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_601
timestamp 1679581782
transform 1 0 58272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_608
timestamp 1679581782
transform 1 0 58944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_615
timestamp 1679581782
transform 1 0 59616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_622
timestamp 1679581782
transform 1 0 60288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_629
timestamp 1679581782
transform 1 0 60960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_636
timestamp 1679581782
transform 1 0 61632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_643
timestamp 1679581782
transform 1 0 62304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_650
timestamp 1679581782
transform 1 0 62976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_657
timestamp 1679581782
transform 1 0 63648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_664
timestamp 1679581782
transform 1 0 64320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_671
timestamp 1679581782
transform 1 0 64992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_678
timestamp 1679581782
transform 1 0 65664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_685
timestamp 1679581782
transform 1 0 66336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_692
timestamp 1679581782
transform 1 0 67008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_699
timestamp 1679581782
transform 1 0 67680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_706
timestamp 1679581782
transform 1 0 68352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_713
timestamp 1679581782
transform 1 0 69024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_720
timestamp 1679581782
transform 1 0 69696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_727
timestamp 1679581782
transform 1 0 70368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_734
timestamp 1679581782
transform 1 0 71040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_741
timestamp 1679581782
transform 1 0 71712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_748
timestamp 1679581782
transform 1 0 72384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_755
timestamp 1679581782
transform 1 0 73056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_762
timestamp 1679581782
transform 1 0 73728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_769
timestamp 1679581782
transform 1 0 74400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_776
timestamp 1679581782
transform 1 0 75072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_783
timestamp 1679581782
transform 1 0 75744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_790
timestamp 1679581782
transform 1 0 76416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_797
timestamp 1679581782
transform 1 0 77088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_804
timestamp 1679581782
transform 1 0 77760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_811
timestamp 1679581782
transform 1 0 78432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_818
timestamp 1679581782
transform 1 0 79104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_825
timestamp 1679581782
transform 1 0 79776 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_832
timestamp 1677580104
transform 1 0 80448 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_834
timestamp 1677579658
transform 1 0 80640 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_217
timestamp 1677580104
transform 1 0 21408 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_293
timestamp 1679577901
transform 1 0 28704 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_1_405
timestamp 1679577901
transform 1 0 39456 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_527
timestamp 1679581782
transform 1 0 51168 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_534
timestamp 1677579658
transform 1 0 51840 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_562
timestamp 1679581782
transform 1 0 54528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_569
timestamp 1679581782
transform 1 0 55200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_576
timestamp 1679581782
transform 1 0 55872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_583
timestamp 1679581782
transform 1 0 56544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_590
timestamp 1679581782
transform 1 0 57216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_597
timestamp 1679581782
transform 1 0 57888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_604
timestamp 1679581782
transform 1 0 58560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_611
timestamp 1679581782
transform 1 0 59232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_618
timestamp 1679581782
transform 1 0 59904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_625
timestamp 1679581782
transform 1 0 60576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_632
timestamp 1679581782
transform 1 0 61248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_639
timestamp 1679581782
transform 1 0 61920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_646
timestamp 1679581782
transform 1 0 62592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_653
timestamp 1679581782
transform 1 0 63264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_660
timestamp 1679581782
transform 1 0 63936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_667
timestamp 1679581782
transform 1 0 64608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_674
timestamp 1679581782
transform 1 0 65280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_681
timestamp 1679581782
transform 1 0 65952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_688
timestamp 1679581782
transform 1 0 66624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_695
timestamp 1679581782
transform 1 0 67296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_702
timestamp 1679581782
transform 1 0 67968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_709
timestamp 1679581782
transform 1 0 68640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_716
timestamp 1679581782
transform 1 0 69312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_723
timestamp 1679581782
transform 1 0 69984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_730
timestamp 1679581782
transform 1 0 70656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_737
timestamp 1679581782
transform 1 0 71328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_744
timestamp 1679581782
transform 1 0 72000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_751
timestamp 1679581782
transform 1 0 72672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_758
timestamp 1679581782
transform 1 0 73344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_765
timestamp 1679581782
transform 1 0 74016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_772
timestamp 1679581782
transform 1 0 74688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_779
timestamp 1679581782
transform 1 0 75360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_786
timestamp 1679581782
transform 1 0 76032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_793
timestamp 1679581782
transform 1 0 76704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_800
timestamp 1679581782
transform 1 0 77376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_807
timestamp 1679581782
transform 1 0 78048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_814
timestamp 1679581782
transform 1 0 78720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_821
timestamp 1679581782
transform 1 0 79392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_828
timestamp 1679581782
transform 1 0 80064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_200
timestamp 1679581782
transform 1 0 19776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_207
timestamp 1679581782
transform 1 0 20448 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_214
timestamp 1677580104
transform 1 0 21120 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_216
timestamp 1677579658
transform 1 0 21312 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_248
timestamp 1679581782
transform 1 0 24384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_255
timestamp 1679581782
transform 1 0 25056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_262
timestamp 1679581782
transform 1 0 25728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_269
timestamp 1679581782
transform 1 0 26400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_276
timestamp 1679577901
transform 1 0 27072 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_280
timestamp 1677580104
transform 1 0 27456 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_292
timestamp 1679577901
transform 1 0 28608 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_296
timestamp 1677580104
transform 1 0 28992 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_308
timestamp 1679581782
transform 1 0 30144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_315
timestamp 1679581782
transform 1 0 30816 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_322
timestamp 1677579658
transform 1 0 31488 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_336
timestamp 1679581782
transform 1 0 32832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_343
timestamp 1679581782
transform 1 0 33504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_350
timestamp 1679577901
transform 1 0 34176 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_354
timestamp 1677580104
transform 1 0 34560 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_360
timestamp 1679581782
transform 1 0 35136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_367
timestamp 1679581782
transform 1 0 35808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_374
timestamp 1679581782
transform 1 0 36480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_381
timestamp 1679581782
transform 1 0 37152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_388
timestamp 1679581782
transform 1 0 37824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_405
timestamp 1679577901
transform 1 0 39456 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_419
timestamp 1679581782
transform 1 0 40800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_426
timestamp 1679581782
transform 1 0 41472 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_433
timestamp 1677579658
transform 1 0 42144 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_445
timestamp 1679581782
transform 1 0 43296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_452
timestamp 1679581782
transform 1 0 43968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_459
timestamp 1679581782
transform 1 0 44640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_490
timestamp 1679581782
transform 1 0 47616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_497
timestamp 1679581782
transform 1 0 48288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_541
timestamp 1679581782
transform 1 0 52512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_548
timestamp 1679581782
transform 1 0 53184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_555
timestamp 1679581782
transform 1 0 53856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_562
timestamp 1679581782
transform 1 0 54528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_569
timestamp 1679581782
transform 1 0 55200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_576
timestamp 1679581782
transform 1 0 55872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_583
timestamp 1679581782
transform 1 0 56544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_590
timestamp 1679581782
transform 1 0 57216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_597
timestamp 1679581782
transform 1 0 57888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_604
timestamp 1679581782
transform 1 0 58560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_611
timestamp 1679581782
transform 1 0 59232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_618
timestamp 1679581782
transform 1 0 59904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_625
timestamp 1679581782
transform 1 0 60576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_632
timestamp 1679581782
transform 1 0 61248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_639
timestamp 1679581782
transform 1 0 61920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_646
timestamp 1679581782
transform 1 0 62592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_653
timestamp 1679581782
transform 1 0 63264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_660
timestamp 1679581782
transform 1 0 63936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_667
timestamp 1679581782
transform 1 0 64608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_674
timestamp 1679581782
transform 1 0 65280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_681
timestamp 1679581782
transform 1 0 65952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_688
timestamp 1679581782
transform 1 0 66624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_695
timestamp 1679581782
transform 1 0 67296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_702
timestamp 1679581782
transform 1 0 67968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_709
timestamp 1679581782
transform 1 0 68640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_716
timestamp 1679581782
transform 1 0 69312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_723
timestamp 1679581782
transform 1 0 69984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_730
timestamp 1679581782
transform 1 0 70656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_737
timestamp 1679581782
transform 1 0 71328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_744
timestamp 1679581782
transform 1 0 72000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_751
timestamp 1679581782
transform 1 0 72672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_758
timestamp 1679581782
transform 1 0 73344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_765
timestamp 1679581782
transform 1 0 74016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_772
timestamp 1679581782
transform 1 0 74688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_779
timestamp 1679581782
transform 1 0 75360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_786
timestamp 1679581782
transform 1 0 76032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_793
timestamp 1679581782
transform 1 0 76704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_800
timestamp 1679581782
transform 1 0 77376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_807
timestamp 1679581782
transform 1 0 78048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_814
timestamp 1679581782
transform 1 0 78720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_821
timestamp 1679581782
transform 1 0 79392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_828
timestamp 1679581782
transform 1 0 80064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 13728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 15744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_165
timestamp 1679577901
transform 1 0 16416 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 17760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679581782
transform 1 0 18432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679581782
transform 1 0 19104 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_200
timestamp 1677580104
transform 1 0 19776 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_202
timestamp 1677579658
transform 1 0 19968 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_213
timestamp 1677579658
transform 1 0 21024 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 24096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679581782
transform 1 0 24768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679581782
transform 1 0 25440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_293
timestamp 1679581782
transform 1 0 28704 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_300
timestamp 1677579658
transform 1 0 29376 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_328
timestamp 1677579658
transform 1 0 32064 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_334
timestamp 1679581782
transform 1 0 32640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_341
timestamp 1679581782
transform 1 0 33312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_348
timestamp 1679581782
transform 1 0 33984 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_355
timestamp 1677579658
transform 1 0 34656 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_362
timestamp 1679581782
transform 1 0 35328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_369
timestamp 1679581782
transform 1 0 36000 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_376
timestamp 1677580104
transform 1 0 36672 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_384
timestamp 1679581782
transform 1 0 37440 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_391
timestamp 1677579658
transform 1 0 38112 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_398
timestamp 1679581782
transform 1 0 38784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_405
timestamp 1679581782
transform 1 0 39456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_412
timestamp 1679581782
transform 1 0 40128 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_419
timestamp 1677579658
transform 1 0 40800 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_425
timestamp 1679581782
transform 1 0 41376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_432
timestamp 1679581782
transform 1 0 42048 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_439
timestamp 1677580104
transform 1 0 42720 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_446
timestamp 1679577901
transform 1 0 43392 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_450
timestamp 1677579658
transform 1 0 43776 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_468
timestamp 1679581782
transform 1 0 45504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_502
timestamp 1679581782
transform 1 0 48768 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_509
timestamp 1677580104
transform 1 0 49440 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_521
timestamp 1679581782
transform 1 0 50592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_528
timestamp 1679581782
transform 1 0 51264 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_535
timestamp 1677580104
transform 1 0 51936 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_537
timestamp 1677579658
transform 1 0 52128 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_565
timestamp 1679581782
transform 1 0 54816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_572
timestamp 1679581782
transform 1 0 55488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_579
timestamp 1679581782
transform 1 0 56160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_586
timestamp 1679581782
transform 1 0 56832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_593
timestamp 1679581782
transform 1 0 57504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_600
timestamp 1679581782
transform 1 0 58176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_607
timestamp 1679581782
transform 1 0 58848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_614
timestamp 1679581782
transform 1 0 59520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_621
timestamp 1679581782
transform 1 0 60192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_628
timestamp 1679581782
transform 1 0 60864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_635
timestamp 1679581782
transform 1 0 61536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_642
timestamp 1679581782
transform 1 0 62208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_649
timestamp 1679581782
transform 1 0 62880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_656
timestamp 1679581782
transform 1 0 63552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_663
timestamp 1679581782
transform 1 0 64224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_670
timestamp 1679581782
transform 1 0 64896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_677
timestamp 1679581782
transform 1 0 65568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_684
timestamp 1679581782
transform 1 0 66240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_691
timestamp 1679581782
transform 1 0 66912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_698
timestamp 1679581782
transform 1 0 67584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_705
timestamp 1679581782
transform 1 0 68256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_712
timestamp 1679581782
transform 1 0 68928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_719
timestamp 1679581782
transform 1 0 69600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_726
timestamp 1679581782
transform 1 0 70272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_733
timestamp 1679581782
transform 1 0 70944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_740
timestamp 1679581782
transform 1 0 71616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_747
timestamp 1679581782
transform 1 0 72288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_754
timestamp 1679581782
transform 1 0 72960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_761
timestamp 1679581782
transform 1 0 73632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_768
timestamp 1679581782
transform 1 0 74304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_775
timestamp 1679581782
transform 1 0 74976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_782
timestamp 1679581782
transform 1 0 75648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_789
timestamp 1679581782
transform 1 0 76320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_796
timestamp 1679581782
transform 1 0 76992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_803
timestamp 1679581782
transform 1 0 77664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_810
timestamp 1679581782
transform 1 0 78336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_817
timestamp 1679581782
transform 1 0 79008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_824
timestamp 1679581782
transform 1 0 79680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_831
timestamp 1679577901
transform 1 0 80352 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_109
timestamp 1679581782
transform 1 0 11040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_116
timestamp 1679581782
transform 1 0 11712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_123
timestamp 1679581782
transform 1 0 12384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679581782
transform 1 0 13056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 15744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_229
timestamp 1679581782
transform 1 0 22560 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_236
timestamp 1677579658
transform 1 0 23232 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_264
timestamp 1677580104
transform 1 0 25920 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_266
timestamp 1677579658
transform 1 0 26112 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_304
timestamp 1677580104
transform 1 0 29760 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_306
timestamp 1677579658
transform 1 0 29952 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_344
timestamp 1679581782
transform 1 0 33600 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_351
timestamp 1677580104
transform 1 0 34272 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_353
timestamp 1677579658
transform 1 0 34464 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_363
timestamp 1679581782
transform 1 0 35424 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_370
timestamp 1677579658
transform 1 0 36096 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_375
timestamp 1679581782
transform 1 0 36576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_382
timestamp 1679581782
transform 1 0 37248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_389
timestamp 1679577901
transform 1 0 37920 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_393
timestamp 1677580104
transform 1 0 38304 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_398
timestamp 1679581782
transform 1 0 38784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_405
timestamp 1679577901
transform 1 0 39456 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_409
timestamp 1677579658
transform 1 0 39840 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_415
timestamp 1677580104
transform 1 0 40416 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_425
timestamp 1679581782
transform 1 0 41376 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_432
timestamp 1677580104
transform 1 0 42048 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_459
timestamp 1679581782
transform 1 0 44640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_466
timestamp 1679577901
transform 1 0 45312 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_480
timestamp 1677580104
transform 1 0 46656 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_482
timestamp 1677579658
transform 1 0 46848 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_547
timestamp 1677579658
transform 1 0 53088 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_585
timestamp 1679581782
transform 1 0 56736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_592
timestamp 1679581782
transform 1 0 57408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_599
timestamp 1679581782
transform 1 0 58080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_606
timestamp 1679581782
transform 1 0 58752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_613
timestamp 1679581782
transform 1 0 59424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_620
timestamp 1679581782
transform 1 0 60096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_627
timestamp 1679581782
transform 1 0 60768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_634
timestamp 1679581782
transform 1 0 61440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_641
timestamp 1679581782
transform 1 0 62112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_648
timestamp 1679581782
transform 1 0 62784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_655
timestamp 1679581782
transform 1 0 63456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_662
timestamp 1679581782
transform 1 0 64128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_669
timestamp 1679581782
transform 1 0 64800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_676
timestamp 1679581782
transform 1 0 65472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_683
timestamp 1679581782
transform 1 0 66144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_690
timestamp 1679581782
transform 1 0 66816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_697
timestamp 1679581782
transform 1 0 67488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_704
timestamp 1679581782
transform 1 0 68160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_711
timestamp 1679581782
transform 1 0 68832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_718
timestamp 1679581782
transform 1 0 69504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_725
timestamp 1679581782
transform 1 0 70176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_732
timestamp 1679581782
transform 1 0 70848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_739
timestamp 1679581782
transform 1 0 71520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_746
timestamp 1679581782
transform 1 0 72192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_753
timestamp 1679581782
transform 1 0 72864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_760
timestamp 1679581782
transform 1 0 73536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_767
timestamp 1679581782
transform 1 0 74208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_774
timestamp 1679581782
transform 1 0 74880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_781
timestamp 1679581782
transform 1 0 75552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_788
timestamp 1679581782
transform 1 0 76224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_795
timestamp 1679581782
transform 1 0 76896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_802
timestamp 1679581782
transform 1 0 77568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_809
timestamp 1679581782
transform 1 0 78240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_816
timestamp 1679581782
transform 1 0 78912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_823
timestamp 1679581782
transform 1 0 79584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_830
timestamp 1679577901
transform 1 0 80256 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_834
timestamp 1677579658
transform 1 0 80640 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_158
timestamp 1677580104
transform 1 0 15744 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_187
timestamp 1679581782
transform 1 0 18528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_194
timestamp 1679581782
transform 1 0 19200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_201
timestamp 1679581782
transform 1 0 19872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_208
timestamp 1679581782
transform 1 0 20544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_225
timestamp 1679581782
transform 1 0 22176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_232
timestamp 1679581782
transform 1 0 22848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_239
timestamp 1679577901
transform 1 0 23520 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_253
timestamp 1677580104
transform 1 0 24864 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_255
timestamp 1677579658
transform 1 0 25056 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_278
timestamp 1679581782
transform 1 0 27264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_285
timestamp 1679581782
transform 1 0 27936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_292
timestamp 1679581782
transform 1 0 28608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_299
timestamp 1679581782
transform 1 0 29280 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_306
timestamp 1677580104
transform 1 0 29952 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_318
timestamp 1679581782
transform 1 0 31104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_336
timestamp 1679581782
transform 1 0 32832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_343
timestamp 1679581782
transform 1 0 33504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_350
timestamp 1679581782
transform 1 0 34176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_357
timestamp 1679581782
transform 1 0 34848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_364
timestamp 1679581782
transform 1 0 35520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_371
timestamp 1679581782
transform 1 0 36192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_382
timestamp 1679581782
transform 1 0 37248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_389
timestamp 1679577901
transform 1 0 37920 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_393
timestamp 1677580104
transform 1 0 38304 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_405
timestamp 1679581782
transform 1 0 39456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_412
timestamp 1679581782
transform 1 0 40128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_419
timestamp 1679581782
transform 1 0 40800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_426
timestamp 1679581782
transform 1 0 41472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_433
timestamp 1679581782
transform 1 0 42144 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_440
timestamp 1677580104
transform 1 0 42816 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_442
timestamp 1677579658
transform 1 0 43008 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_468
timestamp 1679581782
transform 1 0 45504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_475
timestamp 1679577901
transform 1 0 46176 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_479
timestamp 1677580104
transform 1 0 46560 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_485
timestamp 1679581782
transform 1 0 47136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_492
timestamp 1679581782
transform 1 0 47808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_499
timestamp 1679581782
transform 1 0 48480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_506
timestamp 1679581782
transform 1 0 49152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_513
timestamp 1679581782
transform 1 0 49824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_520
timestamp 1679581782
transform 1 0 50496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_527
timestamp 1679577901
transform 1 0 51168 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_541
timestamp 1679581782
transform 1 0 52512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_548
timestamp 1679581782
transform 1 0 53184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_555
timestamp 1679581782
transform 1 0 53856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_562
timestamp 1679581782
transform 1 0 54528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_569
timestamp 1679581782
transform 1 0 55200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_576
timestamp 1679581782
transform 1 0 55872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_583
timestamp 1679581782
transform 1 0 56544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_590
timestamp 1679581782
transform 1 0 57216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_597
timestamp 1679581782
transform 1 0 57888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_604
timestamp 1679581782
transform 1 0 58560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_611
timestamp 1679581782
transform 1 0 59232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_618
timestamp 1679581782
transform 1 0 59904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_625
timestamp 1679581782
transform 1 0 60576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_632
timestamp 1679581782
transform 1 0 61248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_639
timestamp 1679581782
transform 1 0 61920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_646
timestamp 1679581782
transform 1 0 62592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_653
timestamp 1679581782
transform 1 0 63264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_660
timestamp 1679581782
transform 1 0 63936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_667
timestamp 1679581782
transform 1 0 64608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_674
timestamp 1679581782
transform 1 0 65280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_681
timestamp 1679581782
transform 1 0 65952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_688
timestamp 1679581782
transform 1 0 66624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_695
timestamp 1679581782
transform 1 0 67296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_702
timestamp 1679581782
transform 1 0 67968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_709
timestamp 1679581782
transform 1 0 68640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_716
timestamp 1679581782
transform 1 0 69312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_723
timestamp 1679581782
transform 1 0 69984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_730
timestamp 1679581782
transform 1 0 70656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_737
timestamp 1679581782
transform 1 0 71328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_744
timestamp 1679581782
transform 1 0 72000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_751
timestamp 1679581782
transform 1 0 72672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_758
timestamp 1679581782
transform 1 0 73344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_765
timestamp 1679581782
transform 1 0 74016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_772
timestamp 1679581782
transform 1 0 74688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_779
timestamp 1679581782
transform 1 0 75360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_786
timestamp 1679581782
transform 1 0 76032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_793
timestamp 1679581782
transform 1 0 76704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_800
timestamp 1679581782
transform 1 0 77376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_807
timestamp 1679581782
transform 1 0 78048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_814
timestamp 1679581782
transform 1 0 78720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_821
timestamp 1679581782
transform 1 0 79392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_828
timestamp 1679581782
transform 1 0 80064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679581782
transform 1 0 3648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679581782
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679581782
transform 1 0 4992 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_53
timestamp 1677580104
transform 1 0 5664 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_55
timestamp 1677579658
transform 1 0 5856 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_765
timestamp 1679581782
transform 1 0 74016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_772
timestamp 1679581782
transform 1 0 74688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_779
timestamp 1679581782
transform 1 0 75360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_786
timestamp 1679581782
transform 1 0 76032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_793
timestamp 1679581782
transform 1 0 76704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_800
timestamp 1679581782
transform 1 0 77376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_807
timestamp 1679581782
transform 1 0 78048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_814
timestamp 1679581782
transform 1 0 78720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_821
timestamp 1679581782
transform 1 0 79392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_828
timestamp 1679581782
transform 1 0 80064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_765
timestamp 1679581782
transform 1 0 74016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_772
timestamp 1679581782
transform 1 0 74688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_779
timestamp 1679581782
transform 1 0 75360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_786
timestamp 1679581782
transform 1 0 76032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_793
timestamp 1679581782
transform 1 0 76704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_800
timestamp 1679581782
transform 1 0 77376 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_807
timestamp 1677579658
transform 1 0 78048 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_833
timestamp 1677580104
transform 1 0 80544 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_32
timestamp 1679577901
transform 1 0 3648 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_36
timestamp 1677580104
transform 1 0 4032 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_48
timestamp 1679581782
transform 1 0 5184 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_55
timestamp 1677579658
transform 1 0 5856 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_765
timestamp 1679581782
transform 1 0 74016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_772
timestamp 1679581782
transform 1 0 74688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_779
timestamp 1679581782
transform 1 0 75360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_786
timestamp 1679581782
transform 1 0 76032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_793
timestamp 1679581782
transform 1 0 76704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_800
timestamp 1679581782
transform 1 0 77376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_807
timestamp 1679581782
transform 1 0 78048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_814
timestamp 1679581782
transform 1 0 78720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_821
timestamp 1679581782
transform 1 0 79392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_828
timestamp 1679581782
transform 1 0 80064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_25
timestamp 1679577901
transform 1 0 2976 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_765
timestamp 1679581782
transform 1 0 74016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_772
timestamp 1679581782
transform 1 0 74688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_779
timestamp 1679581782
transform 1 0 75360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_786
timestamp 1679581782
transform 1 0 76032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_793
timestamp 1679581782
transform 1 0 76704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_800
timestamp 1679581782
transform 1 0 77376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_807
timestamp 1679581782
transform 1 0 78048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_814
timestamp 1679581782
transform 1 0 78720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_821
timestamp 1679581782
transform 1 0 79392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_828
timestamp 1679581782
transform 1 0 80064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679581782
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679581782
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679581782
transform 1 0 2976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679581782
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679581782
transform 1 0 4320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_46
timestamp 1679581782
transform 1 0 4992 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_53
timestamp 1677580104
transform 1 0 5664 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_55
timestamp 1677579658
transform 1 0 5856 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_765
timestamp 1679581782
transform 1 0 74016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_772
timestamp 1679581782
transform 1 0 74688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_779
timestamp 1679581782
transform 1 0 75360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_786
timestamp 1679581782
transform 1 0 76032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_793
timestamp 1679581782
transform 1 0 76704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_800
timestamp 1679581782
transform 1 0 77376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_807
timestamp 1679581782
transform 1 0 78048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_814
timestamp 1679581782
transform 1 0 78720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_821
timestamp 1679581782
transform 1 0 79392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_828
timestamp 1679581782
transform 1 0 80064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679581782
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_32
timestamp 1677580104
transform 1 0 3648 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_44
timestamp 1679581782
transform 1 0 4800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_51
timestamp 1679577901
transform 1 0 5472 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_55
timestamp 1677579658
transform 1 0 5856 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_765
timestamp 1679581782
transform 1 0 74016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_772
timestamp 1679581782
transform 1 0 74688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_779
timestamp 1679581782
transform 1 0 75360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_786
timestamp 1679581782
transform 1 0 76032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_793
timestamp 1679581782
transform 1 0 76704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_800
timestamp 1679581782
transform 1 0 77376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_807
timestamp 1679581782
transform 1 0 78048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_814
timestamp 1679581782
transform 1 0 78720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_821
timestamp 1679581782
transform 1 0 79392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_828
timestamp 1679581782
transform 1 0 80064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679581782
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679581782
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679581782
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_25
timestamp 1679577901
transform 1 0 2976 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_765
timestamp 1679581782
transform 1 0 74016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_772
timestamp 1679581782
transform 1 0 74688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_779
timestamp 1679581782
transform 1 0 75360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_786
timestamp 1679581782
transform 1 0 76032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_793
timestamp 1679581782
transform 1 0 76704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_800
timestamp 1679581782
transform 1 0 77376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_807
timestamp 1679581782
transform 1 0 78048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_814
timestamp 1679581782
transform 1 0 78720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_821
timestamp 1679581782
transform 1 0 79392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_828
timestamp 1679581782
transform 1 0 80064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_4
timestamp 1679577901
transform 1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_8
timestamp 1677580104
transform 1 0 1344 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_47
timestamp 1679581782
transform 1 0 5088 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_54
timestamp 1677580104
transform 1 0 5760 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_765
timestamp 1679581782
transform 1 0 74016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_772
timestamp 1679581782
transform 1 0 74688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_779
timestamp 1679581782
transform 1 0 75360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_786
timestamp 1679581782
transform 1 0 76032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_793
timestamp 1679581782
transform 1 0 76704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_800
timestamp 1679581782
transform 1 0 77376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_807
timestamp 1679581782
transform 1 0 78048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_814
timestamp 1679581782
transform 1 0 78720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_821
timestamp 1679581782
transform 1 0 79392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_828
timestamp 1679581782
transform 1 0 80064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679581782
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679581782
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679581782
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_32
timestamp 1677579658
transform 1 0 3648 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_43
timestamp 1679581782
transform 1 0 4704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_50
timestamp 1679577901
transform 1 0 5376 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_54
timestamp 1677580104
transform 1 0 5760 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_765
timestamp 1679581782
transform 1 0 74016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_772
timestamp 1679581782
transform 1 0 74688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_779
timestamp 1679581782
transform 1 0 75360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_786
timestamp 1679581782
transform 1 0 76032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_793
timestamp 1679581782
transform 1 0 76704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_800
timestamp 1679581782
transform 1 0 77376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_807
timestamp 1679581782
transform 1 0 78048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_814
timestamp 1679581782
transform 1 0 78720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_821
timestamp 1679581782
transform 1 0 79392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_828
timestamp 1679581782
transform 1 0 80064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679581782
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_25
timestamp 1679577901
transform 1 0 2976 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_765
timestamp 1679581782
transform 1 0 74016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_772
timestamp 1679581782
transform 1 0 74688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_779
timestamp 1679581782
transform 1 0 75360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_786
timestamp 1679581782
transform 1 0 76032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_793
timestamp 1679581782
transform 1 0 76704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_800
timestamp 1679581782
transform 1 0 77376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_807
timestamp 1679581782
transform 1 0 78048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_814
timestamp 1679581782
transform 1 0 78720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_821
timestamp 1679581782
transform 1 0 79392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_828
timestamp 1679581782
transform 1 0 80064 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_0
timestamp 1677580104
transform 1 0 576 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_765
timestamp 1679581782
transform 1 0 74016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_772
timestamp 1679581782
transform 1 0 74688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_779
timestamp 1679581782
transform 1 0 75360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_786
timestamp 1679581782
transform 1 0 76032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_793
timestamp 1679581782
transform 1 0 76704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_800
timestamp 1679581782
transform 1 0 77376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_807
timestamp 1679581782
transform 1 0 78048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_814
timestamp 1679581782
transform 1 0 78720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_821
timestamp 1679581782
transform 1 0 79392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_828
timestamp 1679581782
transform 1 0 80064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_7
timestamp 1677579658
transform 1 0 1248 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_18
timestamp 1679581782
transform 1 0 2304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_25
timestamp 1679577901
transform 1 0 2976 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_29
timestamp 1677579658
transform 1 0 3360 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_40
timestamp 1679581782
transform 1 0 4416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_47
timestamp 1679581782
transform 1 0 5088 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_54
timestamp 1677580104
transform 1 0 5760 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_765
timestamp 1679581782
transform 1 0 74016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_772
timestamp 1679581782
transform 1 0 74688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_779
timestamp 1679581782
transform 1 0 75360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_786
timestamp 1679581782
transform 1 0 76032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_793
timestamp 1679581782
transform 1 0 76704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_800
timestamp 1679581782
transform 1 0 77376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_807
timestamp 1679581782
transform 1 0 78048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_814
timestamp 1679581782
transform 1 0 78720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_821
timestamp 1679581782
transform 1 0 79392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_828
timestamp 1679581782
transform 1 0 80064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_4
timestamp 1679577901
transform 1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_8
timestamp 1677580104
transform 1 0 1344 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_47
timestamp 1679581782
transform 1 0 5088 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_54
timestamp 1677580104
transform 1 0 5760 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_765
timestamp 1679581782
transform 1 0 74016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_772
timestamp 1679581782
transform 1 0 74688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_779
timestamp 1679581782
transform 1 0 75360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_786
timestamp 1679581782
transform 1 0 76032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_793
timestamp 1679581782
transform 1 0 76704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_800
timestamp 1679581782
transform 1 0 77376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_807
timestamp 1679581782
transform 1 0 78048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_814
timestamp 1679581782
transform 1 0 78720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_821
timestamp 1679581782
transform 1 0 79392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_828
timestamp 1679581782
transform 1 0 80064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_4
timestamp 1679577901
transform 1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679581782
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_25
timestamp 1679577901
transform 1 0 2976 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_765
timestamp 1679581782
transform 1 0 74016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_772
timestamp 1679581782
transform 1 0 74688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_779
timestamp 1679581782
transform 1 0 75360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_786
timestamp 1679581782
transform 1 0 76032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_793
timestamp 1679581782
transform 1 0 76704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_800
timestamp 1679581782
transform 1 0 77376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_807
timestamp 1679581782
transform 1 0 78048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_814
timestamp 1679581782
transform 1 0 78720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_821
timestamp 1679581782
transform 1 0 79392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_828
timestamp 1679581782
transform 1 0 80064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_4
timestamp 1679577901
transform 1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_8
timestamp 1677580104
transform 1 0 1344 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_47
timestamp 1679581782
transform 1 0 5088 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_54
timestamp 1677580104
transform 1 0 5760 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_765
timestamp 1679581782
transform 1 0 74016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_772
timestamp 1679581782
transform 1 0 74688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_779
timestamp 1679581782
transform 1 0 75360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_786
timestamp 1679581782
transform 1 0 76032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_793
timestamp 1679581782
transform 1 0 76704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_800
timestamp 1679581782
transform 1 0 77376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_807
timestamp 1679581782
transform 1 0 78048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_814
timestamp 1679581782
transform 1 0 78720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_821
timestamp 1679581782
transform 1 0 79392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_828
timestamp 1679581782
transform 1 0 80064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_8
timestamp 1679581782
transform 1 0 1344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_15
timestamp 1679581782
transform 1 0 2016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_22
timestamp 1679581782
transform 1 0 2688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_765
timestamp 1679581782
transform 1 0 74016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_772
timestamp 1679581782
transform 1 0 74688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_779
timestamp 1679581782
transform 1 0 75360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_786
timestamp 1679581782
transform 1 0 76032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_793
timestamp 1679577901
transform 1 0 76704 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_797
timestamp 1677579658
transform 1 0 77088 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_0
timestamp 1677579658
transform 1 0 576 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_42
timestamp 1679581782
transform 1 0 4608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_49
timestamp 1679581782
transform 1 0 5280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_765
timestamp 1679581782
transform 1 0 74016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_772
timestamp 1679581782
transform 1 0 74688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_779
timestamp 1679581782
transform 1 0 75360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_786
timestamp 1679581782
transform 1 0 76032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_793
timestamp 1679581782
transform 1 0 76704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_800
timestamp 1679581782
transform 1 0 77376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_807
timestamp 1679581782
transform 1 0 78048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_814
timestamp 1679581782
transform 1 0 78720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_821
timestamp 1679581782
transform 1 0 79392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_828
timestamp 1679581782
transform 1 0 80064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_11
timestamp 1677580104
transform 1 0 1632 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_21
timestamp 1679581782
transform 1 0 2592 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_28
timestamp 1677579658
transform 1 0 3264 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_765
timestamp 1679581782
transform 1 0 74016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_772
timestamp 1679581782
transform 1 0 74688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_779
timestamp 1679581782
transform 1 0 75360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_786
timestamp 1679581782
transform 1 0 76032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_793
timestamp 1679581782
transform 1 0 76704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_800
timestamp 1679581782
transform 1 0 77376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_807
timestamp 1679581782
transform 1 0 78048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_814
timestamp 1679581782
transform 1 0 78720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_821
timestamp 1679581782
transform 1 0 79392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_828
timestamp 1679581782
transform 1 0 80064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_4
timestamp 1679577901
transform 1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_8
timestamp 1677579658
transform 1 0 1344 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_23
timestamp 1679581782
transform 1 0 2784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_48
timestamp 1679581782
transform 1 0 5184 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_55
timestamp 1677579658
transform 1 0 5856 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_765
timestamp 1679581782
transform 1 0 74016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_772
timestamp 1679581782
transform 1 0 74688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_779
timestamp 1679581782
transform 1 0 75360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_786
timestamp 1679581782
transform 1 0 76032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_793
timestamp 1679581782
transform 1 0 76704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_800
timestamp 1679581782
transform 1 0 77376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_807
timestamp 1679581782
transform 1 0 78048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_814
timestamp 1679581782
transform 1 0 78720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_821
timestamp 1679581782
transform 1 0 79392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_828
timestamp 1679581782
transform 1 0 80064 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_4
timestamp 1677580104
transform 1 0 960 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_43
timestamp 1679581782
transform 1 0 4704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_50
timestamp 1679577901
transform 1 0 5376 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_54
timestamp 1677580104
transform 1 0 5760 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_765
timestamp 1679581782
transform 1 0 74016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_772
timestamp 1679581782
transform 1 0 74688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_779
timestamp 1679581782
transform 1 0 75360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_786
timestamp 1679581782
transform 1 0 76032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_793
timestamp 1679581782
transform 1 0 76704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_800
timestamp 1679581782
transform 1 0 77376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_807
timestamp 1679581782
transform 1 0 78048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_814
timestamp 1679581782
transform 1 0 78720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_821
timestamp 1679581782
transform 1 0 79392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_828
timestamp 1679581782
transform 1 0 80064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_835
timestamp 1679581782
transform 1 0 80736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_842
timestamp 1679581782
transform 1 0 81408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_849
timestamp 1679581782
transform 1 0 82080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_856
timestamp 1679581782
transform 1 0 82752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_863
timestamp 1679581782
transform 1 0 83424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_870
timestamp 1679581782
transform 1 0 84096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_877
timestamp 1679581782
transform 1 0 84768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_884
timestamp 1679581782
transform 1 0 85440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_891
timestamp 1679581782
transform 1 0 86112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_898
timestamp 1679581782
transform 1 0 86784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_905
timestamp 1679581782
transform 1 0 87456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_912
timestamp 1679581782
transform 1 0 88128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_919
timestamp 1679581782
transform 1 0 88800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_926
timestamp 1679581782
transform 1 0 89472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_933
timestamp 1679581782
transform 1 0 90144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_940
timestamp 1679581782
transform 1 0 90816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_947
timestamp 1679581782
transform 1 0 91488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_954
timestamp 1679581782
transform 1 0 92160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_961
timestamp 1679581782
transform 1 0 92832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_968
timestamp 1679581782
transform 1 0 93504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_975
timestamp 1679581782
transform 1 0 94176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_982
timestamp 1679581782
transform 1 0 94848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_989
timestamp 1679581782
transform 1 0 95520 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_996
timestamp 1677579658
transform 1 0 96192 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_1022
timestamp 1679581782
transform 1 0 98688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_11
timestamp 1677580104
transform 1 0 1632 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_13
timestamp 1677579658
transform 1 0 1824 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_51
timestamp 1679577901
transform 1 0 5472 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_55
timestamp 1677579658
transform 1 0 5856 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_765
timestamp 1679581782
transform 1 0 74016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_772
timestamp 1679581782
transform 1 0 74688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_779
timestamp 1679581782
transform 1 0 75360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_786
timestamp 1679581782
transform 1 0 76032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_793
timestamp 1679581782
transform 1 0 76704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_800
timestamp 1679581782
transform 1 0 77376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_807
timestamp 1679581782
transform 1 0 78048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_814
timestamp 1679581782
transform 1 0 78720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_821
timestamp 1679581782
transform 1 0 79392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_828
timestamp 1679581782
transform 1 0 80064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_835
timestamp 1679581782
transform 1 0 80736 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_842
timestamp 1677579658
transform 1 0 81408 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_853
timestamp 1679581782
transform 1 0 82464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_860
timestamp 1679581782
transform 1 0 83136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_867
timestamp 1679581782
transform 1 0 83808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_874
timestamp 1679581782
transform 1 0 84480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_881
timestamp 1679581782
transform 1 0 85152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_888
timestamp 1679581782
transform 1 0 85824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_895
timestamp 1679581782
transform 1 0 86496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_902
timestamp 1679581782
transform 1 0 87168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_909
timestamp 1679581782
transform 1 0 87840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_916
timestamp 1679581782
transform 1 0 88512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_923
timestamp 1679581782
transform 1 0 89184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_930
timestamp 1679581782
transform 1 0 89856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_937
timestamp 1679581782
transform 1 0 90528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_944
timestamp 1679581782
transform 1 0 91200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_951
timestamp 1679581782
transform 1 0 91872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_958
timestamp 1679581782
transform 1 0 92544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_965
timestamp 1679581782
transform 1 0 93216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_972
timestamp 1679581782
transform 1 0 93888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_979
timestamp 1679581782
transform 1 0 94560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_986
timestamp 1679581782
transform 1 0 95232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_993
timestamp 1679581782
transform 1 0 95904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1000
timestamp 1679581782
transform 1 0 96576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1007
timestamp 1679581782
transform 1 0 97248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1014
timestamp 1679581782
transform 1 0 97920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1021
timestamp 1679581782
transform 1 0 98592 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_1028
timestamp 1677579658
transform 1 0 99264 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_28
timestamp 1677579658
transform 1 0 3264 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_765
timestamp 1679581782
transform 1 0 74016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_772
timestamp 1679581782
transform 1 0 74688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_779
timestamp 1679581782
transform 1 0 75360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_786
timestamp 1679581782
transform 1 0 76032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_793
timestamp 1679581782
transform 1 0 76704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_800
timestamp 1679581782
transform 1 0 77376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_807
timestamp 1679581782
transform 1 0 78048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_814
timestamp 1679581782
transform 1 0 78720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_821
timestamp 1679581782
transform 1 0 79392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_828
timestamp 1679581782
transform 1 0 80064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_835
timestamp 1679581782
transform 1 0 80736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_842
timestamp 1679581782
transform 1 0 81408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_849
timestamp 1679577901
transform 1 0 82080 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_853
timestamp 1677580104
transform 1 0 82464 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_882
timestamp 1679581782
transform 1 0 85248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_889
timestamp 1679581782
transform 1 0 85920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_896
timestamp 1679581782
transform 1 0 86592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_903
timestamp 1679581782
transform 1 0 87264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_910
timestamp 1679581782
transform 1 0 87936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_917
timestamp 1679581782
transform 1 0 88608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_924
timestamp 1679581782
transform 1 0 89280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_931
timestamp 1679581782
transform 1 0 89952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_938
timestamp 1679581782
transform 1 0 90624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_945
timestamp 1679581782
transform 1 0 91296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_952
timestamp 1679581782
transform 1 0 91968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_959
timestamp 1679581782
transform 1 0 92640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_966
timestamp 1679581782
transform 1 0 93312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_973
timestamp 1679581782
transform 1 0 93984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_980
timestamp 1679581782
transform 1 0 94656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_987
timestamp 1679581782
transform 1 0 95328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_994
timestamp 1679581782
transform 1 0 96000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1001
timestamp 1679581782
transform 1 0 96672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1008
timestamp 1679581782
transform 1 0 97344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1015
timestamp 1679581782
transform 1 0 98016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1022
timestamp 1679581782
transform 1 0 98688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_25
timestamp 1679577901
transform 1 0 2976 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_29
timestamp 1677580104
transform 1 0 3360 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_41
timestamp 1679581782
transform 1 0 4512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_48
timestamp 1679581782
transform 1 0 5184 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_55
timestamp 1677579658
transform 1 0 5856 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_765
timestamp 1679581782
transform 1 0 74016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_772
timestamp 1679581782
transform 1 0 74688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_779
timestamp 1679581782
transform 1 0 75360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_786
timestamp 1679581782
transform 1 0 76032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_793
timestamp 1679581782
transform 1 0 76704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_800
timestamp 1679581782
transform 1 0 77376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_807
timestamp 1679581782
transform 1 0 78048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_814
timestamp 1679581782
transform 1 0 78720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_821
timestamp 1679581782
transform 1 0 79392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_828
timestamp 1679581782
transform 1 0 80064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_835
timestamp 1679581782
transform 1 0 80736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_842
timestamp 1679581782
transform 1 0 81408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_849
timestamp 1679581782
transform 1 0 82080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_856
timestamp 1679577901
transform 1 0 82752 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_860
timestamp 1677580104
transform 1 0 83136 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_4
timestamp 1679581782
transform 1 0 960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_11
timestamp 1679581782
transform 1 0 1632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_18
timestamp 1679581782
transform 1 0 2304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_25
timestamp 1679577901
transform 1 0 2976 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_778
timestamp 1679581782
transform 1 0 75264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_785
timestamp 1679581782
transform 1 0 75936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_792
timestamp 1679581782
transform 1 0 76608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_799
timestamp 1679581782
transform 1 0 77280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_806
timestamp 1679581782
transform 1 0 77952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_813
timestamp 1679581782
transform 1 0 78624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_820
timestamp 1679581782
transform 1 0 79296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_827
timestamp 1679581782
transform 1 0 79968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_834
timestamp 1679581782
transform 1 0 80640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_841
timestamp 1679581782
transform 1 0 81312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_848
timestamp 1679581782
transform 1 0 81984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_855
timestamp 1679581782
transform 1 0 82656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_4
timestamp 1679581782
transform 1 0 960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_11
timestamp 1679581782
transform 1 0 1632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_18
timestamp 1679581782
transform 1 0 2304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_25
timestamp 1679581782
transform 1 0 2976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_32
timestamp 1679581782
transform 1 0 3648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_39
timestamp 1679581782
transform 1 0 4320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_46
timestamp 1679581782
transform 1 0 4992 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_53
timestamp 1677580104
transform 1 0 5664 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_55
timestamp 1677579658
transform 1 0 5856 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_778
timestamp 1679581782
transform 1 0 75264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_785
timestamp 1679581782
transform 1 0 75936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_792
timestamp 1679581782
transform 1 0 76608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_799
timestamp 1679581782
transform 1 0 77280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_806
timestamp 1679581782
transform 1 0 77952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_813
timestamp 1679581782
transform 1 0 78624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_820
timestamp 1679581782
transform 1 0 79296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_827
timestamp 1679581782
transform 1 0 79968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_834
timestamp 1679581782
transform 1 0 80640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_841
timestamp 1679581782
transform 1 0 81312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_848
timestamp 1679581782
transform 1 0 81984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_855
timestamp 1679581782
transform 1 0 82656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_4
timestamp 1679581782
transform 1 0 960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_11
timestamp 1679581782
transform 1 0 1632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_18
timestamp 1679581782
transform 1 0 2304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_25
timestamp 1679581782
transform 1 0 2976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_32
timestamp 1679577901
transform 1 0 3648 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_36
timestamp 1677580104
transform 1 0 4032 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_48
timestamp 1679581782
transform 1 0 5184 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_55
timestamp 1677579658
transform 1 0 5856 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_768
timestamp 1679581782
transform 1 0 74304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_775
timestamp 1679581782
transform 1 0 74976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_782
timestamp 1679581782
transform 1 0 75648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_789
timestamp 1679581782
transform 1 0 76320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_796
timestamp 1679581782
transform 1 0 76992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_803
timestamp 1679581782
transform 1 0 77664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_810
timestamp 1679581782
transform 1 0 78336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_817
timestamp 1679581782
transform 1 0 79008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_824
timestamp 1679581782
transform 1 0 79680 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_831
timestamp 1677579658
transform 1 0 80352 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_859
timestamp 1677580104
transform 1 0 83040 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_861
timestamp 1677579658
transform 1 0 83232 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_11
timestamp 1679581782
transform 1 0 1632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_18
timestamp 1679581782
transform 1 0 2304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_25
timestamp 1679577901
transform 1 0 2976 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_765
timestamp 1679581782
transform 1 0 74016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_772
timestamp 1679581782
transform 1 0 74688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_779
timestamp 1679581782
transform 1 0 75360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_786
timestamp 1679581782
transform 1 0 76032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_793
timestamp 1679581782
transform 1 0 76704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_800
timestamp 1679581782
transform 1 0 77376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_807
timestamp 1679581782
transform 1 0 78048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_814
timestamp 1679581782
transform 1 0 78720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_821
timestamp 1679577901
transform 1 0 79392 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679581782
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679581782
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679581782
transform 1 0 1920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679581782
transform 1 0 2592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_28
timestamp 1679581782
transform 1 0 3264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_35
timestamp 1679581782
transform 1 0 3936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_42
timestamp 1679581782
transform 1 0 4608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_49
timestamp 1679581782
transform 1 0 5280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_765
timestamp 1679581782
transform 1 0 74016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_772
timestamp 1679581782
transform 1 0 74688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_779
timestamp 1679581782
transform 1 0 75360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_786
timestamp 1679581782
transform 1 0 76032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_793
timestamp 1679581782
transform 1 0 76704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_800
timestamp 1679581782
transform 1 0 77376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_807
timestamp 1679581782
transform 1 0 78048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_814
timestamp 1679581782
transform 1 0 78720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_821
timestamp 1679581782
transform 1 0 79392 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_838
timestamp 1677579658
transform 1 0 81024 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_849
timestamp 1679581782
transform 1 0 82080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_856
timestamp 1679577901
transform 1 0 82752 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_860
timestamp 1677580104
transform 1 0 83136 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_35
timestamp 1679577901
transform 1 0 3936 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_765
timestamp 1679581782
transform 1 0 74016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_772
timestamp 1679581782
transform 1 0 74688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_779
timestamp 1679581782
transform 1 0 75360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_786
timestamp 1679581782
transform 1 0 76032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_793
timestamp 1679581782
transform 1 0 76704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_800
timestamp 1679581782
transform 1 0 77376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_807
timestamp 1679581782
transform 1 0 78048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_814
timestamp 1679581782
transform 1 0 78720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_821
timestamp 1679581782
transform 1 0 79392 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_828
timestamp 1677580104
transform 1 0 80064 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_830
timestamp 1677579658
transform 1 0 80256 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_858
timestamp 1679577901
transform 1 0 82944 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_28
timestamp 1677579658
transform 1 0 3264 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_765
timestamp 1679581782
transform 1 0 74016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_772
timestamp 1679581782
transform 1 0 74688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_779
timestamp 1679581782
transform 1 0 75360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_786
timestamp 1679581782
transform 1 0 76032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_793
timestamp 1679581782
transform 1 0 76704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_800
timestamp 1679581782
transform 1 0 77376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_807
timestamp 1679581782
transform 1 0 78048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_814
timestamp 1679581782
transform 1 0 78720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_821
timestamp 1679581782
transform 1 0 79392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_828
timestamp 1679581782
transform 1 0 80064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_790
timestamp 1679581782
transform 1 0 76416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_797
timestamp 1679581782
transform 1 0 77088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_804
timestamp 1679581782
transform 1 0 77760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_811
timestamp 1679581782
transform 1 0 78432 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_818
timestamp 1677579658
transform 1 0 79104 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_856
timestamp 1679577901
transform 1 0 82752 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_860
timestamp 1677580104
transform 1 0 83136 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_765
timestamp 1679581782
transform 1 0 74016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_772
timestamp 1679581782
transform 1 0 74688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_779
timestamp 1679581782
transform 1 0 75360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_786
timestamp 1679581782
transform 1 0 76032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_793
timestamp 1679581782
transform 1 0 76704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_800
timestamp 1679581782
transform 1 0 77376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_807
timestamp 1679581782
transform 1 0 78048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_814
timestamp 1679581782
transform 1 0 78720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_821
timestamp 1679577901
transform 1 0 79392 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_825
timestamp 1677579658
transform 1 0 79776 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_846
timestamp 1679581782
transform 1 0 81792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_853
timestamp 1679581782
transform 1 0 82464 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_860
timestamp 1677580104
transform 1 0 83136 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_765
timestamp 1679581782
transform 1 0 74016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_772
timestamp 1679581782
transform 1 0 74688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_779
timestamp 1679581782
transform 1 0 75360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_786
timestamp 1679581782
transform 1 0 76032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_793
timestamp 1679581782
transform 1 0 76704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_800
timestamp 1679581782
transform 1 0 77376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_807
timestamp 1679581782
transform 1 0 78048 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_814
timestamp 1677580104
transform 1 0 78720 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_816
timestamp 1677579658
transform 1 0 78912 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_854
timestamp 1679581782
transform 1 0 82560 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_861
timestamp 1677579658
transform 1 0 83232 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_35
timestamp 1679577901
transform 1 0 3936 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_765
timestamp 1679581782
transform 1 0 74016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_772
timestamp 1679581782
transform 1 0 74688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_779
timestamp 1679581782
transform 1 0 75360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_786
timestamp 1679581782
transform 1 0 76032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_793
timestamp 1679581782
transform 1 0 76704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_800
timestamp 1679581782
transform 1 0 77376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_807
timestamp 1679581782
transform 1 0 78048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_814
timestamp 1679581782
transform 1 0 78720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_821
timestamp 1679577901
transform 1 0 79392 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_825
timestamp 1677579658
transform 1 0 79776 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_830
timestamp 1679577901
transform 1 0 80256 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_834
timestamp 1677579658
transform 1 0 80640 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_28
timestamp 1677579658
transform 1 0 3264 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_765
timestamp 1679581782
transform 1 0 74016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_772
timestamp 1679581782
transform 1 0 74688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_779
timestamp 1679581782
transform 1 0 75360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_786
timestamp 1679581782
transform 1 0 76032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_793
timestamp 1679581782
transform 1 0 76704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_800
timestamp 1679581782
transform 1 0 77376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_807
timestamp 1679581782
transform 1 0 78048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_814
timestamp 1679581782
transform 1 0 78720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_821
timestamp 1679581782
transform 1 0 79392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_828
timestamp 1679577901
transform 1 0 80064 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_832
timestamp 1677579658
transform 1 0 80448 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_843
timestamp 1677579658
transform 1 0 81504 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_848
timestamp 1679581782
transform 1 0 81984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_855
timestamp 1679581782
transform 1 0 82656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_35
timestamp 1679577901
transform 1 0 3936 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_765
timestamp 1679581782
transform 1 0 74016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_772
timestamp 1679581782
transform 1 0 74688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_779
timestamp 1679581782
transform 1 0 75360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_786
timestamp 1679581782
transform 1 0 76032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_793
timestamp 1679581782
transform 1 0 76704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_800
timestamp 1679581782
transform 1 0 77376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_807
timestamp 1679581782
transform 1 0 78048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_814
timestamp 1679581782
transform 1 0 78720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_821
timestamp 1679581782
transform 1 0 79392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_828
timestamp 1679581782
transform 1 0 80064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_49
timestamp 1677579658
transform 1 0 5280 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_54
timestamp 1677580104
transform 1 0 5760 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_765
timestamp 1679581782
transform 1 0 74016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_772
timestamp 1679581782
transform 1 0 74688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_779
timestamp 1679581782
transform 1 0 75360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_786
timestamp 1679581782
transform 1 0 76032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_793
timestamp 1679581782
transform 1 0 76704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_800
timestamp 1679581782
transform 1 0 77376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_807
timestamp 1679581782
transform 1 0 78048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_814
timestamp 1679581782
transform 1 0 78720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_821
timestamp 1679581782
transform 1 0 79392 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_828
timestamp 1677580104
transform 1 0 80064 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_830
timestamp 1677579658
transform 1 0 80256 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_765
timestamp 1679581782
transform 1 0 74016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_772
timestamp 1679581782
transform 1 0 74688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_779
timestamp 1679581782
transform 1 0 75360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_786
timestamp 1679581782
transform 1 0 76032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_793
timestamp 1679581782
transform 1 0 76704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_800
timestamp 1679581782
transform 1 0 77376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_807
timestamp 1679581782
transform 1 0 78048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_814
timestamp 1679581782
transform 1 0 78720 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_821
timestamp 1677580104
transform 1 0 79392 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_843
timestamp 1677580104
transform 1 0 81504 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_849
timestamp 1679581782
transform 1 0 82080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_856
timestamp 1679577901
transform 1 0 82752 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_860
timestamp 1677580104
transform 1 0 83136 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_63
timestamp 1679577901
transform 1 0 6624 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_67
timestamp 1677579658
transform 1 0 7008 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_81
timestamp 1679581782
transform 1 0 8352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_88
timestamp 1679581782
transform 1 0 9024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_95
timestamp 1679581782
transform 1 0 9696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_102
timestamp 1679577901
transform 1 0 10368 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_143
timestamp 1679581782
transform 1 0 14304 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_150
timestamp 1677580104
transform 1 0 14976 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_192
timestamp 1679581782
transform 1 0 19008 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_239
timestamp 1677579658
transform 1 0 23520 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_277
timestamp 1679581782
transform 1 0 27168 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_284
timestamp 1677579658
transform 1 0 27840 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_312
timestamp 1679577901
transform 1 0 30528 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_316
timestamp 1677580104
transform 1 0 30912 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_365
timestamp 1679581782
transform 1 0 35616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_372
timestamp 1679581782
transform 1 0 36288 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_379
timestamp 1677580104
transform 1 0 36960 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_381
timestamp 1677579658
transform 1 0 37152 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_409
timestamp 1679581782
transform 1 0 39840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_416
timestamp 1679577901
transform 1 0 40512 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_420
timestamp 1677579658
transform 1 0 40896 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_426
timestamp 1677579658
transform 1 0 41472 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_431
timestamp 1677580104
transform 1 0 41952 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_436
timestamp 1677580104
transform 1 0 42432 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_467
timestamp 1679581782
transform 1 0 45408 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_474
timestamp 1677580104
transform 1 0 46080 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_476
timestamp 1677579658
transform 1 0 46272 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_524
timestamp 1679577901
transform 1 0 50880 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_554
timestamp 1677580104
transform 1 0 53760 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_556
timestamp 1677579658
transform 1 0 53952 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_584
timestamp 1679581782
transform 1 0 56640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_591
timestamp 1679581782
transform 1 0 57312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_598
timestamp 1679581782
transform 1 0 57984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_605
timestamp 1679581782
transform 1 0 58656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_612
timestamp 1679581782
transform 1 0 59328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_619
timestamp 1679581782
transform 1 0 60000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_626
timestamp 1679581782
transform 1 0 60672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_671
timestamp 1679581782
transform 1 0 64992 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_678
timestamp 1677579658
transform 1 0 65664 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_692
timestamp 1679581782
transform 1 0 67008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_699
timestamp 1679581782
transform 1 0 67680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_706
timestamp 1679581782
transform 1 0 68352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_713
timestamp 1679581782
transform 1 0 69024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_720
timestamp 1679581782
transform 1 0 69696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_727
timestamp 1679581782
transform 1 0 70368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_734
timestamp 1679581782
transform 1 0 71040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_741
timestamp 1679581782
transform 1 0 71712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_748
timestamp 1679581782
transform 1 0 72384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_755
timestamp 1679581782
transform 1 0 73056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_762
timestamp 1679581782
transform 1 0 73728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_769
timestamp 1679581782
transform 1 0 74400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_776
timestamp 1679581782
transform 1 0 75072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_783
timestamp 1679581782
transform 1 0 75744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_790
timestamp 1679581782
transform 1 0 76416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_797
timestamp 1679581782
transform 1 0 77088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_804
timestamp 1679581782
transform 1 0 77760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_811
timestamp 1679581782
transform 1 0 78432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_818
timestamp 1679581782
transform 1 0 79104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_825
timestamp 1679581782
transform 1 0 79776 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_832
timestamp 1677580104
transform 1 0 80448 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_834
timestamp 1677579658
transform 1 0 80640 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_119
timestamp 1677580104
transform 1 0 12000 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_125
timestamp 1679581782
transform 1 0 12576 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_182
timestamp 1677579658
transform 1 0 18048 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_220
timestamp 1679581782
transform 1 0 21696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_227
timestamp 1679581782
transform 1 0 22368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_234
timestamp 1679581782
transform 1 0 23040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_241
timestamp 1679577901
transform 1 0 23712 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_245
timestamp 1677579658
transform 1 0 24096 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_331
timestamp 1679581782
transform 1 0 32352 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_338
timestamp 1677580104
transform 1 0 33024 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_340
timestamp 1677579658
transform 1 0 33216 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_381
timestamp 1677580104
transform 1 0 37152 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_413
timestamp 1677579658
transform 1 0 40224 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_445
timestamp 1677579658
transform 1 0 43296 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_451
timestamp 1677579658
transform 1 0 43872 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_574
timestamp 1679581782
transform 1 0 55680 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_581
timestamp 1679581782
transform 1 0 56352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_588
timestamp 1679581782
transform 1 0 57024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_595
timestamp 1679581782
transform 1 0 57696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_602
timestamp 1679581782
transform 1 0 58368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_609
timestamp 1679581782
transform 1 0 59040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_616
timestamp 1679581782
transform 1 0 59712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679581782
transform 1 0 60384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_630
timestamp 1679581782
transform 1 0 61056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_637
timestamp 1679581782
transform 1 0 61728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_644
timestamp 1679581782
transform 1 0 62400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_651
timestamp 1679581782
transform 1 0 63072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_658
timestamp 1679581782
transform 1 0 63744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_665
timestamp 1679581782
transform 1 0 64416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_672
timestamp 1679581782
transform 1 0 65088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_679
timestamp 1679581782
transform 1 0 65760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_686
timestamp 1679581782
transform 1 0 66432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_693
timestamp 1679581782
transform 1 0 67104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_700
timestamp 1679581782
transform 1 0 67776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_707
timestamp 1679581782
transform 1 0 68448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_714
timestamp 1679581782
transform 1 0 69120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_721
timestamp 1679581782
transform 1 0 69792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_728
timestamp 1679581782
transform 1 0 70464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_735
timestamp 1679581782
transform 1 0 71136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_742
timestamp 1679581782
transform 1 0 71808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_749
timestamp 1679581782
transform 1 0 72480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_756
timestamp 1679581782
transform 1 0 73152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_763
timestamp 1679581782
transform 1 0 73824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_770
timestamp 1679581782
transform 1 0 74496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_777
timestamp 1679581782
transform 1 0 75168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_784
timestamp 1679581782
transform 1 0 75840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_791
timestamp 1679581782
transform 1 0 76512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_798
timestamp 1679581782
transform 1 0 77184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_805
timestamp 1679581782
transform 1 0 77856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_812
timestamp 1679581782
transform 1 0 78528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_819
timestamp 1679581782
transform 1 0 79200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_826
timestamp 1679581782
transform 1 0 79872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_833
timestamp 1679581782
transform 1 0 80544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_840
timestamp 1679581782
transform 1 0 81216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_847
timestamp 1679581782
transform 1 0 81888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_854
timestamp 1679581782
transform 1 0 82560 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_861
timestamp 1677579658
transform 1 0 83232 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_133
timestamp 1677580104
transform 1 0 13344 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_135
timestamp 1677579658
transform 1 0 13536 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_150
timestamp 1677580104
transform 1 0 14976 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_179
timestamp 1679581782
transform 1 0 17760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_186
timestamp 1679577901
transform 1 0 18432 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_197
timestamp 1677579658
transform 1 0 19488 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_216
timestamp 1677580104
transform 1 0 21312 0 1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_46_223
timestamp 1679577901
transform 1 0 21984 0 1 35532
box -48 -56 432 834
use sg13g2_decap_4  FILLER_46_254
timestamp 1679577901
transform 1 0 24960 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_258
timestamp 1677580104
transform 1 0 25344 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_315
timestamp 1677580104
transform 1 0 30816 0 1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_46_356
timestamp 1679577901
transform 1 0 34752 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_360
timestamp 1677580104
transform 1 0 35136 0 1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_46_389
timestamp 1679577901
transform 1 0 37920 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_403
timestamp 1677579658
transform 1 0 39264 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_414
timestamp 1679581782
transform 1 0 40320 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_421
timestamp 1677580104
transform 1 0 40992 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_423
timestamp 1677579658
transform 1 0 41184 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_438
timestamp 1679581782
transform 1 0 42624 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_445
timestamp 1677579658
transform 1 0 43296 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_46_483
timestamp 1679577901
transform 1 0 46944 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_487
timestamp 1677579658
transform 1 0 47328 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_513
timestamp 1679581782
transform 1 0 49824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_520
timestamp 1679581782
transform 1 0 50496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_527
timestamp 1679581782
transform 1 0 51168 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_534
timestamp 1677580104
transform 1 0 51840 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_536
timestamp 1677579658
transform 1 0 52032 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_557
timestamp 1679581782
transform 1 0 54048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_564
timestamp 1679581782
transform 1 0 54720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_571
timestamp 1679581782
transform 1 0 55392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_578
timestamp 1679581782
transform 1 0 56064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_585
timestamp 1679581782
transform 1 0 56736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_592
timestamp 1679581782
transform 1 0 57408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_599
timestamp 1679581782
transform 1 0 58080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_606
timestamp 1679581782
transform 1 0 58752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_613
timestamp 1679581782
transform 1 0 59424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_620
timestamp 1679581782
transform 1 0 60096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_627
timestamp 1679581782
transform 1 0 60768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_634
timestamp 1679581782
transform 1 0 61440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_641
timestamp 1679581782
transform 1 0 62112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_648
timestamp 1679581782
transform 1 0 62784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_655
timestamp 1679581782
transform 1 0 63456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_662
timestamp 1679581782
transform 1 0 64128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_669
timestamp 1679581782
transform 1 0 64800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_676
timestamp 1679581782
transform 1 0 65472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_683
timestamp 1679581782
transform 1 0 66144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_690
timestamp 1679581782
transform 1 0 66816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_697
timestamp 1679581782
transform 1 0 67488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_704
timestamp 1679581782
transform 1 0 68160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_711
timestamp 1679581782
transform 1 0 68832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_718
timestamp 1679581782
transform 1 0 69504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_725
timestamp 1679581782
transform 1 0 70176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_732
timestamp 1679581782
transform 1 0 70848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_739
timestamp 1679577901
transform 1 0 71520 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_743
timestamp 1677579658
transform 1 0 71904 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_757
timestamp 1679581782
transform 1 0 73248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_764
timestamp 1679581782
transform 1 0 73920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_771
timestamp 1679581782
transform 1 0 74592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_778
timestamp 1679581782
transform 1 0 75264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_785
timestamp 1679581782
transform 1 0 75936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_792
timestamp 1679581782
transform 1 0 76608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_799
timestamp 1679581782
transform 1 0 77280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_806
timestamp 1679581782
transform 1 0 77952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_813
timestamp 1679581782
transform 1 0 78624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_820
timestamp 1679581782
transform 1 0 79296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_827
timestamp 1679581782
transform 1 0 79968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_834
timestamp 1679581782
transform 1 0 80640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_841
timestamp 1679581782
transform 1 0 81312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_848
timestamp 1679581782
transform 1 0 81984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_855
timestamp 1679581782
transform 1 0 82656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_175
timestamp 1679577901
transform 1 0 17376 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_214
timestamp 1677579658
transform 1 0 21120 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_222
timestamp 1677579658
transform 1 0 21888 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_231
timestamp 1677579658
transform 1 0 22752 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_245
timestamp 1677580104
transform 1 0 24096 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_252
timestamp 1677580104
transform 1 0 24768 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_261
timestamp 1677580104
transform 1 0 25632 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_286
timestamp 1679581782
transform 1 0 28032 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_293
timestamp 1677580104
transform 1 0 28704 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_295
timestamp 1677579658
transform 1 0 28896 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_323
timestamp 1679581782
transform 1 0 31584 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_330
timestamp 1677579658
transform 1 0 32256 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_368
timestamp 1679581782
transform 1 0 35904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_375
timestamp 1679581782
transform 1 0 36576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_382
timestamp 1679581782
transform 1 0 37248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_389
timestamp 1679577901
transform 1 0 37920 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_393
timestamp 1677579658
transform 1 0 38304 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_455
timestamp 1679577901
transform 1 0 44256 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_459
timestamp 1677580104
transform 1 0 44640 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679581782
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679581782
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679581782
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_861
timestamp 1677579658
transform 1 0 83232 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_189
timestamp 1679577901
transform 1 0 18720 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_193
timestamp 1677579658
transform 1 0 19104 0 1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_48_199
timestamp 1679577901
transform 1 0 19680 0 1 37044
box -48 -56 432 834
use sg13g2_decap_4  FILLER_48_257
timestamp 1679577901
transform 1 0 25248 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_261
timestamp 1677580104
transform 1 0 25632 0 1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_294
timestamp 1677580104
transform 1 0 28800 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_296
timestamp 1677579658
transform 1 0 28992 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_332
timestamp 1679581782
transform 1 0 32448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_339
timestamp 1679581782
transform 1 0 33120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_346
timestamp 1679581782
transform 1 0 33792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_353
timestamp 1679581782
transform 1 0 34464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_360
timestamp 1679581782
transform 1 0 35136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_367
timestamp 1679581782
transform 1 0 35808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_374
timestamp 1679581782
transform 1 0 36480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_381
timestamp 1679577901
transform 1 0 37152 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_385
timestamp 1677580104
transform 1 0 37536 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_414
timestamp 1679581782
transform 1 0 40320 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_421
timestamp 1677579658
transform 1 0 40992 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_459
timestamp 1679581782
transform 1 0 44640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_466
timestamp 1679581782
transform 1 0 45312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_473
timestamp 1679581782
transform 1 0 45984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_480
timestamp 1679581782
transform 1 0 46656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_487
timestamp 1679581782
transform 1 0 47328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_494
timestamp 1679581782
transform 1 0 48000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_501
timestamp 1679581782
transform 1 0 48672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_508
timestamp 1679581782
transform 1 0 49344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_515
timestamp 1679581782
transform 1 0 50016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_522
timestamp 1679581782
transform 1 0 50688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_529
timestamp 1679581782
transform 1 0 51360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_536
timestamp 1679581782
transform 1 0 52032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_543
timestamp 1679581782
transform 1 0 52704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_550
timestamp 1679581782
transform 1 0 53376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_557
timestamp 1679581782
transform 1 0 54048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_564
timestamp 1679581782
transform 1 0 54720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_571
timestamp 1679581782
transform 1 0 55392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_578
timestamp 1679581782
transform 1 0 56064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_585
timestamp 1679581782
transform 1 0 56736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_592
timestamp 1679581782
transform 1 0 57408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_599
timestamp 1679581782
transform 1 0 58080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_606
timestamp 1679581782
transform 1 0 58752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_613
timestamp 1679581782
transform 1 0 59424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_620
timestamp 1679581782
transform 1 0 60096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_627
timestamp 1679581782
transform 1 0 60768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_634
timestamp 1679581782
transform 1 0 61440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_641
timestamp 1679581782
transform 1 0 62112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_648
timestamp 1679581782
transform 1 0 62784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_655
timestamp 1679581782
transform 1 0 63456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_662
timestamp 1679581782
transform 1 0 64128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_669
timestamp 1679581782
transform 1 0 64800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_676
timestamp 1679581782
transform 1 0 65472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_683
timestamp 1679581782
transform 1 0 66144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_690
timestamp 1679581782
transform 1 0 66816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_697
timestamp 1679581782
transform 1 0 67488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_704
timestamp 1679581782
transform 1 0 68160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_711
timestamp 1679581782
transform 1 0 68832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_718
timestamp 1679581782
transform 1 0 69504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_725
timestamp 1679581782
transform 1 0 70176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_732
timestamp 1679581782
transform 1 0 70848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_739
timestamp 1679581782
transform 1 0 71520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_746
timestamp 1679581782
transform 1 0 72192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_753
timestamp 1679581782
transform 1 0 72864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_760
timestamp 1679581782
transform 1 0 73536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_767
timestamp 1679581782
transform 1 0 74208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_774
timestamp 1679581782
transform 1 0 74880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_781
timestamp 1679581782
transform 1 0 75552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_788
timestamp 1679581782
transform 1 0 76224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_795
timestamp 1679581782
transform 1 0 76896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_802
timestamp 1679581782
transform 1 0 77568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_809
timestamp 1679581782
transform 1 0 78240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_816
timestamp 1679581782
transform 1 0 78912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_823
timestamp 1679581782
transform 1 0 79584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_830
timestamp 1679581782
transform 1 0 80256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_837
timestamp 1679581782
transform 1 0 80928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_844
timestamp 1679581782
transform 1 0 81600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_851
timestamp 1679581782
transform 1 0 82272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_858
timestamp 1679577901
transform 1 0 82944 0 1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679581782
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679581782
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679581782
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679581782
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679581782
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679581782
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679581782
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679581782
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679581782
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679581782
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679581782
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679581782
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_207
timestamp 1679577901
transform 1 0 20448 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_211
timestamp 1677579658
transform 1 0 20832 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_217
timestamp 1677580104
transform 1 0 21408 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_219
timestamp 1677579658
transform 1 0 21600 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679581782
transform 1 0 22080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_231
timestamp 1679577901
transform 1 0 22752 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_247
timestamp 1679581782
transform 1 0 24288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_254
timestamp 1679581782
transform 1 0 24960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_261
timestamp 1679581782
transform 1 0 25632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_268
timestamp 1679577901
transform 1 0 26304 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_272
timestamp 1677579658
transform 1 0 26688 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_279
timestamp 1679581782
transform 1 0 27360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_286
timestamp 1679577901
transform 1 0 28032 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_302
timestamp 1679581782
transform 1 0 29568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_309
timestamp 1679581782
transform 1 0 30240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_316
timestamp 1679581782
transform 1 0 30912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_323
timestamp 1679581782
transform 1 0 31584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_330
timestamp 1679581782
transform 1 0 32256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_337
timestamp 1679581782
transform 1 0 32928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_344
timestamp 1679581782
transform 1 0 33600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_351
timestamp 1679581782
transform 1 0 34272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_358
timestamp 1679581782
transform 1 0 34944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_365
timestamp 1679581782
transform 1 0 35616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_372
timestamp 1679581782
transform 1 0 36288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_379
timestamp 1679581782
transform 1 0 36960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_386
timestamp 1679581782
transform 1 0 37632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679581782
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679581782
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_417
timestamp 1677580104
transform 1 0 40608 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_419
timestamp 1677579658
transform 1 0 40800 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_430
timestamp 1679581782
transform 1 0 41856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_437
timestamp 1679581782
transform 1 0 42528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_444
timestamp 1679581782
transform 1 0 43200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_451
timestamp 1679581782
transform 1 0 43872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_458
timestamp 1679581782
transform 1 0 44544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_465
timestamp 1679581782
transform 1 0 45216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_472
timestamp 1679581782
transform 1 0 45888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_479
timestamp 1679581782
transform 1 0 46560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_486
timestamp 1679581782
transform 1 0 47232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_493
timestamp 1679581782
transform 1 0 47904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_500
timestamp 1679581782
transform 1 0 48576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_507
timestamp 1679581782
transform 1 0 49248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_514
timestamp 1679581782
transform 1 0 49920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_521
timestamp 1679581782
transform 1 0 50592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_528
timestamp 1679581782
transform 1 0 51264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_535
timestamp 1679581782
transform 1 0 51936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_542
timestamp 1679581782
transform 1 0 52608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_549
timestamp 1679581782
transform 1 0 53280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_556
timestamp 1679581782
transform 1 0 53952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_563
timestamp 1679581782
transform 1 0 54624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_570
timestamp 1679581782
transform 1 0 55296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_577
timestamp 1679581782
transform 1 0 55968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_584
timestamp 1679581782
transform 1 0 56640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_591
timestamp 1679581782
transform 1 0 57312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_598
timestamp 1679581782
transform 1 0 57984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_605
timestamp 1679581782
transform 1 0 58656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_612
timestamp 1679581782
transform 1 0 59328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_619
timestamp 1679581782
transform 1 0 60000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_626
timestamp 1679581782
transform 1 0 60672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_633
timestamp 1679581782
transform 1 0 61344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_640
timestamp 1679581782
transform 1 0 62016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_647
timestamp 1679581782
transform 1 0 62688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_654
timestamp 1679581782
transform 1 0 63360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_661
timestamp 1679581782
transform 1 0 64032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_668
timestamp 1679581782
transform 1 0 64704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_675
timestamp 1679581782
transform 1 0 65376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_682
timestamp 1679581782
transform 1 0 66048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_689
timestamp 1679581782
transform 1 0 66720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_696
timestamp 1679581782
transform 1 0 67392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_703
timestamp 1679581782
transform 1 0 68064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_710
timestamp 1679581782
transform 1 0 68736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_717
timestamp 1679581782
transform 1 0 69408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_737
timestamp 1679581782
transform 1 0 71328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_744
timestamp 1679581782
transform 1 0 72000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_751
timestamp 1679581782
transform 1 0 72672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_758
timestamp 1679581782
transform 1 0 73344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_765
timestamp 1679581782
transform 1 0 74016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_772
timestamp 1679581782
transform 1 0 74688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_779
timestamp 1679581782
transform 1 0 75360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_786
timestamp 1679581782
transform 1 0 76032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_793
timestamp 1679581782
transform 1 0 76704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_800
timestamp 1679581782
transform 1 0 77376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_807
timestamp 1679581782
transform 1 0 78048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_814
timestamp 1679581782
transform 1 0 78720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_821
timestamp 1679581782
transform 1 0 79392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_828
timestamp 1679581782
transform 1 0 80064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_835
timestamp 1679581782
transform 1 0 80736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_842
timestamp 1679581782
transform 1 0 81408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_849
timestamp 1679581782
transform 1 0 82080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_856
timestamp 1679577901
transform 1 0 82752 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_860
timestamp 1677580104
transform 1 0 83136 0 -1 38556
box -48 -56 240 834
use sg13g2_tielo  heichips25_internal_47
timestamp 1680000637
transform 1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_48
timestamp 1680000637
transform 1 0 576 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_49
timestamp 1680000637
transform 1 0 576 0 -1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_50
timestamp 1680000637
transform 1 0 576 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_51
timestamp 1680000637
transform 1 0 576 0 -1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_52
timestamp 1680000637
transform 1 0 576 0 1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_53
timestamp 1680000637
transform 1 0 576 0 1 21924
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal
timestamp 1680000637
transform 1 0 576 0 1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_54
timestamp 1680000637
transform 1 0 576 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_55
timestamp 1680000637
transform 1 0 576 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_56
timestamp 1680000637
transform 1 0 576 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_57
timestamp 1680000637
transform 1 0 576 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_58
timestamp 1680000637
transform 1 0 576 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_59
timestamp 1680000637
transform 1 0 576 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_60
timestamp 1680000637
transform 1 0 576 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_61
timestamp 1680000637
transform 1 0 576 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 576 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 576 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 576 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 576 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 576 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 576 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 576 0 -1 15876
box -48 -56 432 834
use adc  u_adc
timestamp 0
transform 1 0 82800 0 1 1400
box 0 0 1 1
use sg13g2_buf_16  u_clkbuf_analog_pin0.u_buf
timestamp 1676553496
transform 1 0 78144 0 -1 6804
box -48 -56 2448 834
use sg13g2_buf_16  u_clkbuf_analog_pin1.u_buf
timestamp 1676553496
transform 1 0 96288 0 -1 20412
box -48 -56 2448 834
use delay_line  u_delay_line
timestamp 0
transform 1 0 85400 0 1 24600
box 0 0 1 1
use multimode_dll  u_multimode_dll
timestamp 0
transform 1 0 8000 0 1 7400
box 0 0 1 1
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 712 95476 38600 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 99920 33140 100000 33220 0 FreeSans 320 0 0 0 analog_adc
port 2 nsew signal bidirectional
flabel metal3 s 99920 6596 100000 6676 0 FreeSans 320 0 0 0 analog_pin0
port 3 nsew signal bidirectional
flabel metal3 s 99920 19868 100000 19948 0 FreeSans 320 0 0 0 analog_pin1
port 4 nsew signal bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 5 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 6 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 7 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 8 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 9 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 10 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 11 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 12 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 13 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 14 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 15 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 16 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 17 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 18 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 19 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 20 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 21 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 22 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 23 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 24 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 25 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 26 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 27 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 28 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 29 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 30 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 31 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 32 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 33 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 34 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 35 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 36 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 37 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 38 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 39 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 40 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 41 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 42 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 43 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 44 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 45 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 46 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 47 nsew signal output
rlabel via5 65100 24200 65100 24200 0 VGND
rlabel via5 63860 28960 63860 28960 0 VPWR
rlabel metal2 43968 3486 43968 3486 0 _000_
rlabel metal3 20736 37296 20736 37296 0 _001_
rlabel metal2 22704 36876 22704 36876 0 _002_
rlabel metal2 22464 36162 22464 36162 0 _003_
rlabel metal3 26448 35364 26448 35364 0 _004_
rlabel metal2 26304 37464 26304 37464 0 _005_
rlabel metal2 29040 36792 29040 36792 0 _006_
rlabel metal2 29952 37254 29952 37254 0 _007_
rlabel metal2 24672 34440 24672 34440 0 _008_
rlabel metal2 28032 34650 28032 34650 0 _009_
rlabel metal2 29856 35112 29856 35112 0 _010_
rlabel metal2 32448 36414 32448 36414 0 _011_
rlabel metal2 35424 35658 35424 35658 0 _012_
rlabel metal2 47424 34650 47424 34650 0 _013_
rlabel metal2 50592 34902 50592 34902 0 _014_
rlabel metal2 53184 35364 53184 35364 0 _015_
rlabel metal2 54048 34356 54048 34356 0 _016_
rlabel metal2 48000 34902 48000 34902 0 _017_
rlabel metal3 37536 34650 37536 34650 0 _018_
rlabel metal3 35088 35196 35088 35196 0 _019_
rlabel metal2 32160 34440 32160 34440 0 _020_
rlabel metal2 29568 4116 29568 4116 0 _021_
rlabel metal2 31104 4200 31104 4200 0 _022_
rlabel metal2 46320 3528 46320 3528 0 _023_
rlabel metal2 48000 4200 48000 4200 0 _024_
rlabel metal2 50544 3276 50544 3276 0 _025_
rlabel metal2 52368 3528 52368 3528 0 _026_
rlabel metal2 54240 4200 54240 4200 0 _027_
rlabel metal2 50016 2688 50016 2688 0 _028_
rlabel metal2 52080 1932 52080 1932 0 _029_
rlabel metal2 42528 1638 42528 1638 0 _030_
rlabel metal2 45120 1638 45120 1638 0 _031_
rlabel metal2 34368 1638 34368 1638 0 _032_
rlabel metal2 31776 1638 31776 1638 0 _033_
rlabel metal2 29184 2184 29184 2184 0 _034_
rlabel metal2 28224 1092 28224 1092 0 _035_
rlabel metal2 27264 4200 27264 4200 0 _036_
rlabel metal2 26208 4116 26208 4116 0 _037_
rlabel metal2 23424 4410 23424 4410 0 _038_
rlabel metal3 20496 3276 20496 3276 0 _039_
rlabel metal2 21600 4116 21600 4116 0 _040_
rlabel metal2 22464 1974 22464 1974 0 _041_
rlabel metal2 23616 1848 23616 1848 0 _042_
rlabel metal2 26208 1638 26208 1638 0 _043_
rlabel metal3 40320 2016 40320 2016 0 _044_
rlabel metal3 39024 1092 39024 1092 0 _045_
rlabel metal2 36960 1638 36960 1638 0 _046_
rlabel metal2 3456 19026 3456 19026 0 _047_
rlabel metal2 2976 20832 2976 20832 0 _048_
rlabel metal3 3936 23100 3936 23100 0 _049_
rlabel metal2 5088 25011 5088 25011 0 _050_
rlabel metal2 11808 34440 11808 34440 0 _051_
rlabel metal2 14304 35112 14304 35112 0 _052_
rlabel metal2 15072 35868 15072 35868 0 _053_
rlabel metal3 4320 27636 4320 27636 0 _054_
rlabel metal2 4704 9492 4704 9492 0 _055_
rlabel metal2 2496 11088 2496 11088 0 _056_
rlabel metal2 2208 12789 2208 12789 0 _057_
rlabel metal3 1920 13860 1920 13860 0 _058_
rlabel metal3 1920 15372 1920 15372 0 _059_
rlabel metal2 1728 17808 1728 17808 0 _060_
rlabel metal3 1776 20076 1776 20076 0 _061_
rlabel metal3 4080 19908 4080 19908 0 _062_
rlabel metal3 4320 30492 4320 30492 0 _063_
rlabel metal2 16512 34440 16512 34440 0 _064_
rlabel metal2 21024 34860 21024 34860 0 _065_
rlabel metal2 19200 35112 19200 35112 0 _066_
rlabel metal2 16032 4662 16032 4662 0 _067_
rlabel metal2 17664 3654 17664 3654 0 _068_
rlabel metal2 5088 7686 5088 7686 0 _069_
rlabel metal3 4032 12516 4032 12516 0 _070_
rlabel metal2 3456 13230 3456 13230 0 _071_
rlabel metal3 4224 15540 4224 15540 0 _072_
rlabel metal3 4224 17052 4224 17052 0 _073_
rlabel metal2 78240 16968 78240 16968 0 _074_
rlabel metal2 82752 21294 82752 21294 0 _075_
rlabel metal3 81408 25284 81408 25284 0 _076_
rlabel metal2 80592 24696 80592 24696 0 _077_
rlabel metal3 80688 25956 80688 25956 0 _078_
rlabel metal2 80784 28980 80784 28980 0 _079_
rlabel metal2 80064 29904 80064 29904 0 _080_
rlabel metal2 80256 28392 80256 28392 0 _081_
rlabel metal3 81264 27720 81264 27720 0 _082_
rlabel metal2 80832 31878 80832 31878 0 _083_
rlabel metal3 81120 32844 81120 32844 0 _084_
rlabel metal3 80640 33516 80640 33516 0 _085_
rlabel metal2 44352 35868 44352 35868 0 _086_
rlabel metal2 41952 37494 41952 37494 0 _087_
rlabel metal3 41424 36792 41424 36792 0 _088_
rlabel metal3 38496 37296 38496 37296 0 _089_
rlabel metal2 38496 36414 38496 36414 0 _090_
rlabel metal2 41184 34650 41184 34650 0 _091_
rlabel metal2 43728 35364 43728 35364 0 _092_
rlabel metal2 48672 1848 48672 1848 0 _093_
rlabel metal3 18384 36708 18384 36708 0 _094_
rlabel metal3 23472 36708 23472 36708 0 _095_
rlabel metal3 42960 34188 42960 34188 0 _096_
rlabel metal3 44736 3444 44736 3444 0 _097_
rlabel metal2 43872 4200 43872 4200 0 _098_
rlabel metal2 43008 3696 43008 3696 0 _099_
rlabel metal2 38592 5040 38592 5040 0 _100_
rlabel metal2 41280 4830 41280 4830 0 _101_
rlabel metal2 40128 3822 40128 3822 0 _102_
rlabel metal2 41280 3864 41280 3864 0 _103_
rlabel metal3 38640 3360 38640 3360 0 _104_
rlabel metal2 38496 3486 38496 3486 0 _105_
rlabel metal2 35808 1512 35808 1512 0 _106_
rlabel metal2 34848 2742 34848 2742 0 _107_
rlabel metal2 36480 4410 36480 4410 0 _108_
rlabel metal2 36288 3906 36288 3906 0 _109_
rlabel metal2 39360 4872 39360 4872 0 _110_
rlabel metal2 39168 4872 39168 4872 0 _111_
rlabel metal3 21792 37254 21792 37254 0 _112_
rlabel metal2 20640 35868 20640 35868 0 _113_
rlabel via2 26688 36876 26688 36876 0 _114_
rlabel metal3 27120 38220 27120 38220 0 _115_
rlabel metal2 21792 37031 21792 37031 0 _116_
rlabel metal2 19392 36076 19392 36076 0 _117_
rlabel metal3 21648 38388 21648 38388 0 _118_
rlabel metal2 21216 36540 21216 36540 0 _119_
rlabel metal3 23760 36540 23760 36540 0 _120_
rlabel metal2 26208 36540 26208 36540 0 _121_
rlabel metal2 26784 36750 26784 36750 0 _122_
rlabel metal2 28896 38304 28896 38304 0 _123_
rlabel metal2 26064 36876 26064 36876 0 _124_
rlabel metal2 29376 37674 29376 37674 0 _125_
rlabel metal2 41088 34650 41088 34650 0 _126_
rlabel metal2 42912 34608 42912 34608 0 _127_
rlabel metal4 98880 8376 98880 8376 0 adc_data\[0\]
rlabel metal2 31680 2268 31680 2268 0 adc_data\[1\]
rlabel metal2 32736 1932 32736 1932 0 adc_data\[2\]
rlabel metal2 81984 2520 81984 2520 0 adc_data\[3\]
rlabel metal2 35904 1008 35904 1008 0 adc_data\[4\]
rlabel via4 98760 9235 98760 9235 0 adc_data\[5\]
rlabel metal4 98760 8964 98760 8964 0 adc_data\[6\]
rlabel metal2 43392 2604 43392 2604 0 adc_data\[7\]
rlabel metal4 82944 20526 82944 20526 0 analog_adc
rlabel metal3 80496 6384 80496 6384 0 analog_pin0
rlabel metal3 98402 19908 98402 19908 0 analog_pin1
rlabel metal3 3582 36708 3582 36708 0 clk
rlabel metal2 40800 6762 40800 6762 0 clk0_out
rlabel metal2 82752 12600 82752 12600 0 clk1_out
rlabel metal2 37645 7235 37645 7235 0 clk2_out
rlabel metal3 85056 33369 85056 33369 0 clk_delayed
rlabel metal2 43872 4788 43872 4788 0 clk_regs
rlabel metal2 63360 33222 63360 33222 0 clknet_0_clk
rlabel metal2 19872 34440 19872 34440 0 clknet_0_clk_regs
rlabel via2 26382 7140 26382 7140 0 clknet_1_0__leaf_clk
rlabel metal3 98830 9399 98830 9399 0 clknet_1_1__leaf_clk
rlabel metal2 18720 4452 18720 4452 0 clknet_4_0_0_clk_regs
rlabel metal3 81744 21588 81744 21588 0 clknet_4_10_0_clk_regs
rlabel metal2 66912 34272 66912 34272 0 clknet_4_11_0_clk_regs
rlabel metal2 33408 34440 33408 34440 0 clknet_4_12_0_clk_regs
rlabel metal2 70608 37968 70608 37968 0 clknet_4_13_0_clk_regs
rlabel metal2 46368 2394 46368 2394 0 clknet_4_14_0_clk_regs
rlabel metal3 42480 1932 42480 1932 0 clknet_4_15_0_clk_regs
rlabel metal2 4800 13188 4800 13188 0 clknet_4_1_0_clk_regs
rlabel metal3 17808 4032 17808 4032 0 clknet_4_2_0_clk_regs
rlabel metal2 40032 1470 40032 1470 0 clknet_4_3_0_clk_regs
rlabel metal2 4752 18564 4752 18564 0 clknet_4_4_0_clk_regs
rlabel metal2 4752 21588 4752 21588 0 clknet_4_5_0_clk_regs
rlabel metal2 22272 34440 22272 34440 0 clknet_4_6_0_clk_regs
rlabel metal2 17472 35616 17472 35616 0 clknet_4_7_0_clk_regs
rlabel metal4 59808 4410 59808 4410 0 clknet_4_8_0_clk_regs
rlabel metal2 45312 35238 45312 35238 0 clknet_4_9_0_clk_regs
rlabel metal2 29574 31752 29574 31752 0 data\[0\]
rlabel metal2 39744 34062 39744 34062 0 data\[10\]
rlabel metal2 35232 34230 35232 34230 0 data\[11\]
rlabel metal3 10464 5292 10464 5292 0 data\[12\]
rlabel metal2 30720 4578 30720 4578 0 data\[13\]
rlabel metal3 46176 4074 46176 4074 0 data\[14\]
rlabel metal2 47424 5040 47424 5040 0 data\[15\]
rlabel metal2 47232 5700 47232 5700 0 data\[16\]
rlabel metal2 46944 5322 46944 5322 0 data\[17\]
rlabel metal2 47136 6078 47136 6078 0 data\[18\]
rlabel metal2 47376 6048 47376 6048 0 data\[19\]
rlabel metal2 29833 31752 29833 31752 0 data\[1\]
rlabel metal3 40032 2688 40032 2688 0 data\[20\]
rlabel metal2 42528 1134 42528 1134 0 data\[21\]
rlabel metal3 41568 1092 41568 1092 0 data\[22\]
rlabel metal2 44832 1176 44832 1176 0 data\[23\]
rlabel metal3 33216 1092 33216 1092 0 data\[24\]
rlabel metal2 34176 2142 34176 2142 0 data\[25\]
rlabel metal2 31584 2394 31584 2394 0 data\[26\]
rlabel metal2 26688 3402 26688 3402 0 data\[27\]
rlabel metal3 26400 4116 26400 4116 0 data\[28\]
rlabel metal2 26112 5166 26112 5166 0 data\[29\]
rlabel metal2 32185 31752 32185 31752 0 data\[2\]
rlabel metal2 24480 4452 24480 4452 0 data\[30\]
rlabel metal2 21696 4578 21696 4578 0 data\[31\]
rlabel metal2 21792 5166 21792 5166 0 data\[32\]
rlabel metal3 23904 2688 23904 2688 0 data\[33\]
rlabel metal2 23136 2058 23136 2058 0 data\[34\]
rlabel metal2 26208 1176 26208 1176 0 data\[35\]
rlabel metal2 40416 2688 40416 2688 0 data\[36\]
rlabel metal2 39072 2730 39072 2730 0 data\[37\]
rlabel metal2 4032 19404 4032 19404 0 data\[38\]
rlabel metal2 5952 18480 5952 18480 0 data\[39\]
rlabel metal2 31494 31752 31494 31752 0 data\[3\]
rlabel metal2 5376 19740 5376 19740 0 data\[40\]
rlabel metal2 5904 22848 5904 22848 0 data\[41\]
rlabel metal2 15181 31447 15181 31447 0 data\[42\]
rlabel metal2 18816 32970 18816 32970 0 data\[43\]
rlabel metal2 24006 31752 24006 31752 0 data\[44\]
rlabel metal3 17664 35742 17664 35742 0 data\[45\]
rlabel metal2 4032 11256 4032 11256 0 data\[46\]
rlabel metal3 4032 9492 4032 9492 0 data\[47\]
rlabel metal2 4992 11844 4992 11844 0 data\[48\]
rlabel metal2 3264 12642 3264 12642 0 data\[49\]
rlabel metal3 42432 35700 42432 35700 0 data\[4\]
rlabel metal2 1824 15204 1824 15204 0 data\[50\]
rlabel metal2 4032 16674 4032 16674 0 data\[51\]
rlabel metal2 1248 17808 1248 17808 0 data\[52\]
rlabel metal2 4224 19824 4224 19824 0 data\[53\]
rlabel metal3 5616 21504 5616 21504 0 data\[54\]
rlabel metal3 16134 31360 16134 31360 0 data\[55\]
rlabel metal2 18912 34398 18912 34398 0 data\[56\]
rlabel metal2 23622 31752 23622 31752 0 data\[57\]
rlabel metal2 18720 35322 18720 35322 0 data\[58\]
rlabel metal2 18432 6162 18432 6162 0 data\[59\]
rlabel metal2 47136 34356 47136 34356 0 data\[5\]
rlabel metal2 19920 4284 19920 4284 0 data\[60\]
rlabel metal2 4224 12222 4224 12222 0 data\[61\]
rlabel metal2 4320 11760 4320 11760 0 data\[62\]
rlabel metal2 5856 12852 5856 12852 0 data\[63\]
rlabel metal2 5856 16128 5856 16128 0 data\[64\]
rlabel metal2 5856 16758 5856 16758 0 data\[65\]
rlabel metal3 81312 20748 81312 20748 0 data\[66\]
rlabel metal2 82080 20790 82080 20790 0 data\[67\]
rlabel metal2 83232 25746 83232 25746 0 data\[68\]
rlabel metal2 80400 25200 80400 25200 0 data\[69\]
rlabel metal2 52992 33348 52992 33348 0 data\[6\]
rlabel metal2 82896 27048 82896 27048 0 data\[70\]
rlabel metal2 83376 30828 83376 30828 0 data\[71\]
rlabel metal3 82992 30072 82992 30072 0 data\[72\]
rlabel metal2 81312 28854 81312 28854 0 data\[73\]
rlabel metal2 83232 27762 83232 27762 0 data\[74\]
rlabel metal2 83280 32340 83280 32340 0 data\[75\]
rlabel metal2 83184 32676 83184 32676 0 data\[76\]
rlabel metal2 43968 35700 43968 35700 0 data\[77\]
rlabel metal2 43872 35700 43872 35700 0 data\[78\]
rlabel metal2 41664 37254 41664 37254 0 data\[79\]
rlabel metal2 53568 35616 53568 35616 0 data\[7\]
rlabel metal3 42480 38220 42480 38220 0 data\[80\]
rlabel metal2 38880 37830 38880 37830 0 data\[81\]
rlabel metal3 41376 35868 41376 35868 0 data\[82\]
rlabel metal2 43200 34314 43200 34314 0 data\[83\]
rlabel metal2 45216 3528 45216 3528 0 data\[84\]
rlabel metal2 47328 2184 47328 2184 0 data\[85\]
rlabel metal2 46848 33978 46848 33978 0 data\[8\]
rlabel metal2 46944 34734 46944 34734 0 data\[9\]
rlabel metal2 32928 34881 32928 34881 0 delaynet_0_clk
rlabel metal2 2592 7044 2592 7044 0 ena
rlabel metal3 462 15708 462 15708 0 net
rlabel metal3 3168 37968 3168 37968 0 net1
rlabel metal3 2160 9828 2160 9828 0 net10
rlabel metal3 1728 12432 1728 12432 0 net11
rlabel metal2 624 14784 624 14784 0 net12
rlabel metal4 672 9702 672 9702 0 net13
rlabel metal3 4272 17976 4272 17976 0 net14
rlabel via2 1632 18648 1632 18648 0 net15
rlabel metal2 4416 7098 4416 7098 0 net16
rlabel metal2 3744 22302 3744 22302 0 net17
rlabel metal3 20496 35868 20496 35868 0 net18
rlabel metal2 25728 4410 25728 4410 0 net19
rlabel metal2 816 23268 816 23268 0 net2
rlabel metal2 26400 3318 26400 3318 0 net20
rlabel metal3 39792 37212 39792 37212 0 net21
rlabel metal2 41376 34566 41376 34566 0 net22
rlabel metal3 5664 19320 5664 19320 0 net23
rlabel metal2 42480 2436 42480 2436 0 net24
rlabel metal2 46752 35070 46752 35070 0 net25
rlabel metal2 81312 26040 81312 26040 0 net26
rlabel metal2 80736 30954 80736 30954 0 net27
rlabel metal2 41568 35574 41568 35574 0 net28
rlabel metal2 21696 36498 21696 36498 0 net29
rlabel metal3 1008 24024 1008 24024 0 net3
rlabel metal3 2976 18396 2976 18396 0 net30
rlabel metal2 1920 18564 1920 18564 0 net31
rlabel metal3 2496 18480 2496 18480 0 net32
rlabel metal3 3600 20748 3600 20748 0 net33
rlabel metal2 19584 35028 19584 35028 0 net34
rlabel metal3 26256 3444 26256 3444 0 net35
rlabel metal2 26976 4830 26976 4830 0 net36
rlabel metal3 26016 4704 26016 4704 0 net37
rlabel metal2 29472 36792 29472 36792 0 net38
rlabel metal2 23664 37968 23664 37968 0 net39
rlabel metal2 960 24444 960 24444 0 net4
rlabel metal2 41472 36792 41472 36792 0 net40
rlabel metal3 2592 19320 2592 19320 0 net41
rlabel metal2 46656 3108 46656 3108 0 net42
rlabel metal2 44832 35448 44832 35448 0 net43
rlabel metal3 82032 24612 82032 24612 0 net44
rlabel metal2 81216 31962 81216 31962 0 net45
rlabel metal2 45504 35910 45504 35910 0 net46
rlabel metal3 654 16548 654 16548 0 net47
rlabel metal3 462 17388 462 17388 0 net48
rlabel metal3 462 18228 462 18228 0 net49
rlabel metal3 1104 25116 1104 25116 0 net5
rlabel metal3 462 19068 462 19068 0 net50
rlabel metal3 462 19908 462 19908 0 net51
rlabel metal3 462 20748 462 20748 0 net52
rlabel metal3 462 21588 462 21588 0 net53
rlabel metal3 462 2268 462 2268 0 net54
rlabel metal3 462 3108 462 3108 0 net55
rlabel metal3 462 3948 462 3948 0 net56
rlabel metal3 462 4788 462 4788 0 net57
rlabel metal3 462 5628 462 5628 0 net58
rlabel metal3 462 6468 462 6468 0 net59
rlabel metal3 21504 4662 21504 4662 0 net6
rlabel metal3 462 7308 462 7308 0 net60
rlabel metal3 414 8148 414 8148 0 net61
rlabel metal3 816 10248 816 10248 0 net7
rlabel metal3 912 10920 912 10920 0 net8
rlabel metal2 40992 4200 40992 4200 0 net9
rlabel metal2 31776 5364 31776 5364 0 osc_out
rlabel metal3 366 37548 366 37548 0 rst_n
rlabel metal2 34784 7319 34784 7319 0 stable
rlabel metal3 45264 3528 45264 3528 0 u_custom_cells.u_latch0.D
rlabel metal2 47424 2898 47424 2898 0 u_custom_cells.u_latch0.Q
rlabel metal2 22560 37128 22560 37128 0 u_shift_reg.bit_count\[0\]
rlabel metal3 22368 36750 22368 36750 0 u_shift_reg.bit_count\[1\]
rlabel metal2 22944 36792 22944 36792 0 u_shift_reg.bit_count\[2\]
rlabel metal3 26736 36708 26736 36708 0 u_shift_reg.bit_count\[3\]
rlabel metal2 27744 36624 27744 36624 0 u_shift_reg.bit_count\[4\]
rlabel metal3 30480 38220 30480 38220 0 u_shift_reg.bit_count\[5\]
rlabel metal3 28272 37380 28272 37380 0 u_shift_reg.bit_count\[6\]
rlabel metal2 19248 37380 19248 37380 0 u_shift_reg.locked
rlabel metal3 366 22428 366 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 462 8988 462 8988 0 uio_out[0]
rlabel metal3 462 9828 462 9828 0 uio_out[1]
rlabel metal3 462 10668 462 10668 0 uio_out[2]
rlabel metal3 462 11508 462 11508 0 uio_out[3]
rlabel metal3 654 12348 654 12348 0 uio_out[4]
rlabel metal2 816 12684 816 12684 0 uio_out[5]
rlabel metal3 462 14028 462 14028 0 uio_out[6]
rlabel metal3 462 14868 462 14868 0 uio_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
