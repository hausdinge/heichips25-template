magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771577402
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 99360 38576
rect 576 38512 99360 38536
rect 643 38156 701 38157
rect 643 38116 652 38156
rect 692 38116 701 38156
rect 643 38115 701 38116
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 576 37820 99360 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 99360 37820
rect 576 37756 99360 37780
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 99360 37064
rect 576 37000 99360 37024
rect 576 36308 99360 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 99360 36308
rect 576 36244 99360 36268
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 99360 35552
rect 576 35488 99360 35512
rect 576 34796 99360 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 99360 34796
rect 576 34732 99360 34756
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 99360 34040
rect 576 33976 99360 34000
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 99360 33284
rect 576 33220 99360 33244
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 99360 32528
rect 576 32464 99360 32488
rect 576 31772 99360 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 99360 31772
rect 576 31708 99360 31732
rect 576 31016 99360 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 99360 31016
rect 576 30952 99360 30976
rect 576 30260 99360 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 99360 30260
rect 576 30196 99360 30220
rect 576 29504 99360 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 99360 29504
rect 576 29440 99360 29464
rect 576 28748 99360 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 99360 28748
rect 576 28684 99360 28708
rect 576 27992 99360 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 99360 27992
rect 576 27928 99360 27952
rect 576 27236 99360 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 99360 27236
rect 576 27172 99360 27196
rect 576 26480 99360 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 99360 26480
rect 576 26416 99360 26440
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 99360 25724
rect 576 25660 99360 25684
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 99360 24968
rect 576 24904 99360 24928
rect 576 24212 99360 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 99360 24212
rect 576 24148 99360 24172
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 99360 23456
rect 576 23392 99360 23416
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 843 22868 885 22877
rect 843 22828 844 22868
rect 884 22828 885 22868
rect 843 22819 885 22828
rect 576 22700 99360 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 99360 22700
rect 576 22636 99360 22660
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 576 21880 99360 21904
rect 4971 21692 5013 21701
rect 4971 21652 4972 21692
rect 5012 21652 5013 21692
rect 4971 21643 5013 21652
rect 5347 21608 5405 21609
rect 5347 21568 5356 21608
rect 5396 21568 5405 21608
rect 5347 21567 5405 21568
rect 6211 21608 6269 21609
rect 6211 21568 6220 21608
rect 6260 21568 6269 21608
rect 6211 21567 6269 21568
rect 7363 21356 7421 21357
rect 7363 21316 7372 21356
rect 7412 21316 7421 21356
rect 7363 21315 7421 21316
rect 576 21188 99360 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 576 21124 99360 21148
rect 3243 21020 3285 21029
rect 3243 20980 3244 21020
rect 3284 20980 3285 21020
rect 3243 20971 3285 20980
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 5355 20936 5397 20945
rect 5355 20896 5356 20936
rect 5396 20896 5397 20936
rect 5355 20887 5397 20896
rect 2571 20768 2613 20777
rect 2571 20728 2572 20768
rect 2612 20728 2613 20768
rect 2571 20719 2613 20728
rect 2667 20768 2709 20777
rect 2667 20728 2668 20768
rect 2708 20728 2709 20768
rect 2667 20719 2709 20728
rect 2763 20768 2805 20777
rect 2763 20728 2764 20768
rect 2804 20728 2805 20768
rect 2763 20719 2805 20728
rect 2859 20768 2901 20777
rect 2859 20728 2860 20768
rect 2900 20728 2901 20768
rect 2859 20719 2901 20728
rect 3243 20768 3285 20777
rect 3243 20728 3244 20768
rect 3284 20728 3285 20768
rect 3243 20719 3285 20728
rect 3435 20768 3477 20777
rect 3435 20728 3436 20768
rect 3476 20728 3477 20768
rect 3435 20719 3477 20728
rect 3523 20768 3581 20769
rect 3523 20728 3532 20768
rect 3572 20728 3581 20768
rect 3523 20727 3581 20728
rect 5547 20768 5589 20777
rect 5547 20728 5548 20768
rect 5588 20728 5589 20768
rect 5547 20719 5589 20728
rect 6211 20768 6269 20769
rect 6211 20728 6220 20768
rect 6260 20728 6269 20768
rect 6211 20727 6269 20728
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 576 20368 99360 20392
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 576 19676 99360 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 576 19612 99360 19636
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 99360 18920
rect 576 18856 99360 18880
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 576 18164 99360 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 99360 18164
rect 576 18100 99360 18124
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 7659 17744 7701 17753
rect 7659 17704 7660 17744
rect 7700 17704 7701 17744
rect 7659 17695 7701 17704
rect 8035 17744 8093 17745
rect 8035 17704 8044 17744
rect 8084 17704 8093 17744
rect 8035 17703 8093 17704
rect 8899 17744 8957 17745
rect 8899 17704 8908 17744
rect 8948 17704 8957 17744
rect 8899 17703 8957 17704
rect 10051 17576 10109 17577
rect 10051 17536 10060 17576
rect 10100 17536 10109 17576
rect 10051 17535 10109 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 99360 17408
rect 576 17344 99360 17368
rect 8131 17240 8189 17241
rect 8131 17200 8140 17240
rect 8180 17200 8189 17240
rect 8131 17199 8189 17200
rect 8803 17072 8861 17073
rect 8803 17032 8812 17072
rect 8852 17032 8861 17072
rect 8803 17031 8861 17032
rect 10147 17072 10205 17073
rect 10147 17032 10156 17072
rect 10196 17032 10205 17072
rect 10147 17031 10205 17032
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 7947 16904 7989 16913
rect 7947 16864 7948 16904
rect 7988 16864 7989 16904
rect 7947 16855 7989 16864
rect 9475 16820 9533 16821
rect 9475 16780 9484 16820
rect 9524 16780 9533 16820
rect 9475 16779 9533 16780
rect 576 16652 99360 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 99360 16652
rect 576 16588 99360 16612
rect 8427 16484 8469 16493
rect 8427 16444 8428 16484
rect 8468 16444 8469 16484
rect 8427 16435 8469 16444
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 8427 16232 8469 16241
rect 8427 16192 8428 16232
rect 8468 16192 8469 16232
rect 8427 16183 8469 16192
rect 8619 16232 8661 16241
rect 8619 16192 8620 16232
rect 8660 16192 8661 16232
rect 8619 16183 8661 16192
rect 8707 16232 8765 16233
rect 8707 16192 8716 16232
rect 8756 16192 8765 16232
rect 8707 16191 8765 16192
rect 9003 16232 9045 16241
rect 9003 16192 9004 16232
rect 9044 16192 9045 16232
rect 9003 16183 9045 16192
rect 9099 16232 9141 16241
rect 9099 16192 9100 16232
rect 9140 16192 9141 16232
rect 9099 16183 9141 16192
rect 9195 16232 9237 16241
rect 9195 16192 9196 16232
rect 9236 16192 9237 16232
rect 9195 16183 9237 16192
rect 8899 16064 8957 16065
rect 8899 16024 8908 16064
rect 8948 16024 8957 16064
rect 8899 16023 8957 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 99360 15896
rect 576 15832 99360 15856
rect 9003 15728 9045 15737
rect 9003 15688 9004 15728
rect 9044 15688 9045 15728
rect 9003 15679 9045 15688
rect 10915 15560 10973 15561
rect 10915 15520 10924 15560
rect 10964 15520 10973 15560
rect 10915 15519 10973 15520
rect 835 15476 893 15477
rect 835 15436 844 15476
rect 884 15436 893 15476
rect 835 15435 893 15436
rect 9571 15476 9629 15477
rect 9571 15436 9580 15476
rect 9620 15436 9629 15476
rect 9571 15435 9629 15436
rect 13611 15392 13653 15401
rect 13611 15352 13612 15392
rect 13652 15352 13653 15392
rect 13611 15343 13653 15352
rect 651 15308 693 15317
rect 651 15268 652 15308
rect 692 15268 693 15308
rect 651 15259 693 15268
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 99360 15140
rect 576 15076 99360 15100
rect 835 14804 893 14805
rect 835 14764 844 14804
rect 884 14764 893 14804
rect 835 14763 893 14764
rect 13507 14720 13565 14721
rect 13507 14680 13516 14720
rect 13556 14680 13565 14720
rect 13507 14679 13565 14680
rect 14371 14720 14429 14721
rect 14371 14680 14380 14720
rect 14420 14680 14429 14720
rect 14371 14679 14429 14680
rect 13131 14636 13173 14645
rect 13131 14596 13132 14636
rect 13172 14596 13173 14636
rect 13131 14587 13173 14596
rect 651 14552 693 14561
rect 651 14512 652 14552
rect 692 14512 693 14552
rect 651 14503 693 14512
rect 15523 14552 15581 14553
rect 15523 14512 15532 14552
rect 15572 14512 15581 14552
rect 15523 14511 15581 14512
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 99360 14384
rect 576 14320 99360 14344
rect 11299 14216 11357 14217
rect 11299 14176 11308 14216
rect 11348 14176 11357 14216
rect 11299 14175 11357 14176
rect 3907 14048 3965 14049
rect 3907 14008 3916 14048
rect 3956 14008 3965 14048
rect 3907 14007 3965 14008
rect 4771 14048 4829 14049
rect 4771 14008 4780 14048
rect 4820 14008 4829 14048
rect 4771 14007 4829 14008
rect 5163 14048 5205 14057
rect 5163 14008 5164 14048
rect 5204 14008 5205 14048
rect 5163 13999 5205 14008
rect 11107 14048 11165 14049
rect 11107 14008 11116 14048
rect 11156 14008 11165 14048
rect 11107 14007 11165 14008
rect 11211 14048 11253 14057
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 11403 14048 11445 14057
rect 11403 14008 11404 14048
rect 11444 14008 11445 14048
rect 11403 13999 11445 14008
rect 13515 14048 13557 14057
rect 13515 14008 13516 14048
rect 13556 14008 13557 14048
rect 13515 13999 13557 14008
rect 14179 14048 14237 14049
rect 14179 14008 14188 14048
rect 14228 14008 14237 14048
rect 14179 14007 14237 14008
rect 2755 13796 2813 13797
rect 2755 13756 2764 13796
rect 2804 13756 2813 13796
rect 2755 13755 2813 13756
rect 576 13628 99360 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 99360 13628
rect 576 13564 99360 13588
rect 4011 13376 4053 13385
rect 4011 13336 4012 13376
rect 4052 13336 4053 13376
rect 4011 13327 4053 13336
rect 835 13292 893 13293
rect 835 13252 844 13292
rect 884 13252 893 13292
rect 835 13251 893 13252
rect 3619 13208 3677 13209
rect 3619 13168 3628 13208
rect 3668 13168 3677 13208
rect 3619 13167 3677 13168
rect 10155 13208 10197 13217
rect 10155 13168 10156 13208
rect 10196 13168 10197 13208
rect 10155 13159 10197 13168
rect 10251 13208 10293 13217
rect 10251 13168 10252 13208
rect 10292 13168 10293 13208
rect 10251 13159 10293 13168
rect 10347 13208 10389 13217
rect 10347 13168 10348 13208
rect 10388 13168 10389 13208
rect 10347 13159 10389 13168
rect 10443 13208 10485 13217
rect 10443 13168 10444 13208
rect 10484 13168 10485 13208
rect 10443 13159 10485 13168
rect 651 13040 693 13049
rect 651 13000 652 13040
rect 692 13000 693 13040
rect 651 12991 693 13000
rect 2947 13040 3005 13041
rect 2947 13000 2956 13040
rect 2996 13000 3005 13040
rect 2947 12999 3005 13000
rect 576 12872 99360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 99360 12872
rect 576 12808 99360 12832
rect 9859 12536 9917 12537
rect 9859 12496 9868 12536
rect 9908 12496 9917 12536
rect 9859 12495 9917 12496
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 11299 12452 11357 12453
rect 11299 12412 11308 12452
rect 11348 12412 11357 12452
rect 11299 12411 11357 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 576 12116 99360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 99360 12116
rect 576 12052 99360 12076
rect 2571 11864 2613 11873
rect 2571 11824 2572 11864
rect 2612 11824 2613 11864
rect 2571 11815 2613 11824
rect 4491 11864 4533 11873
rect 4491 11824 4492 11864
rect 4532 11824 4533 11864
rect 4491 11815 4533 11824
rect 8515 11864 8573 11865
rect 8515 11824 8524 11864
rect 8564 11824 8573 11864
rect 8515 11823 8573 11824
rect 9963 11864 10005 11873
rect 9963 11824 9964 11864
rect 10004 11824 10005 11864
rect 9963 11815 10005 11824
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 2275 11696 2333 11697
rect 2275 11656 2284 11696
rect 2324 11656 2333 11696
rect 2275 11655 2333 11656
rect 2379 11696 2421 11705
rect 2379 11656 2380 11696
rect 2420 11656 2421 11696
rect 2379 11647 2421 11656
rect 2571 11696 2613 11705
rect 2571 11656 2572 11696
rect 2612 11656 2613 11696
rect 2571 11647 2613 11656
rect 2955 11696 2997 11705
rect 2955 11656 2956 11696
rect 2996 11656 2997 11696
rect 2955 11647 2997 11656
rect 3051 11696 3093 11705
rect 3051 11656 3052 11696
rect 3092 11656 3093 11696
rect 3051 11647 3093 11656
rect 3427 11696 3485 11697
rect 3427 11656 3436 11696
rect 3476 11656 3485 11696
rect 3427 11655 3485 11656
rect 4107 11696 4149 11705
rect 4107 11656 4108 11696
rect 4148 11656 4149 11696
rect 4107 11647 4149 11656
rect 4299 11696 4341 11705
rect 4299 11656 4300 11696
rect 4340 11656 4341 11696
rect 4299 11647 4341 11656
rect 4395 11696 4437 11705
rect 4395 11656 4396 11696
rect 4436 11656 4437 11696
rect 4395 11647 4437 11656
rect 4587 11696 4629 11705
rect 4587 11656 4588 11696
rect 4628 11656 4629 11696
rect 4587 11647 4629 11656
rect 8715 11696 8757 11705
rect 8715 11656 8716 11696
rect 8756 11656 8757 11696
rect 8715 11647 8757 11656
rect 8811 11696 8853 11705
rect 8811 11656 8812 11696
rect 8852 11656 8853 11696
rect 8811 11647 8853 11656
rect 8907 11696 8949 11705
rect 8907 11656 8908 11696
rect 8948 11656 8949 11696
rect 8907 11647 8949 11656
rect 9003 11696 9045 11705
rect 9003 11656 9004 11696
rect 9044 11656 9045 11696
rect 9003 11647 9045 11656
rect 9667 11696 9725 11697
rect 9667 11656 9676 11696
rect 9716 11656 9725 11696
rect 9667 11655 9725 11656
rect 9771 11696 9813 11705
rect 9771 11656 9772 11696
rect 9812 11656 9813 11696
rect 9771 11647 9813 11656
rect 9963 11696 10005 11705
rect 9963 11656 9964 11696
rect 10004 11656 10005 11696
rect 9963 11647 10005 11656
rect 10819 11696 10877 11697
rect 10819 11656 10828 11696
rect 10868 11656 10877 11696
rect 10819 11655 10877 11656
rect 12067 11696 12125 11697
rect 12067 11656 12076 11696
rect 12116 11656 12125 11696
rect 12067 11655 12125 11656
rect 13419 11696 13461 11705
rect 13419 11656 13420 11696
rect 13460 11656 13461 11696
rect 13419 11647 13461 11656
rect 14083 11696 14141 11697
rect 14083 11656 14092 11696
rect 14132 11656 14141 11696
rect 14083 11655 14141 11656
rect 3235 11612 3293 11613
rect 3235 11572 3244 11612
rect 3284 11572 3293 11612
rect 3235 11571 3293 11572
rect 10155 11612 10197 11621
rect 10155 11572 10156 11612
rect 10196 11572 10197 11612
rect 10155 11563 10197 11572
rect 12747 11612 12789 11621
rect 12747 11572 12748 11612
rect 12788 11572 12789 11612
rect 12747 11563 12789 11572
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 2947 11528 3005 11529
rect 2947 11488 2956 11528
rect 2996 11488 3005 11528
rect 2947 11487 3005 11488
rect 576 11360 99360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 99360 11360
rect 576 11296 99360 11320
rect 9187 11192 9245 11193
rect 9187 11152 9196 11192
rect 9236 11152 9245 11192
rect 9187 11151 9245 11152
rect 9475 11192 9533 11193
rect 9475 11152 9484 11192
rect 9524 11152 9533 11192
rect 9475 11151 9533 11152
rect 9771 11192 9813 11201
rect 9771 11152 9772 11192
rect 9812 11152 9813 11192
rect 9771 11143 9813 11152
rect 16483 11192 16541 11193
rect 16483 11152 16492 11192
rect 16532 11152 16541 11192
rect 16483 11151 16541 11152
rect 14091 11108 14133 11117
rect 14091 11068 14092 11108
rect 14132 11068 14133 11108
rect 14091 11059 14133 11068
rect 9283 11024 9341 11025
rect 9283 10984 9292 11024
rect 9332 10984 9341 11024
rect 9283 10983 9341 10984
rect 9675 11024 9717 11033
rect 9675 10984 9676 11024
rect 9716 10984 9717 11024
rect 9675 10975 9717 10984
rect 9867 11024 9909 11033
rect 9867 10984 9868 11024
rect 9908 10984 9909 11024
rect 9867 10975 9909 10984
rect 9963 11024 10005 11033
rect 9963 10984 9964 11024
rect 10004 10984 10005 11024
rect 9963 10975 10005 10984
rect 14467 11024 14525 11025
rect 14467 10984 14476 11024
rect 14516 10984 14525 11024
rect 14467 10983 14525 10984
rect 15331 11024 15389 11025
rect 15331 10984 15340 11024
rect 15380 10984 15389 11024
rect 15331 10983 15389 10984
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 576 10604 99360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 99360 10604
rect 576 10540 99360 10564
rect 14571 10352 14613 10361
rect 14571 10312 14572 10352
rect 14612 10312 14613 10352
rect 14571 10303 14613 10312
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 576 9848 99360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 99360 9848
rect 576 9784 99360 9808
rect 4203 9680 4245 9689
rect 4203 9640 4204 9680
rect 4244 9640 4245 9680
rect 4203 9631 4245 9640
rect 12459 9680 12501 9689
rect 12459 9640 12460 9680
rect 12500 9640 12501 9680
rect 12459 9631 12501 9640
rect 4099 9512 4157 9513
rect 4099 9472 4108 9512
rect 4148 9472 4157 9512
rect 4099 9471 4157 9472
rect 10531 9512 10589 9513
rect 10531 9472 10540 9512
rect 10580 9472 10589 9512
rect 10531 9471 10589 9472
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 2851 9428 2909 9429
rect 2851 9388 2860 9428
rect 2900 9388 2909 9428
rect 2851 9387 2909 9388
rect 651 9260 693 9269
rect 651 9220 652 9260
rect 692 9220 693 9260
rect 651 9211 693 9220
rect 2667 9260 2709 9269
rect 2667 9220 2668 9260
rect 2708 9220 2709 9260
rect 2667 9211 2709 9220
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 2283 8840 2325 8849
rect 2283 8800 2284 8840
rect 2324 8800 2325 8840
rect 2283 8791 2325 8800
rect 7371 8840 7413 8849
rect 7371 8800 7372 8840
rect 7412 8800 7413 8840
rect 7371 8791 7413 8800
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 2467 8756 2525 8757
rect 2467 8716 2476 8756
rect 2516 8716 2525 8756
rect 2467 8715 2525 8716
rect 2851 8756 2909 8757
rect 2851 8716 2860 8756
rect 2900 8716 2909 8756
rect 2851 8715 2909 8716
rect 7179 8697 7221 8706
rect 7083 8672 7125 8681
rect 7083 8632 7084 8672
rect 7124 8632 7125 8672
rect 7179 8657 7180 8697
rect 7220 8657 7221 8697
rect 7179 8648 7221 8657
rect 7083 8623 7125 8632
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 2667 8504 2709 8513
rect 2667 8464 2668 8504
rect 2708 8464 2709 8504
rect 2667 8455 2709 8464
rect 7075 8504 7133 8505
rect 7075 8464 7084 8504
rect 7124 8464 7133 8504
rect 7075 8463 7133 8464
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 9187 8168 9245 8169
rect 9187 8128 9196 8168
rect 9236 8128 9245 8168
rect 9187 8127 9245 8128
rect 8419 8000 8477 8001
rect 8419 7960 8428 8000
rect 8468 7960 8477 8000
rect 8419 7959 8477 7960
rect 8523 8000 8565 8009
rect 8523 7960 8524 8000
rect 8564 7960 8565 8000
rect 8523 7951 8565 7960
rect 8707 8000 8765 8001
rect 8707 7960 8716 8000
rect 8756 7960 8765 8000
rect 8707 7959 8765 7960
rect 8803 8000 8861 8001
rect 8803 7960 8812 8000
rect 8852 7960 8861 8000
rect 8803 7959 8861 7960
rect 9003 8000 9045 8009
rect 9003 7960 9004 8000
rect 9044 7960 9045 8000
rect 9003 7951 9045 7960
rect 9099 8000 9141 8009
rect 9099 7960 9100 8000
rect 9140 7960 9141 8000
rect 9099 7951 9141 7960
rect 9246 8000 9304 8001
rect 9246 7960 9255 8000
rect 9295 7960 9304 8000
rect 9246 7959 9304 7960
rect 10435 8000 10493 8001
rect 10435 7960 10444 8000
rect 10484 7960 10493 8000
rect 10435 7959 10493 7960
rect 12067 8000 12125 8001
rect 12067 7960 12076 8000
rect 12116 7960 12125 8000
rect 12067 7959 12125 7960
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 2851 7916 2909 7917
rect 2851 7876 2860 7916
rect 2900 7876 2909 7916
rect 2851 7875 2909 7876
rect 11403 7916 11445 7925
rect 11403 7876 11404 7916
rect 11444 7876 11445 7916
rect 11403 7867 11445 7876
rect 12267 7832 12309 7841
rect 12267 7792 12268 7832
rect 12308 7792 12309 7832
rect 12267 7783 12309 7792
rect 651 7748 693 7757
rect 651 7708 652 7748
rect 692 7708 693 7748
rect 651 7699 693 7708
rect 2667 7748 2709 7757
rect 2667 7708 2668 7748
rect 2708 7708 2709 7748
rect 2667 7699 2709 7708
rect 11107 7748 11165 7749
rect 11107 7708 11116 7748
rect 11156 7708 11165 7748
rect 11107 7707 11165 7708
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 5547 7412 5589 7421
rect 5547 7372 5548 7412
rect 5588 7372 5589 7412
rect 5547 7363 5589 7372
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 5251 7160 5309 7161
rect 5251 7120 5260 7160
rect 5300 7120 5309 7160
rect 5251 7119 5309 7120
rect 5355 7160 5397 7169
rect 5355 7120 5356 7160
rect 5396 7120 5397 7160
rect 5355 7111 5397 7120
rect 5539 7160 5597 7161
rect 5539 7120 5548 7160
rect 5588 7120 5597 7160
rect 5539 7119 5597 7120
rect 11691 7160 11733 7169
rect 11691 7120 11692 7160
rect 11732 7120 11733 7160
rect 11691 7111 11733 7120
rect 12067 7160 12125 7161
rect 12067 7120 12076 7160
rect 12116 7120 12125 7160
rect 12067 7119 12125 7120
rect 12931 7160 12989 7161
rect 12931 7120 12940 7160
rect 12980 7120 12989 7160
rect 12931 7119 12989 7120
rect 651 6992 693 7001
rect 651 6952 652 6992
rect 692 6952 693 6992
rect 651 6943 693 6952
rect 14083 6992 14141 6993
rect 14083 6952 14092 6992
rect 14132 6952 14141 6992
rect 14083 6951 14141 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 4771 6488 4829 6489
rect 4771 6448 4780 6488
rect 4820 6448 4829 6488
rect 4771 6447 4829 6448
rect 4971 6488 5013 6497
rect 4971 6448 4972 6488
rect 5012 6448 5013 6488
rect 4971 6439 5013 6448
rect 2851 6404 2909 6405
rect 2851 6364 2860 6404
rect 2900 6364 2909 6404
rect 2851 6363 2909 6364
rect 2667 6236 2709 6245
rect 2667 6196 2668 6236
rect 2708 6196 2709 6236
rect 2667 6187 2709 6196
rect 4875 6236 4917 6245
rect 4875 6196 4876 6236
rect 4916 6196 4917 6236
rect 4875 6187 4917 6196
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 835 5732 893 5733
rect 835 5692 844 5732
rect 884 5692 893 5732
rect 835 5691 893 5692
rect 4963 5648 5021 5649
rect 4963 5608 4972 5648
rect 5012 5608 5021 5648
rect 4963 5607 5021 5608
rect 651 5480 693 5489
rect 651 5440 652 5480
rect 692 5440 693 5480
rect 651 5431 693 5440
rect 4291 5480 4349 5481
rect 4291 5440 4300 5480
rect 4340 5440 4349 5480
rect 4291 5439 4349 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 4003 5144 4061 5145
rect 4003 5104 4012 5144
rect 4052 5104 4061 5144
rect 4003 5103 4061 5104
rect 3811 4976 3869 4977
rect 3811 4936 3820 4976
rect 3860 4936 3869 4976
rect 3811 4935 3869 4936
rect 3915 4976 3957 4985
rect 3915 4936 3916 4976
rect 3956 4936 3957 4976
rect 3915 4927 3957 4936
rect 4107 4976 4149 4985
rect 4107 4936 4108 4976
rect 4148 4936 4149 4976
rect 4107 4927 4149 4936
rect 4299 4976 4341 4985
rect 4299 4936 4300 4976
rect 4340 4936 4341 4976
rect 4299 4927 4341 4936
rect 4491 4976 4533 4985
rect 4491 4936 4492 4976
rect 4532 4936 4533 4976
rect 4491 4927 4533 4936
rect 9195 4976 9237 4985
rect 9195 4936 9196 4976
rect 9236 4936 9237 4976
rect 9195 4927 9237 4936
rect 9291 4976 9333 4985
rect 9291 4936 9292 4976
rect 9332 4936 9333 4976
rect 9291 4927 9333 4936
rect 9387 4976 9429 4985
rect 9387 4936 9388 4976
rect 9428 4936 9429 4976
rect 9387 4927 9429 4936
rect 9483 4976 9525 4985
rect 9483 4936 9484 4976
rect 9524 4936 9525 4976
rect 9483 4927 9525 4936
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 2851 4892 2909 4893
rect 2851 4852 2860 4892
rect 2900 4852 2909 4892
rect 2851 4851 2909 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 2667 4808 2709 4817
rect 2667 4768 2668 4808
rect 2708 4768 2709 4808
rect 2667 4759 2709 4768
rect 4491 4724 4533 4733
rect 4491 4684 4492 4724
rect 4532 4684 4533 4724
rect 4491 4675 4533 4684
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 2667 4304 2709 4313
rect 2667 4264 2668 4304
rect 2708 4264 2709 4304
rect 2667 4255 2709 4264
rect 5155 4304 5213 4305
rect 5155 4264 5164 4304
rect 5204 4264 5213 4304
rect 5155 4263 5213 4264
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 2851 4220 2909 4221
rect 2851 4180 2860 4220
rect 2900 4180 2909 4220
rect 2851 4179 2909 4180
rect 4771 4136 4829 4137
rect 4771 4096 4780 4136
rect 4820 4096 4829 4136
rect 4771 4095 4829 4096
rect 5827 4136 5885 4137
rect 5827 4096 5836 4136
rect 5876 4096 5885 4136
rect 5827 4095 5885 4096
rect 9291 4136 9333 4145
rect 9291 4096 9292 4136
rect 9332 4096 9333 4136
rect 9291 4087 9333 4096
rect 9483 4136 9525 4145
rect 9483 4096 9484 4136
rect 9524 4096 9525 4136
rect 9483 4087 9525 4096
rect 9571 4136 9629 4137
rect 9571 4096 9580 4136
rect 9620 4096 9629 4136
rect 9571 4095 9629 4096
rect 10635 4136 10677 4145
rect 10635 4096 10636 4136
rect 10676 4096 10677 4136
rect 10635 4087 10677 4096
rect 11299 4136 11357 4137
rect 11299 4096 11308 4136
rect 11348 4096 11357 4136
rect 11299 4095 11357 4096
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 4099 3968 4157 3969
rect 4099 3928 4108 3968
rect 4148 3928 4157 3968
rect 4099 3927 4157 3928
rect 9379 3968 9437 3969
rect 9379 3928 9388 3968
rect 9428 3928 9437 3968
rect 9379 3927 9437 3928
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 11587 3632 11645 3633
rect 11587 3592 11596 3632
rect 11636 3592 11645 3632
rect 11587 3591 11645 3592
rect 9195 3548 9237 3557
rect 9195 3508 9196 3548
rect 9236 3508 9237 3548
rect 9195 3499 9237 3508
rect 9571 3464 9629 3465
rect 9571 3424 9580 3464
rect 9620 3424 9629 3464
rect 9571 3423 9629 3424
rect 10435 3464 10493 3465
rect 10435 3424 10444 3464
rect 10484 3424 10493 3464
rect 10435 3423 10493 3424
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 4107 3296 4149 3305
rect 4107 3256 4108 3296
rect 4148 3256 4149 3296
rect 4107 3247 4149 3256
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 6019 2876 6077 2877
rect 6019 2836 6028 2876
rect 6068 2836 6077 2876
rect 6019 2835 6077 2836
rect 2667 2792 2709 2801
rect 2667 2752 2668 2792
rect 2708 2752 2709 2792
rect 2667 2743 2709 2752
rect 9675 2792 9717 2801
rect 9675 2752 9676 2792
rect 9716 2752 9717 2792
rect 9675 2743 9717 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 2851 2708 2909 2709
rect 2851 2668 2860 2708
rect 2900 2668 2909 2708
rect 2851 2667 2909 2668
rect 3627 2624 3669 2633
rect 3627 2584 3628 2624
rect 3668 2584 3669 2624
rect 3627 2575 3669 2584
rect 4003 2624 4061 2625
rect 4003 2584 4012 2624
rect 4052 2584 4061 2624
rect 4003 2583 4061 2584
rect 4867 2624 4925 2625
rect 4867 2584 4876 2624
rect 4916 2584 4925 2624
rect 4867 2583 4925 2584
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 652 38116 692 38156
rect 844 37948 884 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 652 22996 692 23036
rect 844 22828 884 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 652 22408 692 22448
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 4972 21652 5012 21692
rect 5356 21568 5396 21608
rect 6220 21568 6260 21608
rect 7372 21316 7412 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 3244 20980 3284 21020
rect 652 20896 692 20936
rect 5356 20896 5396 20936
rect 2572 20728 2612 20768
rect 2668 20728 2708 20768
rect 2764 20728 2804 20768
rect 2860 20728 2900 20768
rect 3244 20728 3284 20768
rect 3436 20728 3476 20768
rect 3532 20728 3572 20768
rect 5548 20728 5588 20768
rect 6220 20728 6260 20768
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 652 19888 692 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 652 19384 692 19424
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 652 18376 692 18416
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 652 17872 692 17912
rect 7660 17704 7700 17744
rect 8044 17704 8084 17744
rect 8908 17704 8948 17744
rect 10060 17536 10100 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 8140 17200 8180 17240
rect 8812 17032 8852 17072
rect 10156 17032 10196 17072
rect 652 16864 692 16904
rect 7948 16864 7988 16904
rect 9484 16780 9524 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 8428 16444 8468 16484
rect 652 16360 692 16400
rect 8428 16192 8468 16232
rect 8620 16192 8660 16232
rect 8716 16192 8756 16232
rect 9004 16192 9044 16232
rect 9100 16192 9140 16232
rect 9196 16192 9236 16232
rect 8908 16024 8948 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 9004 15688 9044 15728
rect 10924 15520 10964 15560
rect 844 15436 884 15476
rect 9580 15436 9620 15476
rect 13612 15352 13652 15392
rect 652 15268 692 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 844 14764 884 14804
rect 13516 14680 13556 14720
rect 14380 14680 14420 14720
rect 13132 14596 13172 14636
rect 652 14512 692 14552
rect 15532 14512 15572 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 11308 14176 11348 14216
rect 3916 14008 3956 14048
rect 4780 14008 4820 14048
rect 5164 14008 5204 14048
rect 11116 14008 11156 14048
rect 11212 14008 11252 14048
rect 11404 14008 11444 14048
rect 13516 14008 13556 14048
rect 14188 14008 14228 14048
rect 2764 13756 2804 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4012 13336 4052 13376
rect 844 13252 884 13292
rect 3628 13168 3668 13208
rect 10156 13168 10196 13208
rect 10252 13168 10292 13208
rect 10348 13168 10388 13208
rect 10444 13168 10484 13208
rect 652 13000 692 13040
rect 2956 13000 2996 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 9868 12496 9908 12536
rect 844 12412 884 12452
rect 11308 12412 11348 12452
rect 652 12328 692 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 2572 11824 2612 11864
rect 4492 11824 4532 11864
rect 8524 11824 8564 11864
rect 9964 11824 10004 11864
rect 844 11740 884 11780
rect 2284 11656 2324 11696
rect 2380 11656 2420 11696
rect 2572 11656 2612 11696
rect 2956 11656 2996 11696
rect 3052 11656 3092 11696
rect 3436 11656 3476 11696
rect 4108 11656 4148 11696
rect 4300 11656 4340 11696
rect 4396 11656 4436 11696
rect 4588 11656 4628 11696
rect 8716 11656 8756 11696
rect 8812 11656 8852 11696
rect 8908 11656 8948 11696
rect 9004 11656 9044 11696
rect 9676 11656 9716 11696
rect 9772 11656 9812 11696
rect 9964 11656 10004 11696
rect 10828 11656 10868 11696
rect 12076 11656 12116 11696
rect 13420 11656 13460 11696
rect 14092 11656 14132 11696
rect 3244 11572 3284 11612
rect 10156 11572 10196 11612
rect 12748 11572 12788 11612
rect 652 11488 692 11528
rect 2956 11488 2996 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 9196 11152 9236 11192
rect 9484 11152 9524 11192
rect 9772 11152 9812 11192
rect 16492 11152 16532 11192
rect 14092 11068 14132 11108
rect 9292 10984 9332 11024
rect 9676 10984 9716 11024
rect 9868 10984 9908 11024
rect 9964 10984 10004 11024
rect 14476 10984 14516 11024
rect 15340 10984 15380 11024
rect 844 10900 884 10940
rect 652 10732 692 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 14572 10312 14612 10352
rect 844 10228 884 10268
rect 652 9976 692 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 4204 9640 4244 9680
rect 12460 9640 12500 9680
rect 4108 9472 4148 9512
rect 10540 9472 10580 9512
rect 844 9388 884 9428
rect 2860 9388 2900 9428
rect 652 9220 692 9260
rect 2668 9220 2708 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 2284 8800 2324 8840
rect 7372 8800 7412 8840
rect 844 8716 884 8756
rect 2476 8716 2516 8756
rect 2860 8716 2900 8756
rect 7084 8632 7124 8672
rect 7180 8657 7220 8697
rect 652 8464 692 8504
rect 2668 8464 2708 8504
rect 7084 8464 7124 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 9196 8128 9236 8168
rect 8428 7960 8468 8000
rect 8524 7960 8564 8000
rect 8716 7960 8756 8000
rect 8812 7960 8852 8000
rect 9004 7960 9044 8000
rect 9100 7960 9140 8000
rect 9255 7960 9295 8000
rect 10444 7960 10484 8000
rect 12076 7960 12116 8000
rect 844 7876 884 7916
rect 2860 7876 2900 7916
rect 11404 7876 11444 7916
rect 12268 7792 12308 7832
rect 652 7708 692 7748
rect 2668 7708 2708 7748
rect 11116 7708 11156 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 5548 7372 5588 7412
rect 844 7204 884 7244
rect 5260 7120 5300 7160
rect 5356 7120 5396 7160
rect 5548 7120 5588 7160
rect 11692 7120 11732 7160
rect 12076 7120 12116 7160
rect 12940 7120 12980 7160
rect 652 6952 692 6992
rect 14092 6952 14132 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 4780 6448 4820 6488
rect 4972 6448 5012 6488
rect 2860 6364 2900 6404
rect 2668 6196 2708 6236
rect 4876 6196 4916 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 844 5692 884 5732
rect 4972 5608 5012 5648
rect 652 5440 692 5480
rect 4300 5440 4340 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 4012 5104 4052 5144
rect 3820 4936 3860 4976
rect 3916 4936 3956 4976
rect 4108 4936 4148 4976
rect 4300 4936 4340 4976
rect 4492 4936 4532 4976
rect 9196 4936 9236 4976
rect 9292 4936 9332 4976
rect 9388 4936 9428 4976
rect 9484 4936 9524 4976
rect 844 4852 884 4892
rect 2860 4852 2900 4892
rect 652 4768 692 4808
rect 2668 4768 2708 4808
rect 4492 4684 4532 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 2668 4264 2708 4304
rect 5164 4264 5204 4304
rect 844 4180 884 4220
rect 2860 4180 2900 4220
rect 4780 4096 4820 4136
rect 5836 4096 5876 4136
rect 9292 4096 9332 4136
rect 9484 4096 9524 4136
rect 9580 4096 9620 4136
rect 10636 4096 10676 4136
rect 11308 4096 11348 4136
rect 652 3928 692 3968
rect 4108 3928 4148 3968
rect 9388 3928 9428 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 11596 3592 11636 3632
rect 9196 3508 9236 3548
rect 9580 3424 9620 3464
rect 10444 3424 10484 3464
rect 844 3340 884 3380
rect 4108 3256 4148 3296
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 6028 2836 6068 2876
rect 2668 2752 2708 2792
rect 9676 2752 9716 2792
rect 844 2668 884 2708
rect 2860 2668 2900 2708
rect 3628 2584 3668 2624
rect 4012 2584 4052 2624
rect 4876 2584 4916 2624
rect 652 2416 692 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 652 38156 692 38165
rect 652 37577 692 38116
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 2187 37988 2229 37997
rect 2187 37948 2188 37988
rect 2228 37948 2229 37988
rect 2187 37939 2229 37948
rect 844 37854 884 37939
rect 651 37568 693 37577
rect 651 37528 652 37568
rect 692 37528 693 37568
rect 651 37519 693 37528
rect 652 23036 692 23045
rect 556 22996 652 23036
rect 556 22457 596 22996
rect 652 22987 692 22996
rect 844 22868 884 22877
rect 555 22448 597 22457
rect 555 22408 556 22448
rect 596 22408 597 22448
rect 555 22399 597 22408
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 844 20777 884 22828
rect 2188 20945 2228 37939
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 9867 36728 9909 36737
rect 9867 36688 9868 36728
rect 9908 36688 9909 36728
rect 9867 36679 9909 36688
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3531 21692 3573 21701
rect 3531 21652 3532 21692
rect 3572 21652 3573 21692
rect 3531 21643 3573 21652
rect 4971 21692 5013 21701
rect 4971 21652 4972 21692
rect 5012 21652 5013 21692
rect 4971 21643 5013 21652
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 3244 21020 3284 21029
rect 3532 21020 3572 21643
rect 4972 21558 5012 21643
rect 5356 21608 5396 21617
rect 3284 20980 3572 21020
rect 3244 20971 3284 20980
rect 2187 20936 2229 20945
rect 2187 20896 2188 20936
rect 2228 20896 2229 20936
rect 2187 20887 2229 20896
rect 2763 20936 2805 20945
rect 2763 20896 2764 20936
rect 2804 20896 2805 20936
rect 2763 20887 2805 20896
rect 3723 20936 3765 20945
rect 3723 20896 3724 20936
rect 3764 20896 3765 20936
rect 3723 20887 3765 20896
rect 5356 20936 5396 21568
rect 6219 21608 6261 21617
rect 6219 21568 6220 21608
rect 6260 21568 6261 21608
rect 6219 21559 6261 21568
rect 8907 21608 8949 21617
rect 8907 21568 8908 21608
rect 8948 21568 8949 21608
rect 8907 21559 8949 21568
rect 6220 21474 6260 21559
rect 6219 21356 6261 21365
rect 6219 21316 6220 21356
rect 6260 21316 6261 21356
rect 6219 21307 6261 21316
rect 7371 21356 7413 21365
rect 7371 21316 7372 21356
rect 7412 21316 7413 21356
rect 7371 21307 7413 21316
rect 5356 20887 5396 20896
rect 2667 20852 2709 20861
rect 2667 20812 2668 20852
rect 2708 20812 2709 20852
rect 2667 20803 2709 20812
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 843 20768 885 20777
rect 843 20728 844 20768
rect 884 20728 885 20768
rect 843 20719 885 20728
rect 2379 20768 2421 20777
rect 2379 20728 2380 20768
rect 2420 20728 2421 20768
rect 2379 20719 2421 20728
rect 2571 20768 2613 20777
rect 2571 20728 2572 20768
rect 2612 20728 2613 20768
rect 2571 20719 2613 20728
rect 2668 20768 2708 20803
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19794 692 19879
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 652 15737 692 16360
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 844 15476 884 15485
rect 652 15308 692 15317
rect 652 14897 692 15268
rect 844 15233 884 15436
rect 843 15224 885 15233
rect 843 15184 844 15224
rect 884 15184 885 15224
rect 843 15175 885 15184
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 843 14804 885 14813
rect 843 14764 844 14804
rect 884 14764 885 14804
rect 843 14755 885 14764
rect 2187 14804 2229 14813
rect 2187 14764 2188 14804
rect 2228 14764 2229 14804
rect 2187 14755 2229 14764
rect 844 14670 884 14755
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 843 13292 885 13301
rect 843 13252 844 13292
rect 884 13252 885 13292
rect 843 13243 885 13252
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 844 13158 884 13243
rect 652 12991 692 13000
rect 843 12452 885 12461
rect 843 12412 844 12452
rect 884 12412 885 12452
rect 843 12403 885 12412
rect 2091 12452 2133 12461
rect 2091 12412 2092 12452
rect 2132 12412 2133 12452
rect 2091 12403 2133 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 652 12234 692 12319
rect 844 12318 884 12403
rect 844 11780 884 11789
rect 884 11740 1076 11780
rect 844 11731 884 11740
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 843 10940 885 10949
rect 843 10900 844 10940
rect 884 10900 885 10940
rect 843 10891 885 10900
rect 844 10806 884 10891
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 652 10638 692 10723
rect 843 10268 885 10277
rect 843 10228 844 10268
rect 884 10228 885 10268
rect 843 10219 885 10228
rect 844 10134 884 10219
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 843 9428 885 9437
rect 843 9388 844 9428
rect 884 9388 885 9428
rect 843 9379 885 9388
rect 844 9294 884 9379
rect 652 9260 692 9269
rect 652 9017 692 9220
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 747 8840 789 8849
rect 747 8800 748 8840
rect 788 8800 789 8840
rect 747 8791 789 8800
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 652 7748 692 7757
rect 652 7337 692 7708
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 748 7244 788 8791
rect 843 8756 885 8765
rect 843 8716 844 8756
rect 884 8716 885 8756
rect 843 8707 885 8716
rect 844 8622 884 8707
rect 939 8672 981 8681
rect 939 8632 940 8672
rect 980 8632 981 8672
rect 939 8623 981 8632
rect 844 7916 884 7925
rect 940 7916 980 8623
rect 884 7876 980 7916
rect 844 7867 884 7876
rect 939 7748 981 7757
rect 939 7708 940 7748
rect 980 7708 981 7748
rect 939 7699 981 7708
rect 844 7244 884 7253
rect 748 7204 844 7244
rect 844 7195 884 7204
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 843 6236 885 6245
rect 843 6196 844 6236
rect 884 6196 885 6236
rect 843 6187 885 6196
rect 844 5732 884 6187
rect 844 5683 884 5692
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 844 4892 884 4903
rect 844 4817 884 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 843 4808 885 4817
rect 843 4768 844 4808
rect 884 4768 885 4808
rect 843 4759 885 4768
rect 652 4674 692 4759
rect 843 4304 885 4313
rect 843 4264 844 4304
rect 884 4264 885 4304
rect 843 4255 885 4264
rect 844 4220 884 4255
rect 844 4169 884 4180
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 844 3380 884 3389
rect 940 3380 980 7699
rect 1036 4901 1076 11740
rect 1131 10940 1173 10949
rect 1131 10900 1132 10940
rect 1172 10900 1173 10940
rect 1131 10891 1173 10900
rect 1035 4892 1077 4901
rect 1035 4852 1036 4892
rect 1076 4852 1077 4892
rect 1035 4843 1077 4852
rect 1132 4397 1172 10891
rect 2092 6413 2132 12403
rect 2188 12209 2228 14755
rect 2187 12200 2229 12209
rect 2187 12160 2188 12200
rect 2228 12160 2229 12200
rect 2187 12151 2229 12160
rect 2188 8933 2228 12151
rect 2283 11780 2325 11789
rect 2283 11740 2284 11780
rect 2324 11740 2325 11780
rect 2283 11731 2325 11740
rect 2284 11696 2324 11731
rect 2284 9437 2324 11656
rect 2380 11696 2420 20719
rect 2572 20634 2612 20719
rect 2668 20717 2708 20728
rect 2764 20768 2804 20887
rect 2764 20719 2804 20728
rect 2859 20768 2901 20777
rect 2859 20728 2860 20768
rect 2900 20728 2901 20768
rect 2859 20719 2901 20728
rect 3243 20768 3285 20777
rect 3243 20728 3244 20768
rect 3284 20728 3285 20768
rect 3243 20719 3285 20728
rect 3436 20768 3476 20779
rect 2860 20634 2900 20719
rect 3244 20634 3284 20719
rect 3436 20693 3476 20728
rect 3531 20768 3573 20777
rect 3531 20728 3532 20768
rect 3572 20728 3573 20768
rect 3531 20719 3573 20728
rect 3435 20684 3477 20693
rect 3435 20644 3436 20684
rect 3476 20644 3477 20684
rect 3435 20635 3477 20644
rect 3532 20634 3572 20719
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 3724 16157 3764 20887
rect 5547 20768 5589 20777
rect 5547 20728 5548 20768
rect 5588 20728 5589 20768
rect 5547 20719 5589 20728
rect 6220 20768 6260 21307
rect 7372 21222 7412 21307
rect 5548 20634 5588 20719
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3723 16148 3765 16157
rect 3723 16108 3724 16148
rect 3764 16108 3765 16148
rect 3723 16099 3765 16108
rect 4107 16148 4149 16157
rect 4107 16108 4108 16148
rect 4148 16108 4149 16148
rect 4107 16099 4149 16108
rect 2859 15224 2901 15233
rect 2859 15184 2860 15224
rect 2900 15184 2901 15224
rect 2859 15175 2901 15184
rect 2764 13796 2804 13805
rect 2475 13292 2517 13301
rect 2475 13252 2476 13292
rect 2516 13252 2517 13292
rect 2475 13243 2517 13252
rect 2476 11957 2516 13243
rect 2764 13217 2804 13756
rect 2763 13208 2805 13217
rect 2763 13168 2764 13208
rect 2804 13168 2805 13208
rect 2763 13159 2805 13168
rect 2475 11948 2517 11957
rect 2475 11908 2476 11948
rect 2516 11908 2517 11948
rect 2475 11899 2517 11908
rect 2380 11537 2420 11656
rect 2379 11528 2421 11537
rect 2379 11488 2380 11528
rect 2420 11488 2421 11528
rect 2379 11479 2421 11488
rect 2283 9428 2325 9437
rect 2283 9388 2284 9428
rect 2324 9388 2420 9428
rect 2283 9379 2325 9388
rect 2187 8924 2229 8933
rect 2187 8884 2188 8924
rect 2228 8884 2229 8924
rect 2187 8875 2229 8884
rect 2283 8840 2325 8849
rect 2283 8800 2284 8840
rect 2324 8800 2325 8840
rect 2283 8791 2325 8800
rect 2284 8706 2324 8791
rect 2380 7220 2420 9388
rect 2476 8756 2516 11899
rect 2572 11873 2612 11958
rect 2571 11864 2613 11873
rect 2571 11824 2572 11864
rect 2612 11824 2613 11864
rect 2571 11815 2613 11824
rect 2571 11696 2613 11705
rect 2571 11656 2572 11696
rect 2612 11656 2613 11696
rect 2571 11647 2613 11656
rect 2572 11562 2612 11647
rect 2764 10277 2804 13159
rect 2763 10268 2805 10277
rect 2763 10228 2764 10268
rect 2804 10228 2805 10268
rect 2763 10219 2805 10228
rect 2668 9260 2708 9269
rect 2668 8765 2708 9220
rect 2476 8707 2516 8716
rect 2667 8756 2709 8765
rect 2667 8716 2668 8756
rect 2708 8716 2709 8756
rect 2667 8707 2709 8716
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 2572 8504 2612 8623
rect 2668 8504 2708 8513
rect 2572 8464 2668 8504
rect 2668 8455 2708 8464
rect 2764 7916 2804 10219
rect 2860 9428 2900 15175
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 3915 14048 3957 14057
rect 3915 14008 3916 14048
rect 3956 14008 3957 14048
rect 3915 13999 3957 14008
rect 3916 13914 3956 13999
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4011 13376 4053 13385
rect 4011 13336 4012 13376
rect 4052 13336 4053 13376
rect 4011 13327 4053 13336
rect 4012 13242 4052 13327
rect 3627 13208 3669 13217
rect 3627 13168 3628 13208
rect 3668 13168 3669 13208
rect 3627 13159 3669 13168
rect 3628 13074 3668 13159
rect 2956 13040 2996 13049
rect 2956 11705 2996 13000
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3435 11864 3477 11873
rect 4108 11864 4148 16099
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4780 14048 4820 14057
rect 5164 14048 5204 14057
rect 4780 13385 4820 14008
rect 4876 14008 5164 14048
rect 4779 13376 4821 13385
rect 4779 13336 4780 13376
rect 4820 13336 4821 13376
rect 4779 13327 4821 13336
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4876 12704 4916 14008
rect 5164 13999 5204 14008
rect 3435 11824 3436 11864
rect 3476 11824 3477 11864
rect 3435 11815 3477 11824
rect 4012 11824 4148 11864
rect 4492 12664 4916 12704
rect 4492 11864 4532 12664
rect 3051 11780 3093 11789
rect 3051 11740 3052 11780
rect 3092 11740 3093 11780
rect 3051 11731 3093 11740
rect 2955 11696 2997 11705
rect 2955 11656 2956 11696
rect 2996 11656 2997 11696
rect 2955 11647 2997 11656
rect 3052 11696 3092 11731
rect 3052 11645 3092 11656
rect 3243 11696 3285 11705
rect 3243 11656 3244 11696
rect 3284 11656 3285 11696
rect 3243 11647 3285 11656
rect 3436 11696 3476 11815
rect 3436 11647 3476 11656
rect 3244 11612 3284 11647
rect 3244 11561 3284 11572
rect 2955 11528 2997 11537
rect 2955 11488 2956 11528
rect 2996 11488 2997 11528
rect 2955 11479 2997 11488
rect 2956 11394 2996 11479
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 4012 9512 4052 11824
rect 4492 11815 4532 11824
rect 6220 11789 6260 20728
rect 7948 17872 8180 17912
rect 7660 17744 7700 17753
rect 7948 17744 7988 17872
rect 7700 17704 7988 17744
rect 8044 17744 8084 17753
rect 7660 17695 7700 17704
rect 8044 17300 8084 17704
rect 7948 17260 8084 17300
rect 7948 16904 7988 17260
rect 8140 17240 8180 17872
rect 8140 17191 8180 17200
rect 8908 17744 8948 21559
rect 7948 16855 7988 16864
rect 8812 17072 8852 17081
rect 8428 16493 8468 16578
rect 8812 16493 8852 17032
rect 8427 16484 8469 16493
rect 8427 16444 8428 16484
rect 8468 16444 8469 16484
rect 8427 16435 8469 16444
rect 8811 16484 8853 16493
rect 8811 16444 8812 16484
rect 8852 16444 8853 16484
rect 8811 16435 8853 16444
rect 8428 16232 8468 16241
rect 8428 16073 8468 16192
rect 8619 16232 8661 16241
rect 8619 16192 8620 16232
rect 8660 16192 8661 16232
rect 8619 16183 8661 16192
rect 8716 16232 8756 16241
rect 8908 16232 8948 17704
rect 9484 16820 9524 16829
rect 9196 16780 9484 16820
rect 8620 16098 8660 16183
rect 8427 16064 8469 16073
rect 8427 16024 8428 16064
rect 8468 16024 8469 16064
rect 8427 16015 8469 16024
rect 8716 15560 8756 16192
rect 8812 16192 8948 16232
rect 9004 16232 9044 16243
rect 9196 16241 9236 16780
rect 9484 16771 9524 16780
rect 8812 15728 8852 16192
rect 9004 16157 9044 16192
rect 9100 16232 9140 16241
rect 9003 16148 9045 16157
rect 9003 16108 9004 16148
rect 9044 16108 9045 16148
rect 9003 16099 9045 16108
rect 8907 16064 8949 16073
rect 8907 16024 8908 16064
rect 8948 16024 8949 16064
rect 8907 16015 8949 16024
rect 8908 15930 8948 16015
rect 9004 15728 9044 15737
rect 8812 15688 9004 15728
rect 9004 15679 9044 15688
rect 9100 15560 9140 16192
rect 9195 16232 9237 16241
rect 9195 16192 9196 16232
rect 9236 16192 9237 16232
rect 9195 16183 9237 16192
rect 9196 16098 9236 16183
rect 8716 15520 9140 15560
rect 8907 11948 8949 11957
rect 8907 11908 8908 11948
rect 8948 11908 8949 11948
rect 8907 11899 8949 11908
rect 8524 11864 8564 11875
rect 8524 11789 8564 11824
rect 6219 11780 6261 11789
rect 6219 11740 6220 11780
rect 6260 11740 6261 11780
rect 6219 11731 6261 11740
rect 8523 11780 8565 11789
rect 8523 11740 8524 11780
rect 8564 11740 8565 11780
rect 8523 11731 8565 11740
rect 4108 11696 4148 11705
rect 4300 11696 4340 11705
rect 4148 11656 4300 11696
rect 4108 11647 4148 11656
rect 4300 11647 4340 11656
rect 4395 11696 4437 11705
rect 4395 11656 4396 11696
rect 4436 11656 4437 11696
rect 4395 11647 4437 11656
rect 4588 11696 4628 11705
rect 8716 11696 8756 11705
rect 4628 11656 4820 11696
rect 4588 11647 4628 11656
rect 4396 11562 4436 11647
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4780 10025 4820 11656
rect 8716 11033 8756 11656
rect 8811 11696 8853 11705
rect 8811 11656 8812 11696
rect 8852 11656 8853 11696
rect 8811 11647 8853 11656
rect 8908 11696 8948 11899
rect 9100 11789 9140 15520
rect 9580 15476 9620 15485
rect 9580 14729 9620 15436
rect 9579 14720 9621 14729
rect 9579 14680 9580 14720
rect 9620 14680 9621 14720
rect 9579 14671 9621 14680
rect 9580 14057 9620 14671
rect 9579 14048 9621 14057
rect 9579 14008 9580 14048
rect 9620 14008 9621 14048
rect 9579 13999 9621 14008
rect 9675 12956 9717 12965
rect 9675 12916 9676 12956
rect 9716 12916 9717 12956
rect 9675 12907 9717 12916
rect 9099 11780 9141 11789
rect 9099 11740 9100 11780
rect 9140 11740 9141 11780
rect 9099 11731 9141 11740
rect 8908 11647 8948 11656
rect 9003 11696 9045 11705
rect 9676 11696 9716 12907
rect 9868 12536 9908 36679
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 10060 17576 10100 17585
rect 10060 17072 10100 17536
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 10156 17072 10196 17100
rect 10060 17032 10156 17072
rect 10060 15233 10100 17032
rect 10156 17023 10196 17032
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 10251 16148 10293 16157
rect 10251 16108 10252 16148
rect 10292 16108 10293 16148
rect 10251 16099 10293 16108
rect 10059 15224 10101 15233
rect 10059 15184 10060 15224
rect 10100 15184 10101 15224
rect 10059 15175 10101 15184
rect 10155 13208 10197 13217
rect 10155 13168 10156 13208
rect 10196 13168 10197 13208
rect 10155 13159 10197 13168
rect 10252 13208 10292 16099
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 10924 15560 10964 15569
rect 10443 14048 10485 14057
rect 10443 14008 10444 14048
rect 10484 14008 10485 14048
rect 10443 13999 10485 14008
rect 10252 13159 10292 13168
rect 10348 13208 10388 13217
rect 10156 13074 10196 13159
rect 10348 12965 10388 13168
rect 10444 13208 10484 13999
rect 10444 13159 10484 13168
rect 10347 12956 10389 12965
rect 10347 12916 10348 12956
rect 10388 12916 10389 12956
rect 10347 12907 10389 12916
rect 9868 12487 9908 12496
rect 10924 12452 10964 15520
rect 13612 15392 13652 15401
rect 13516 15352 13612 15392
rect 13516 14720 13556 15352
rect 13612 15343 13652 15352
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 13516 14671 13556 14680
rect 14379 14720 14421 14729
rect 14379 14680 14380 14720
rect 14420 14680 14421 14720
rect 14379 14671 14421 14680
rect 13132 14636 13172 14645
rect 13132 14225 13172 14596
rect 14380 14586 14420 14671
rect 15532 14552 15572 14561
rect 11307 14216 11349 14225
rect 11307 14176 11308 14216
rect 11348 14176 11349 14216
rect 11307 14167 11349 14176
rect 13131 14216 13173 14225
rect 13131 14176 13132 14216
rect 13172 14176 13173 14216
rect 13131 14167 13173 14176
rect 11308 14082 11348 14167
rect 15532 14057 15572 14512
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 11116 14048 11156 14057
rect 11116 12965 11156 14008
rect 11211 14048 11253 14057
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 11404 14048 11444 14057
rect 11212 13914 11252 13999
rect 11404 13217 11444 14008
rect 13515 14048 13557 14057
rect 13515 14008 13516 14048
rect 13556 14008 13557 14048
rect 13515 13999 13557 14008
rect 14187 14048 14229 14057
rect 14187 14008 14188 14048
rect 14228 14008 14229 14048
rect 14187 13999 14229 14008
rect 15531 14048 15573 14057
rect 15531 14008 15532 14048
rect 15572 14008 15573 14048
rect 15531 13999 15573 14008
rect 13516 13914 13556 13999
rect 11403 13208 11445 13217
rect 11403 13168 11404 13208
rect 11444 13168 11445 13208
rect 11403 13159 11445 13168
rect 11115 12956 11157 12965
rect 11115 12916 11116 12956
rect 11156 12916 11157 12956
rect 11115 12907 11157 12916
rect 11308 12452 11348 12461
rect 10924 12412 11308 12452
rect 9771 11948 9813 11957
rect 9771 11908 9772 11948
rect 9812 11908 9813 11948
rect 9771 11899 9813 11908
rect 9003 11656 9004 11696
rect 9044 11656 9045 11696
rect 9003 11647 9045 11656
rect 9484 11656 9676 11696
rect 8812 11562 8852 11647
rect 9004 11562 9044 11647
rect 9195 11612 9237 11621
rect 9195 11572 9196 11612
rect 9236 11572 9237 11612
rect 9195 11563 9237 11572
rect 9196 11192 9236 11563
rect 9100 11152 9196 11192
rect 8715 11024 8757 11033
rect 8715 10984 8716 11024
rect 8756 10984 8757 11024
rect 8715 10975 8757 10984
rect 4203 10016 4245 10025
rect 4203 9976 4204 10016
rect 4244 9976 4245 10016
rect 4203 9967 4245 9976
rect 4779 10016 4821 10025
rect 4779 9976 4780 10016
rect 4820 9976 4821 10016
rect 4779 9967 4821 9976
rect 4204 9680 4244 9967
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4204 9631 4244 9640
rect 4107 9512 4149 9521
rect 4012 9472 4108 9512
rect 4148 9472 4149 9512
rect 4107 9463 4149 9472
rect 4779 9512 4821 9521
rect 4779 9472 4780 9512
rect 4820 9472 4821 9512
rect 4779 9463 4821 9472
rect 2860 9379 2900 9388
rect 4108 9378 4148 9463
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 2859 8924 2901 8933
rect 2859 8884 2860 8924
rect 2900 8884 2901 8924
rect 2859 8875 2901 8884
rect 2860 8756 2900 8875
rect 2860 8707 2900 8716
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 2860 7916 2900 7925
rect 2764 7876 2860 7916
rect 2860 7867 2900 7876
rect 2667 7748 2709 7757
rect 2667 7708 2668 7748
rect 2708 7708 2709 7748
rect 2667 7699 2709 7708
rect 2668 7614 2708 7699
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 2380 7180 2804 7220
rect 2091 6404 2133 6413
rect 2091 6364 2092 6404
rect 2132 6364 2133 6404
rect 2091 6355 2133 6364
rect 2667 6236 2709 6245
rect 2667 6196 2668 6236
rect 2708 6196 2709 6236
rect 2667 6187 2709 6196
rect 2668 6102 2708 6187
rect 2667 4808 2709 4817
rect 2667 4768 2668 4808
rect 2708 4768 2709 4808
rect 2667 4759 2709 4768
rect 2668 4674 2708 4759
rect 1131 4388 1173 4397
rect 1131 4348 1132 4388
rect 1172 4348 1173 4388
rect 1131 4339 1173 4348
rect 2667 4304 2709 4313
rect 2667 4264 2668 4304
rect 2708 4264 2709 4304
rect 2667 4255 2709 4264
rect 2668 4170 2708 4255
rect 884 3340 980 3380
rect 844 3331 884 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 843 2792 885 2801
rect 843 2752 844 2792
rect 884 2752 885 2792
rect 843 2743 885 2752
rect 2667 2792 2709 2801
rect 2667 2752 2668 2792
rect 2708 2752 2709 2792
rect 2667 2743 2709 2752
rect 844 2708 884 2743
rect 844 2657 884 2668
rect 2668 2658 2708 2743
rect 2764 2708 2804 7180
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 4780 6497 4820 9463
rect 5355 8840 5397 8849
rect 5355 8800 5356 8840
rect 5396 8800 5397 8840
rect 5355 8791 5397 8800
rect 7179 8840 7221 8849
rect 7179 8800 7180 8840
rect 7220 8800 7221 8840
rect 7179 8791 7221 8800
rect 7371 8840 7413 8849
rect 7371 8800 7372 8840
rect 7412 8800 7413 8840
rect 7371 8791 7413 8800
rect 4971 7412 5013 7421
rect 4971 7372 4972 7412
rect 5012 7372 5013 7412
rect 4971 7363 5013 7372
rect 4779 6488 4821 6497
rect 4779 6448 4780 6488
rect 4820 6448 4821 6488
rect 4779 6439 4821 6448
rect 4972 6488 5012 7363
rect 4972 6439 5012 6448
rect 5260 7160 5300 7169
rect 2859 6404 2901 6413
rect 2859 6364 2860 6404
rect 2900 6364 2901 6404
rect 2859 6355 2901 6364
rect 2860 6270 2900 6355
rect 4780 6354 4820 6439
rect 4876 6236 4916 6245
rect 4780 6196 4876 6236
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4300 5480 4340 5489
rect 4204 5440 4300 5480
rect 4011 5144 4053 5153
rect 4011 5104 4012 5144
rect 4052 5104 4053 5144
rect 4204 5144 4244 5440
rect 4300 5431 4340 5440
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 4204 5104 4340 5144
rect 4011 5095 4053 5104
rect 4012 5010 4052 5095
rect 3819 4976 3861 4985
rect 3819 4936 3820 4976
rect 3860 4936 3861 4976
rect 3819 4927 3861 4936
rect 3916 4976 3956 4985
rect 2859 4892 2901 4901
rect 2859 4852 2860 4892
rect 2900 4852 2901 4892
rect 2859 4843 2901 4852
rect 2860 4758 2900 4843
rect 3820 4842 3860 4927
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 3916 4397 3956 4936
rect 4108 4976 4148 4985
rect 4108 4481 4148 4936
rect 4300 4976 4340 5104
rect 4300 4927 4340 4936
rect 4492 4976 4532 4985
rect 4780 4976 4820 6196
rect 4876 6187 4916 6196
rect 4972 5648 5012 5657
rect 4972 5153 5012 5608
rect 4971 5144 5013 5153
rect 4971 5104 4972 5144
rect 5012 5104 5013 5144
rect 4971 5095 5013 5104
rect 5260 4985 5300 7120
rect 5356 7160 5396 8791
rect 7084 8681 7124 8766
rect 7180 8697 7220 8791
rect 7372 8706 7412 8791
rect 5643 8672 5685 8681
rect 5643 8632 5644 8672
rect 5684 8632 5685 8672
rect 5643 8623 5685 8632
rect 7083 8672 7125 8681
rect 7083 8632 7084 8672
rect 7124 8632 7125 8672
rect 7180 8648 7220 8657
rect 8715 8672 8757 8681
rect 7083 8623 7125 8632
rect 8715 8632 8716 8672
rect 8756 8632 8757 8672
rect 8715 8623 8757 8632
rect 5547 7412 5589 7421
rect 5547 7372 5548 7412
rect 5588 7372 5589 7412
rect 5547 7363 5589 7372
rect 5548 7278 5588 7363
rect 4532 4936 4820 4976
rect 5259 4976 5301 4985
rect 5259 4936 5260 4976
rect 5300 4936 5301 4976
rect 4492 4927 4532 4936
rect 5259 4927 5301 4936
rect 4492 4724 4532 4733
rect 4532 4684 4820 4724
rect 4492 4675 4532 4684
rect 4107 4472 4149 4481
rect 4107 4432 4108 4472
rect 4148 4432 4149 4472
rect 4107 4423 4149 4432
rect 2859 4388 2901 4397
rect 2859 4348 2860 4388
rect 2900 4348 2901 4388
rect 2859 4339 2901 4348
rect 3915 4388 3957 4397
rect 3915 4348 3916 4388
rect 3956 4348 3957 4388
rect 3915 4339 3957 4348
rect 2860 4220 2900 4339
rect 2860 4171 2900 4180
rect 4780 4136 4820 4684
rect 5163 4472 5205 4481
rect 5163 4432 5164 4472
rect 5204 4432 5205 4472
rect 5163 4423 5205 4432
rect 5164 4304 5204 4423
rect 5356 4313 5396 7120
rect 5548 7160 5588 7169
rect 5644 7160 5684 8623
rect 7084 8504 7124 8513
rect 7084 8093 7124 8464
rect 8428 8093 8468 8124
rect 7083 8084 7125 8093
rect 7083 8044 7084 8084
rect 7124 8044 7125 8084
rect 7083 8035 7125 8044
rect 8427 8084 8469 8093
rect 8427 8044 8428 8084
rect 8468 8044 8469 8084
rect 8427 8035 8469 8044
rect 8428 8000 8468 8035
rect 8428 7925 8468 7960
rect 8523 8000 8565 8009
rect 8523 7960 8524 8000
rect 8564 7960 8565 8000
rect 8523 7951 8565 7960
rect 8716 8000 8756 8623
rect 8716 7951 8756 7960
rect 8811 8000 8853 8009
rect 8811 7960 8812 8000
rect 8852 7960 8853 8000
rect 8811 7951 8853 7960
rect 9004 8000 9044 8009
rect 8427 7916 8469 7925
rect 8427 7876 8428 7916
rect 8468 7876 8469 7916
rect 8427 7867 8469 7876
rect 8524 7866 8564 7951
rect 8812 7866 8852 7951
rect 9004 7421 9044 7960
rect 9100 8000 9140 11152
rect 9196 11143 9236 11152
rect 9484 11192 9524 11656
rect 9676 11647 9716 11656
rect 9772 11696 9812 11899
rect 9964 11873 10004 11958
rect 9963 11864 10005 11873
rect 9963 11824 9964 11864
rect 10004 11824 10005 11864
rect 9963 11815 10005 11824
rect 10827 11864 10869 11873
rect 10827 11824 10828 11864
rect 10868 11824 10869 11864
rect 10827 11815 10869 11824
rect 9867 11780 9909 11789
rect 9867 11740 9868 11780
rect 9908 11740 9909 11780
rect 9867 11731 9909 11740
rect 9772 11647 9812 11656
rect 9868 11444 9908 11731
rect 9963 11696 10005 11705
rect 9963 11656 9964 11696
rect 10004 11656 10005 11696
rect 9963 11647 10005 11656
rect 10828 11696 10868 11815
rect 10828 11647 10868 11656
rect 9964 11562 10004 11647
rect 10156 11612 10196 11621
rect 10060 11572 10156 11612
rect 9868 11404 10004 11444
rect 9484 11143 9524 11152
rect 9771 11192 9813 11201
rect 9771 11152 9772 11192
rect 9812 11152 9813 11192
rect 9771 11143 9813 11152
rect 9772 11058 9812 11143
rect 9291 11024 9333 11033
rect 9291 10984 9292 11024
rect 9332 10984 9333 11024
rect 9291 10975 9333 10984
rect 9676 11024 9716 11033
rect 9292 8849 9332 10975
rect 9676 10025 9716 10984
rect 9868 11024 9908 11033
rect 9868 10856 9908 10984
rect 9964 11024 10004 11404
rect 9964 10975 10004 10984
rect 10060 10856 10100 11572
rect 10156 11563 10196 11572
rect 9868 10816 10100 10856
rect 9675 10016 9717 10025
rect 9675 9976 9676 10016
rect 9716 9976 9717 10016
rect 9675 9967 9717 9976
rect 9291 8840 9333 8849
rect 9291 8800 9292 8840
rect 9332 8800 9333 8840
rect 9291 8791 9333 8800
rect 9196 8177 9236 8262
rect 9195 8168 9237 8177
rect 9195 8128 9196 8168
rect 9236 8128 9237 8168
rect 9195 8119 9237 8128
rect 9292 8009 9332 8791
rect 9676 8681 9716 9967
rect 10540 9512 10580 9521
rect 11308 9512 11348 12412
rect 14091 12200 14133 12209
rect 14091 12160 14092 12200
rect 14132 12160 14133 12200
rect 14091 12151 14133 12160
rect 14092 11705 14132 12151
rect 14188 11957 14228 13999
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 14187 11948 14229 11957
rect 14187 11908 14188 11948
rect 14228 11908 14229 11948
rect 14187 11899 14229 11908
rect 12076 11696 12116 11705
rect 12076 11201 12116 11656
rect 13419 11696 13461 11705
rect 13419 11656 13420 11696
rect 13460 11656 13461 11696
rect 13419 11647 13461 11656
rect 14091 11696 14133 11705
rect 14091 11656 14092 11696
rect 14132 11656 14133 11696
rect 14091 11647 14133 11656
rect 16491 11696 16533 11705
rect 16491 11656 16492 11696
rect 16532 11656 16533 11696
rect 16491 11647 16533 11656
rect 12747 11612 12789 11621
rect 12747 11572 12748 11612
rect 12788 11572 12789 11612
rect 12747 11563 12789 11572
rect 12748 11478 12788 11563
rect 13420 11562 13460 11647
rect 13995 11612 14037 11621
rect 13995 11572 13996 11612
rect 14036 11572 14037 11612
rect 13995 11563 14037 11572
rect 12075 11192 12117 11201
rect 12075 11152 12076 11192
rect 12116 11152 12117 11192
rect 12075 11143 12117 11152
rect 13996 11108 14036 11563
rect 14092 11562 14132 11647
rect 16492 11192 16532 11647
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 16492 11143 16532 11152
rect 14092 11108 14132 11117
rect 13996 11068 14092 11108
rect 14092 11059 14132 11068
rect 14476 11024 14516 11033
rect 14476 10352 14516 10984
rect 15340 11024 15380 11033
rect 14572 10352 14612 10361
rect 14476 10312 14572 10352
rect 14572 10303 14612 10312
rect 15340 9689 15380 10984
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 12459 9680 12501 9689
rect 12459 9640 12460 9680
rect 12500 9640 12501 9680
rect 12459 9631 12501 9640
rect 12939 9680 12981 9689
rect 12939 9640 12940 9680
rect 12980 9640 12981 9680
rect 12939 9631 12981 9640
rect 15339 9680 15381 9689
rect 15339 9640 15340 9680
rect 15380 9640 15381 9680
rect 15339 9631 15381 9640
rect 12460 9546 12500 9631
rect 10580 9472 11348 9512
rect 10540 9463 10580 9472
rect 12940 8681 12980 9631
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 9675 8672 9717 8681
rect 9675 8632 9676 8672
rect 9716 8632 9717 8672
rect 9675 8623 9717 8632
rect 10539 8672 10581 8681
rect 10539 8632 10540 8672
rect 10580 8632 10581 8672
rect 10539 8623 10581 8632
rect 12939 8672 12981 8681
rect 12939 8632 12940 8672
rect 12980 8632 12981 8672
rect 12939 8623 12981 8632
rect 10443 8168 10485 8177
rect 10443 8128 10444 8168
rect 10484 8128 10485 8168
rect 10443 8119 10485 8128
rect 9003 7412 9045 7421
rect 9003 7372 9004 7412
rect 9044 7372 9045 7412
rect 9003 7363 9045 7372
rect 5588 7120 5684 7160
rect 5548 4481 5588 7120
rect 9100 4985 9140 7960
rect 9255 8000 9332 8009
rect 9295 7960 9332 8000
rect 10444 8000 10484 8119
rect 9255 7951 9295 7960
rect 10444 7951 10484 7960
rect 10540 7220 10580 8623
rect 12076 8000 12116 8009
rect 11980 7960 12076 8000
rect 11403 7916 11445 7925
rect 11403 7876 11404 7916
rect 11444 7876 11445 7916
rect 11403 7867 11445 7876
rect 11404 7782 11444 7867
rect 11115 7748 11157 7757
rect 11115 7708 11116 7748
rect 11156 7708 11157 7748
rect 11115 7699 11157 7708
rect 11691 7748 11733 7757
rect 11691 7708 11692 7748
rect 11732 7708 11733 7748
rect 11691 7699 11733 7708
rect 11116 7614 11156 7699
rect 10444 7180 10580 7220
rect 9291 6488 9333 6497
rect 9291 6448 9292 6488
rect 9332 6448 9333 6488
rect 9291 6439 9333 6448
rect 9099 4976 9141 4985
rect 9099 4936 9100 4976
rect 9140 4936 9141 4976
rect 9099 4927 9141 4936
rect 9196 4976 9236 4985
rect 5835 4892 5877 4901
rect 5835 4852 5836 4892
rect 5876 4852 5877 4892
rect 5835 4843 5877 4852
rect 5547 4472 5589 4481
rect 5547 4432 5548 4472
rect 5588 4432 5589 4472
rect 5547 4423 5589 4432
rect 5164 4255 5204 4264
rect 5355 4304 5397 4313
rect 5355 4264 5356 4304
rect 5396 4264 5397 4304
rect 5355 4255 5397 4264
rect 4780 4087 4820 4096
rect 5836 4136 5876 4843
rect 9196 4136 9236 4936
rect 9292 4976 9332 6439
rect 9292 4927 9332 4936
rect 9387 4976 9429 4985
rect 9387 4936 9388 4976
rect 9428 4936 9429 4976
rect 9387 4927 9429 4936
rect 9484 4976 9524 4985
rect 9388 4842 9428 4927
rect 9484 4145 9524 4936
rect 9579 4976 9621 4985
rect 9579 4936 9580 4976
rect 9620 4936 9621 4976
rect 9579 4927 9621 4936
rect 9292 4136 9332 4145
rect 5876 4096 6068 4136
rect 9196 4096 9292 4136
rect 5836 4087 5876 4096
rect 4108 3968 4148 3977
rect 3628 3928 4108 3968
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 2860 2708 2900 2717
rect 2764 2668 2860 2708
rect 2860 2659 2900 2668
rect 3628 2624 3668 3928
rect 4108 3919 4148 3928
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 4108 3296 4148 3305
rect 3628 2575 3668 2584
rect 4012 3256 4108 3296
rect 4012 2624 4052 3256
rect 4108 3247 4148 3256
rect 6028 2876 6068 4096
rect 9292 4087 9332 4096
rect 9483 4136 9525 4145
rect 9483 4096 9484 4136
rect 9524 4096 9525 4136
rect 9483 4087 9525 4096
rect 9580 4136 9620 4927
rect 9580 4087 9620 4096
rect 9484 4002 9524 4087
rect 9388 3968 9428 3977
rect 9196 3928 9388 3968
rect 9196 3548 9236 3928
rect 9388 3919 9428 3928
rect 9196 3499 9236 3508
rect 9580 3464 9620 3473
rect 10444 3464 10484 7180
rect 11692 7160 11732 7699
rect 11692 7111 11732 7120
rect 11980 7001 12020 7960
rect 12076 7951 12116 7960
rect 12268 7832 12308 7841
rect 12268 7220 12308 7792
rect 12076 7180 12308 7220
rect 12076 7160 12116 7180
rect 12076 7111 12116 7120
rect 12940 7160 12980 8623
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 12940 7111 12980 7120
rect 11979 6992 12021 7001
rect 11979 6952 11980 6992
rect 12020 6952 12021 6992
rect 11979 6943 12021 6952
rect 14091 6992 14133 7001
rect 14091 6952 14092 6992
rect 14132 6952 14133 6992
rect 14091 6943 14133 6952
rect 11980 6413 12020 6943
rect 14092 6858 14132 6943
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 11979 6404 12021 6413
rect 11979 6364 11980 6404
rect 12020 6364 12021 6404
rect 11979 6355 12021 6364
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 11307 4304 11349 4313
rect 11307 4264 11308 4304
rect 11348 4264 11349 4304
rect 11307 4255 11349 4264
rect 11595 4304 11637 4313
rect 11595 4264 11596 4304
rect 11636 4264 11637 4304
rect 11595 4255 11637 4264
rect 10635 4136 10677 4145
rect 10635 4096 10636 4136
rect 10676 4096 10677 4136
rect 10635 4087 10677 4096
rect 11308 4136 11348 4255
rect 11308 4087 11348 4096
rect 10636 4002 10676 4087
rect 11596 3632 11636 4255
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 11596 3583 11636 3592
rect 9620 3424 9716 3464
rect 9580 3415 9620 3424
rect 6028 2827 6068 2836
rect 9676 2792 9716 3424
rect 9676 2743 9716 2752
rect 10444 2633 10484 3424
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 4012 2575 4052 2584
rect 4875 2624 4917 2633
rect 4875 2584 4876 2624
rect 4916 2584 4917 2624
rect 4875 2575 4917 2584
rect 10443 2624 10485 2633
rect 10443 2584 10444 2624
rect 10484 2584 10485 2624
rect 10443 2575 10485 2584
rect 4876 2490 4916 2575
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 844 37948 884 37988
rect 2188 37948 2228 37988
rect 652 37528 692 37568
rect 556 22408 596 22448
rect 652 21568 692 21608
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 9868 36688 9908 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3532 21652 3572 21692
rect 4972 21652 5012 21692
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 2188 20896 2228 20936
rect 2764 20896 2804 20936
rect 3724 20896 3764 20936
rect 6220 21568 6260 21608
rect 8908 21568 8948 21608
rect 6220 21316 6260 21356
rect 7372 21316 7412 21356
rect 2668 20812 2708 20852
rect 652 20728 692 20768
rect 844 20728 884 20768
rect 2380 20728 2420 20768
rect 2572 20728 2612 20768
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 652 15688 692 15728
rect 844 15184 884 15224
rect 652 14848 692 14888
rect 844 14764 884 14804
rect 2188 14764 2228 14804
rect 652 14008 692 14048
rect 844 13252 884 13292
rect 652 13168 692 13208
rect 844 12412 884 12452
rect 2092 12412 2132 12452
rect 652 12328 692 12368
rect 652 11488 692 11528
rect 844 10900 884 10940
rect 652 10732 692 10772
rect 844 10228 884 10268
rect 652 9808 692 9848
rect 844 9388 884 9428
rect 652 8968 692 9008
rect 748 8800 788 8840
rect 652 8128 692 8168
rect 652 7288 692 7328
rect 844 8716 884 8756
rect 940 8632 980 8672
rect 940 7708 980 7748
rect 652 6448 692 6488
rect 844 6196 884 6236
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 844 4768 884 4808
rect 844 4264 884 4304
rect 652 3928 692 3968
rect 1132 10900 1172 10940
rect 1036 4852 1076 4892
rect 2188 12160 2228 12200
rect 2284 11740 2324 11780
rect 2860 20728 2900 20768
rect 3244 20728 3284 20768
rect 3532 20728 3572 20768
rect 3436 20644 3476 20684
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 5548 20728 5588 20768
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3724 16108 3764 16148
rect 4108 16108 4148 16148
rect 2860 15184 2900 15224
rect 2476 13252 2516 13292
rect 2764 13168 2804 13208
rect 2476 11908 2516 11948
rect 2380 11488 2420 11528
rect 2284 9388 2324 9428
rect 2188 8884 2228 8924
rect 2284 8800 2324 8840
rect 2572 11824 2612 11864
rect 2572 11656 2612 11696
rect 2764 10228 2804 10268
rect 2668 8716 2708 8756
rect 2572 8632 2612 8672
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 3916 14008 3956 14048
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4012 13336 4052 13376
rect 3628 13168 3668 13208
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 4780 13336 4820 13376
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3436 11824 3476 11864
rect 3052 11740 3092 11780
rect 2956 11656 2996 11696
rect 3244 11656 3284 11696
rect 2956 11488 2996 11528
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 8428 16444 8468 16484
rect 8812 16444 8852 16484
rect 8620 16192 8660 16232
rect 8428 16024 8468 16064
rect 9004 16108 9044 16148
rect 8908 16024 8948 16064
rect 9196 16192 9236 16232
rect 8908 11908 8948 11948
rect 6220 11740 6260 11780
rect 8524 11740 8564 11780
rect 4396 11656 4436 11696
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8812 11656 8852 11696
rect 9580 14680 9620 14720
rect 9580 14008 9620 14048
rect 9676 12916 9716 12956
rect 9100 11740 9140 11780
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 10252 16108 10292 16148
rect 10060 15184 10100 15224
rect 10156 13168 10196 13208
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 10444 14008 10484 14048
rect 10348 12916 10388 12956
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 14380 14680 14420 14720
rect 11308 14176 11348 14216
rect 13132 14176 13172 14216
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 11212 14008 11252 14048
rect 13516 14008 13556 14048
rect 14188 14008 14228 14048
rect 15532 14008 15572 14048
rect 11404 13168 11444 13208
rect 11116 12916 11156 12956
rect 9772 11908 9812 11948
rect 9004 11656 9044 11696
rect 9196 11572 9236 11612
rect 8716 10984 8756 11024
rect 4204 9976 4244 10016
rect 4780 9976 4820 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 4108 9472 4148 9512
rect 4780 9472 4820 9512
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 2860 8884 2900 8924
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 2668 7708 2708 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 2092 6364 2132 6404
rect 2668 6196 2708 6236
rect 2668 4768 2708 4808
rect 1132 4348 1172 4388
rect 2668 4264 2708 4304
rect 652 3172 692 3212
rect 844 2752 884 2792
rect 2668 2752 2708 2792
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 5356 8800 5396 8840
rect 7180 8800 7220 8840
rect 7372 8800 7412 8840
rect 4972 7372 5012 7412
rect 4780 6448 4820 6488
rect 2860 6364 2900 6404
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4012 5104 4052 5144
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3820 4936 3860 4976
rect 2860 4852 2900 4892
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4972 5104 5012 5144
rect 5644 8632 5684 8672
rect 7084 8632 7124 8672
rect 8716 8632 8756 8672
rect 5548 7372 5588 7412
rect 5260 4936 5300 4976
rect 4108 4432 4148 4472
rect 2860 4348 2900 4388
rect 3916 4348 3956 4388
rect 5164 4432 5204 4472
rect 7084 8044 7124 8084
rect 8428 8044 8468 8084
rect 8524 7960 8564 8000
rect 8812 7960 8852 8000
rect 8428 7876 8468 7916
rect 9964 11824 10004 11864
rect 10828 11824 10868 11864
rect 9868 11740 9908 11780
rect 9964 11656 10004 11696
rect 9772 11152 9812 11192
rect 9292 10984 9332 11024
rect 9676 9976 9716 10016
rect 9292 8800 9332 8840
rect 9196 8128 9236 8168
rect 14092 12160 14132 12200
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 14188 11908 14228 11948
rect 13420 11656 13460 11696
rect 14092 11656 14132 11696
rect 16492 11656 16532 11696
rect 12748 11572 12788 11612
rect 13996 11572 14036 11612
rect 12076 11152 12116 11192
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 12460 9640 12500 9680
rect 12940 9640 12980 9680
rect 15340 9640 15380 9680
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 9676 8632 9716 8672
rect 10540 8632 10580 8672
rect 12940 8632 12980 8672
rect 10444 8128 10484 8168
rect 9004 7372 9044 7412
rect 11404 7876 11444 7916
rect 11116 7708 11156 7748
rect 11692 7708 11732 7748
rect 9292 6448 9332 6488
rect 9100 4936 9140 4976
rect 5836 4852 5876 4892
rect 5548 4432 5588 4472
rect 5356 4264 5396 4304
rect 9388 4936 9428 4976
rect 9580 4936 9620 4976
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 9484 4096 9524 4136
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 11980 6952 12020 6992
rect 14092 6952 14132 6992
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 11980 6364 12020 6404
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 11308 4264 11348 4304
rect 11596 4264 11636 4304
rect 10636 4096 10676 4136
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4876 2584 4916 2624
rect 10444 2584 10484 2624
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 95063 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 95449 38576
rect 835 37948 844 37988
rect 884 37948 2188 37988
rect 2228 37948 2237 37988
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 93823 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 94209 37820
rect 0 37568 80 37588
rect 0 37528 652 37568
rect 692 37528 701 37568
rect 0 37508 80 37528
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 95063 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 95449 37064
rect 0 36728 80 36748
rect 0 36688 9868 36728
rect 9908 36688 9917 36728
rect 0 36668 80 36688
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 93823 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 94209 36308
rect 0 35828 80 35908
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 95063 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 95449 35552
rect 0 34988 80 35068
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 93823 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 94209 34796
rect 0 34148 80 34228
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 95063 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 95449 34040
rect 0 33308 80 33388
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 93823 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 94209 33284
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 95063 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 95449 32528
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 93823 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 94209 31772
rect 0 31628 80 31708
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 95063 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 95449 31016
rect 0 30788 80 30868
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 93823 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 94209 30260
rect 0 29948 80 30028
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 95063 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 95449 29504
rect 0 29108 80 29188
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 93823 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 94209 28748
rect 0 28268 80 28348
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 95063 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 95449 27992
rect 0 27428 80 27508
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 93823 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 94209 27236
rect 0 26588 80 26668
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 95063 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 95449 26480
rect 0 25748 80 25828
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 93823 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 94209 25724
rect 0 24908 80 24988
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 95063 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 95449 24968
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 93823 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 94209 24212
rect 0 24068 80 24148
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 95063 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 95449 23456
rect 0 23228 80 23308
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 93823 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 94209 22700
rect 0 22448 80 22468
rect 0 22408 556 22448
rect 596 22408 605 22448
rect 0 22388 80 22408
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 3523 21652 3532 21692
rect 3572 21652 4972 21692
rect 5012 21652 5021 21692
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 6211 21568 6220 21608
rect 6260 21568 8908 21608
rect 8948 21568 8957 21608
rect 0 21548 80 21568
rect 6211 21316 6220 21356
rect 6260 21316 7372 21356
rect 7412 21316 7421 21356
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 2179 20896 2188 20936
rect 2228 20896 2764 20936
rect 2804 20896 3724 20936
rect 3764 20896 3773 20936
rect 2659 20812 2668 20852
rect 2708 20812 3572 20852
rect 0 20768 80 20788
rect 3532 20768 3572 20812
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 835 20728 844 20768
rect 884 20728 2380 20768
rect 2420 20728 2572 20768
rect 2612 20728 2621 20768
rect 2851 20728 2860 20768
rect 2900 20728 3244 20768
rect 3284 20728 3293 20768
rect 3523 20728 3532 20768
rect 3572 20728 5548 20768
rect 5588 20728 5597 20768
rect 0 20708 80 20728
rect 2572 20684 2612 20728
rect 2572 20644 3436 20684
rect 3476 20644 3485 20684
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 0 19868 80 19888
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 0 19028 80 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 95063 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 95449 18920
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 93823 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 94209 18164
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 95063 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 95449 17408
rect 0 17348 80 17368
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 93823 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 94209 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 0 16508 80 16528
rect 8419 16444 8428 16484
rect 8468 16444 8812 16484
rect 8852 16444 8861 16484
rect 8611 16192 8620 16232
rect 8660 16192 9196 16232
rect 9236 16192 9245 16232
rect 3715 16108 3724 16148
rect 3764 16108 4108 16148
rect 4148 16108 9004 16148
rect 9044 16108 10252 16148
rect 10292 16108 10301 16148
rect 8419 16024 8428 16064
rect 8468 16024 8908 16064
rect 8948 16024 8957 16064
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 95063 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 95449 15896
rect 0 15728 80 15748
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 0 15668 80 15688
rect 835 15184 844 15224
rect 884 15184 2860 15224
rect 2900 15184 10060 15224
rect 10100 15184 10109 15224
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 93823 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 94209 15140
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 0 14828 80 14848
rect 835 14764 844 14804
rect 884 14764 2188 14804
rect 2228 14764 2237 14804
rect 9571 14680 9580 14720
rect 9620 14680 14380 14720
rect 14420 14680 14429 14720
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 95063 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 95449 14384
rect 11299 14176 11308 14216
rect 11348 14176 13132 14216
rect 13172 14176 13181 14216
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 3907 14008 3916 14048
rect 3956 14008 9580 14048
rect 9620 14008 9629 14048
rect 10435 14008 10444 14048
rect 10484 14008 11212 14048
rect 11252 14008 13516 14048
rect 13556 14008 13565 14048
rect 14179 14008 14188 14048
rect 14228 14008 15532 14048
rect 15572 14008 15581 14048
rect 0 13988 80 14008
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 93823 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 94209 13628
rect 4003 13336 4012 13376
rect 4052 13336 4780 13376
rect 4820 13336 4829 13376
rect 835 13252 844 13292
rect 884 13252 2476 13292
rect 2516 13252 2525 13292
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 2755 13168 2764 13208
rect 2804 13168 3628 13208
rect 3668 13168 3677 13208
rect 10147 13168 10156 13208
rect 10196 13168 11404 13208
rect 11444 13168 11453 13208
rect 0 13148 80 13168
rect 9667 12916 9676 12956
rect 9716 12916 10348 12956
rect 10388 12916 11116 12956
rect 11156 12916 11165 12956
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 95063 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 95449 12872
rect 835 12412 844 12452
rect 884 12412 2092 12452
rect 2132 12412 2141 12452
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 0 12308 80 12328
rect 2179 12160 2188 12200
rect 2228 12160 14092 12200
rect 14132 12160 14141 12200
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 93823 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 94209 12116
rect 2467 11908 2476 11948
rect 2516 11908 8908 11948
rect 8948 11908 9772 11948
rect 9812 11908 14188 11948
rect 14228 11908 14237 11948
rect 2563 11824 2572 11864
rect 2612 11824 3436 11864
rect 3476 11824 3485 11864
rect 9955 11824 9964 11864
rect 10004 11824 10828 11864
rect 10868 11824 10877 11864
rect 2275 11740 2284 11780
rect 2324 11740 3052 11780
rect 3092 11740 6220 11780
rect 6260 11740 6269 11780
rect 8515 11740 8524 11780
rect 8564 11740 9100 11780
rect 9140 11740 9868 11780
rect 9908 11740 9917 11780
rect 2563 11656 2572 11696
rect 2612 11656 2956 11696
rect 2996 11656 3005 11696
rect 3235 11656 3244 11696
rect 3284 11656 4396 11696
rect 4436 11656 8812 11696
rect 8852 11656 8861 11696
rect 8995 11656 9004 11696
rect 9044 11656 9964 11696
rect 10004 11656 13420 11696
rect 13460 11656 13469 11696
rect 14083 11656 14092 11696
rect 14132 11656 16492 11696
rect 16532 11656 16541 11696
rect 8812 11612 8852 11656
rect 8812 11572 9196 11612
rect 9236 11572 9245 11612
rect 12739 11572 12748 11612
rect 12788 11572 13996 11612
rect 14036 11572 14045 11612
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 2371 11488 2380 11528
rect 2420 11488 2956 11528
rect 2996 11488 3005 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 95063 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 95449 11360
rect 9763 11152 9772 11192
rect 9812 11152 12076 11192
rect 12116 11152 12125 11192
rect 8707 10984 8716 11024
rect 8756 10984 9292 11024
rect 9332 10984 9341 11024
rect 835 10900 844 10940
rect 884 10900 1132 10940
rect 1172 10900 1181 10940
rect 643 10732 652 10772
rect 692 10732 701 10772
rect 0 10688 80 10708
rect 652 10688 692 10732
rect 0 10648 692 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 93823 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 94209 10604
rect 835 10228 844 10268
rect 884 10228 2764 10268
rect 2804 10228 2813 10268
rect 4195 9976 4204 10016
rect 4244 9976 4780 10016
rect 4820 9976 9676 10016
rect 9716 9976 9725 10016
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 95063 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 95449 9848
rect 0 9788 80 9808
rect 12451 9640 12460 9680
rect 12500 9640 12940 9680
rect 12980 9640 15340 9680
rect 15380 9640 15389 9680
rect 4099 9472 4108 9512
rect 4148 9472 4780 9512
rect 4820 9472 4829 9512
rect 835 9388 844 9428
rect 884 9388 2284 9428
rect 2324 9388 2333 9428
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 2179 8884 2188 8924
rect 2228 8884 2860 8924
rect 2900 8884 2909 8924
rect 739 8800 748 8840
rect 788 8800 2284 8840
rect 2324 8800 2333 8840
rect 5347 8800 5356 8840
rect 5396 8800 7180 8840
rect 7220 8800 7229 8840
rect 7363 8800 7372 8840
rect 7412 8800 9292 8840
rect 9332 8800 9341 8840
rect 835 8716 844 8756
rect 884 8716 2668 8756
rect 2708 8716 2717 8756
rect 931 8632 940 8672
rect 980 8632 2572 8672
rect 2612 8632 2621 8672
rect 5635 8632 5644 8672
rect 5684 8632 7084 8672
rect 7124 8632 7133 8672
rect 8707 8632 8716 8672
rect 8756 8632 9676 8672
rect 9716 8632 9725 8672
rect 10531 8632 10540 8672
rect 10580 8632 12940 8672
rect 12980 8632 12989 8672
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 9187 8128 9196 8168
rect 9236 8128 10444 8168
rect 10484 8128 10493 8168
rect 0 8108 80 8128
rect 7075 8044 7084 8084
rect 7124 8044 8428 8084
rect 8468 8044 8477 8084
rect 8515 7960 8524 8000
rect 8564 7960 8812 8000
rect 8852 7960 8861 8000
rect 8419 7876 8428 7916
rect 8468 7876 11404 7916
rect 11444 7876 11453 7916
rect 931 7708 940 7748
rect 980 7708 2668 7748
rect 2708 7708 2717 7748
rect 11107 7708 11116 7748
rect 11156 7708 11692 7748
rect 11732 7708 11741 7748
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 4963 7372 4972 7412
rect 5012 7372 5548 7412
rect 5588 7372 9004 7412
rect 9044 7372 9053 7412
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 0 7268 80 7288
rect 11971 6952 11980 6992
rect 12020 6952 14092 6992
rect 14132 6952 14141 6992
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 4771 6448 4780 6488
rect 4820 6448 9292 6488
rect 9332 6448 9341 6488
rect 0 6428 80 6448
rect 2083 6364 2092 6404
rect 2132 6364 2860 6404
rect 2900 6364 11980 6404
rect 12020 6364 12029 6404
rect 835 6196 844 6236
rect 884 6196 2668 6236
rect 2708 6196 2717 6236
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 0 5588 80 5608
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 4003 5104 4012 5144
rect 4052 5104 4972 5144
rect 5012 5104 5021 5144
rect 3811 4936 3820 4976
rect 3860 4936 5260 4976
rect 5300 4936 9100 4976
rect 9140 4936 9388 4976
rect 9428 4936 9580 4976
rect 9620 4936 9629 4976
rect 1027 4852 1036 4892
rect 1076 4852 2860 4892
rect 2900 4852 5836 4892
rect 5876 4852 5885 4892
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 835 4768 844 4808
rect 884 4768 2668 4808
rect 2708 4768 2717 4808
rect 0 4748 80 4768
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 4099 4432 4108 4472
rect 4148 4432 5164 4472
rect 5204 4432 5548 4472
rect 5588 4432 5597 4472
rect 1123 4348 1132 4388
rect 1172 4348 2860 4388
rect 2900 4348 3916 4388
rect 3956 4348 4340 4388
rect 4300 4304 4340 4348
rect 835 4264 844 4304
rect 884 4264 2668 4304
rect 2708 4264 2717 4304
rect 4300 4264 5356 4304
rect 5396 4264 11308 4304
rect 11348 4264 11596 4304
rect 11636 4264 11645 4304
rect 9475 4096 9484 4136
rect 9524 4096 10636 4136
rect 10676 4096 10685 4136
rect 0 3968 80 3988
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 0 3908 80 3928
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 835 2752 844 2792
rect 884 2752 2668 2792
rect 2708 2752 2717 2792
rect 4867 2584 4876 2624
rect 4916 2584 10444 2624
rect 10484 2584 10493 2624
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 0 2228 80 2248
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal5 >>
rect 4343 38576 4390 38618
rect 4514 38576 4558 38618
rect 4682 38576 4729 38618
rect 4343 38536 4352 38576
rect 4514 38536 4516 38576
rect 4556 38536 4558 38576
rect 4720 38536 4729 38576
rect 4343 38494 4390 38536
rect 4514 38494 4558 38536
rect 4682 38494 4729 38536
rect 19463 38576 19510 38618
rect 19634 38576 19678 38618
rect 19802 38576 19849 38618
rect 19463 38536 19472 38576
rect 19634 38536 19636 38576
rect 19676 38536 19678 38576
rect 19840 38536 19849 38576
rect 19463 38494 19510 38536
rect 19634 38494 19678 38536
rect 19802 38494 19849 38536
rect 34583 38576 34630 38618
rect 34754 38576 34798 38618
rect 34922 38576 34969 38618
rect 34583 38536 34592 38576
rect 34754 38536 34756 38576
rect 34796 38536 34798 38576
rect 34960 38536 34969 38576
rect 34583 38494 34630 38536
rect 34754 38494 34798 38536
rect 34922 38494 34969 38536
rect 49703 38576 49750 38618
rect 49874 38576 49918 38618
rect 50042 38576 50089 38618
rect 49703 38536 49712 38576
rect 49874 38536 49876 38576
rect 49916 38536 49918 38576
rect 50080 38536 50089 38576
rect 49703 38494 49750 38536
rect 49874 38494 49918 38536
rect 50042 38494 50089 38536
rect 64823 38576 64870 38618
rect 64994 38576 65038 38618
rect 65162 38576 65209 38618
rect 64823 38536 64832 38576
rect 64994 38536 64996 38576
rect 65036 38536 65038 38576
rect 65200 38536 65209 38576
rect 64823 38494 64870 38536
rect 64994 38494 65038 38536
rect 65162 38494 65209 38536
rect 79943 38576 79990 38618
rect 80114 38576 80158 38618
rect 80282 38576 80329 38618
rect 79943 38536 79952 38576
rect 80114 38536 80116 38576
rect 80156 38536 80158 38576
rect 80320 38536 80329 38576
rect 79943 38494 79990 38536
rect 80114 38494 80158 38536
rect 80282 38494 80329 38536
rect 95063 38576 95110 38618
rect 95234 38576 95278 38618
rect 95402 38576 95449 38618
rect 95063 38536 95072 38576
rect 95234 38536 95236 38576
rect 95276 38536 95278 38576
rect 95440 38536 95449 38576
rect 95063 38494 95110 38536
rect 95234 38494 95278 38536
rect 95402 38494 95449 38536
rect 3103 37820 3150 37862
rect 3274 37820 3318 37862
rect 3442 37820 3489 37862
rect 3103 37780 3112 37820
rect 3274 37780 3276 37820
rect 3316 37780 3318 37820
rect 3480 37780 3489 37820
rect 3103 37738 3150 37780
rect 3274 37738 3318 37780
rect 3442 37738 3489 37780
rect 18223 37820 18270 37862
rect 18394 37820 18438 37862
rect 18562 37820 18609 37862
rect 18223 37780 18232 37820
rect 18394 37780 18396 37820
rect 18436 37780 18438 37820
rect 18600 37780 18609 37820
rect 18223 37738 18270 37780
rect 18394 37738 18438 37780
rect 18562 37738 18609 37780
rect 33343 37820 33390 37862
rect 33514 37820 33558 37862
rect 33682 37820 33729 37862
rect 33343 37780 33352 37820
rect 33514 37780 33516 37820
rect 33556 37780 33558 37820
rect 33720 37780 33729 37820
rect 33343 37738 33390 37780
rect 33514 37738 33558 37780
rect 33682 37738 33729 37780
rect 48463 37820 48510 37862
rect 48634 37820 48678 37862
rect 48802 37820 48849 37862
rect 48463 37780 48472 37820
rect 48634 37780 48636 37820
rect 48676 37780 48678 37820
rect 48840 37780 48849 37820
rect 48463 37738 48510 37780
rect 48634 37738 48678 37780
rect 48802 37738 48849 37780
rect 63583 37820 63630 37862
rect 63754 37820 63798 37862
rect 63922 37820 63969 37862
rect 63583 37780 63592 37820
rect 63754 37780 63756 37820
rect 63796 37780 63798 37820
rect 63960 37780 63969 37820
rect 63583 37738 63630 37780
rect 63754 37738 63798 37780
rect 63922 37738 63969 37780
rect 78703 37820 78750 37862
rect 78874 37820 78918 37862
rect 79042 37820 79089 37862
rect 78703 37780 78712 37820
rect 78874 37780 78876 37820
rect 78916 37780 78918 37820
rect 79080 37780 79089 37820
rect 78703 37738 78750 37780
rect 78874 37738 78918 37780
rect 79042 37738 79089 37780
rect 93823 37820 93870 37862
rect 93994 37820 94038 37862
rect 94162 37820 94209 37862
rect 93823 37780 93832 37820
rect 93994 37780 93996 37820
rect 94036 37780 94038 37820
rect 94200 37780 94209 37820
rect 93823 37738 93870 37780
rect 93994 37738 94038 37780
rect 94162 37738 94209 37780
rect 4343 37064 4390 37106
rect 4514 37064 4558 37106
rect 4682 37064 4729 37106
rect 4343 37024 4352 37064
rect 4514 37024 4516 37064
rect 4556 37024 4558 37064
rect 4720 37024 4729 37064
rect 4343 36982 4390 37024
rect 4514 36982 4558 37024
rect 4682 36982 4729 37024
rect 19463 37064 19510 37106
rect 19634 37064 19678 37106
rect 19802 37064 19849 37106
rect 19463 37024 19472 37064
rect 19634 37024 19636 37064
rect 19676 37024 19678 37064
rect 19840 37024 19849 37064
rect 19463 36982 19510 37024
rect 19634 36982 19678 37024
rect 19802 36982 19849 37024
rect 34583 37064 34630 37106
rect 34754 37064 34798 37106
rect 34922 37064 34969 37106
rect 34583 37024 34592 37064
rect 34754 37024 34756 37064
rect 34796 37024 34798 37064
rect 34960 37024 34969 37064
rect 34583 36982 34630 37024
rect 34754 36982 34798 37024
rect 34922 36982 34969 37024
rect 49703 37064 49750 37106
rect 49874 37064 49918 37106
rect 50042 37064 50089 37106
rect 49703 37024 49712 37064
rect 49874 37024 49876 37064
rect 49916 37024 49918 37064
rect 50080 37024 50089 37064
rect 49703 36982 49750 37024
rect 49874 36982 49918 37024
rect 50042 36982 50089 37024
rect 64823 37064 64870 37106
rect 64994 37064 65038 37106
rect 65162 37064 65209 37106
rect 64823 37024 64832 37064
rect 64994 37024 64996 37064
rect 65036 37024 65038 37064
rect 65200 37024 65209 37064
rect 64823 36982 64870 37024
rect 64994 36982 65038 37024
rect 65162 36982 65209 37024
rect 79943 37064 79990 37106
rect 80114 37064 80158 37106
rect 80282 37064 80329 37106
rect 79943 37024 79952 37064
rect 80114 37024 80116 37064
rect 80156 37024 80158 37064
rect 80320 37024 80329 37064
rect 79943 36982 79990 37024
rect 80114 36982 80158 37024
rect 80282 36982 80329 37024
rect 95063 37064 95110 37106
rect 95234 37064 95278 37106
rect 95402 37064 95449 37106
rect 95063 37024 95072 37064
rect 95234 37024 95236 37064
rect 95276 37024 95278 37064
rect 95440 37024 95449 37064
rect 95063 36982 95110 37024
rect 95234 36982 95278 37024
rect 95402 36982 95449 37024
rect 3103 36308 3150 36350
rect 3274 36308 3318 36350
rect 3442 36308 3489 36350
rect 3103 36268 3112 36308
rect 3274 36268 3276 36308
rect 3316 36268 3318 36308
rect 3480 36268 3489 36308
rect 3103 36226 3150 36268
rect 3274 36226 3318 36268
rect 3442 36226 3489 36268
rect 18223 36308 18270 36350
rect 18394 36308 18438 36350
rect 18562 36308 18609 36350
rect 18223 36268 18232 36308
rect 18394 36268 18396 36308
rect 18436 36268 18438 36308
rect 18600 36268 18609 36308
rect 18223 36226 18270 36268
rect 18394 36226 18438 36268
rect 18562 36226 18609 36268
rect 33343 36308 33390 36350
rect 33514 36308 33558 36350
rect 33682 36308 33729 36350
rect 33343 36268 33352 36308
rect 33514 36268 33516 36308
rect 33556 36268 33558 36308
rect 33720 36268 33729 36308
rect 33343 36226 33390 36268
rect 33514 36226 33558 36268
rect 33682 36226 33729 36268
rect 48463 36308 48510 36350
rect 48634 36308 48678 36350
rect 48802 36308 48849 36350
rect 48463 36268 48472 36308
rect 48634 36268 48636 36308
rect 48676 36268 48678 36308
rect 48840 36268 48849 36308
rect 48463 36226 48510 36268
rect 48634 36226 48678 36268
rect 48802 36226 48849 36268
rect 63583 36308 63630 36350
rect 63754 36308 63798 36350
rect 63922 36308 63969 36350
rect 63583 36268 63592 36308
rect 63754 36268 63756 36308
rect 63796 36268 63798 36308
rect 63960 36268 63969 36308
rect 63583 36226 63630 36268
rect 63754 36226 63798 36268
rect 63922 36226 63969 36268
rect 78703 36308 78750 36350
rect 78874 36308 78918 36350
rect 79042 36308 79089 36350
rect 78703 36268 78712 36308
rect 78874 36268 78876 36308
rect 78916 36268 78918 36308
rect 79080 36268 79089 36308
rect 78703 36226 78750 36268
rect 78874 36226 78918 36268
rect 79042 36226 79089 36268
rect 93823 36308 93870 36350
rect 93994 36308 94038 36350
rect 94162 36308 94209 36350
rect 93823 36268 93832 36308
rect 93994 36268 93996 36308
rect 94036 36268 94038 36308
rect 94200 36268 94209 36308
rect 93823 36226 93870 36268
rect 93994 36226 94038 36268
rect 94162 36226 94209 36268
rect 4343 35552 4390 35594
rect 4514 35552 4558 35594
rect 4682 35552 4729 35594
rect 4343 35512 4352 35552
rect 4514 35512 4516 35552
rect 4556 35512 4558 35552
rect 4720 35512 4729 35552
rect 4343 35470 4390 35512
rect 4514 35470 4558 35512
rect 4682 35470 4729 35512
rect 19463 35552 19510 35594
rect 19634 35552 19678 35594
rect 19802 35552 19849 35594
rect 19463 35512 19472 35552
rect 19634 35512 19636 35552
rect 19676 35512 19678 35552
rect 19840 35512 19849 35552
rect 19463 35470 19510 35512
rect 19634 35470 19678 35512
rect 19802 35470 19849 35512
rect 34583 35552 34630 35594
rect 34754 35552 34798 35594
rect 34922 35552 34969 35594
rect 34583 35512 34592 35552
rect 34754 35512 34756 35552
rect 34796 35512 34798 35552
rect 34960 35512 34969 35552
rect 34583 35470 34630 35512
rect 34754 35470 34798 35512
rect 34922 35470 34969 35512
rect 49703 35552 49750 35594
rect 49874 35552 49918 35594
rect 50042 35552 50089 35594
rect 49703 35512 49712 35552
rect 49874 35512 49876 35552
rect 49916 35512 49918 35552
rect 50080 35512 50089 35552
rect 49703 35470 49750 35512
rect 49874 35470 49918 35512
rect 50042 35470 50089 35512
rect 64823 35552 64870 35594
rect 64994 35552 65038 35594
rect 65162 35552 65209 35594
rect 64823 35512 64832 35552
rect 64994 35512 64996 35552
rect 65036 35512 65038 35552
rect 65200 35512 65209 35552
rect 64823 35470 64870 35512
rect 64994 35470 65038 35512
rect 65162 35470 65209 35512
rect 79943 35552 79990 35594
rect 80114 35552 80158 35594
rect 80282 35552 80329 35594
rect 79943 35512 79952 35552
rect 80114 35512 80116 35552
rect 80156 35512 80158 35552
rect 80320 35512 80329 35552
rect 79943 35470 79990 35512
rect 80114 35470 80158 35512
rect 80282 35470 80329 35512
rect 95063 35552 95110 35594
rect 95234 35552 95278 35594
rect 95402 35552 95449 35594
rect 95063 35512 95072 35552
rect 95234 35512 95236 35552
rect 95276 35512 95278 35552
rect 95440 35512 95449 35552
rect 95063 35470 95110 35512
rect 95234 35470 95278 35512
rect 95402 35470 95449 35512
rect 3103 34796 3150 34838
rect 3274 34796 3318 34838
rect 3442 34796 3489 34838
rect 3103 34756 3112 34796
rect 3274 34756 3276 34796
rect 3316 34756 3318 34796
rect 3480 34756 3489 34796
rect 3103 34714 3150 34756
rect 3274 34714 3318 34756
rect 3442 34714 3489 34756
rect 18223 34796 18270 34838
rect 18394 34796 18438 34838
rect 18562 34796 18609 34838
rect 18223 34756 18232 34796
rect 18394 34756 18396 34796
rect 18436 34756 18438 34796
rect 18600 34756 18609 34796
rect 18223 34714 18270 34756
rect 18394 34714 18438 34756
rect 18562 34714 18609 34756
rect 33343 34796 33390 34838
rect 33514 34796 33558 34838
rect 33682 34796 33729 34838
rect 33343 34756 33352 34796
rect 33514 34756 33516 34796
rect 33556 34756 33558 34796
rect 33720 34756 33729 34796
rect 33343 34714 33390 34756
rect 33514 34714 33558 34756
rect 33682 34714 33729 34756
rect 48463 34796 48510 34838
rect 48634 34796 48678 34838
rect 48802 34796 48849 34838
rect 48463 34756 48472 34796
rect 48634 34756 48636 34796
rect 48676 34756 48678 34796
rect 48840 34756 48849 34796
rect 48463 34714 48510 34756
rect 48634 34714 48678 34756
rect 48802 34714 48849 34756
rect 63583 34796 63630 34838
rect 63754 34796 63798 34838
rect 63922 34796 63969 34838
rect 63583 34756 63592 34796
rect 63754 34756 63756 34796
rect 63796 34756 63798 34796
rect 63960 34756 63969 34796
rect 63583 34714 63630 34756
rect 63754 34714 63798 34756
rect 63922 34714 63969 34756
rect 78703 34796 78750 34838
rect 78874 34796 78918 34838
rect 79042 34796 79089 34838
rect 78703 34756 78712 34796
rect 78874 34756 78876 34796
rect 78916 34756 78918 34796
rect 79080 34756 79089 34796
rect 78703 34714 78750 34756
rect 78874 34714 78918 34756
rect 79042 34714 79089 34756
rect 93823 34796 93870 34838
rect 93994 34796 94038 34838
rect 94162 34796 94209 34838
rect 93823 34756 93832 34796
rect 93994 34756 93996 34796
rect 94036 34756 94038 34796
rect 94200 34756 94209 34796
rect 93823 34714 93870 34756
rect 93994 34714 94038 34756
rect 94162 34714 94209 34756
rect 4343 34040 4390 34082
rect 4514 34040 4558 34082
rect 4682 34040 4729 34082
rect 4343 34000 4352 34040
rect 4514 34000 4516 34040
rect 4556 34000 4558 34040
rect 4720 34000 4729 34040
rect 4343 33958 4390 34000
rect 4514 33958 4558 34000
rect 4682 33958 4729 34000
rect 19463 34040 19510 34082
rect 19634 34040 19678 34082
rect 19802 34040 19849 34082
rect 19463 34000 19472 34040
rect 19634 34000 19636 34040
rect 19676 34000 19678 34040
rect 19840 34000 19849 34040
rect 19463 33958 19510 34000
rect 19634 33958 19678 34000
rect 19802 33958 19849 34000
rect 34583 34040 34630 34082
rect 34754 34040 34798 34082
rect 34922 34040 34969 34082
rect 34583 34000 34592 34040
rect 34754 34000 34756 34040
rect 34796 34000 34798 34040
rect 34960 34000 34969 34040
rect 34583 33958 34630 34000
rect 34754 33958 34798 34000
rect 34922 33958 34969 34000
rect 49703 34040 49750 34082
rect 49874 34040 49918 34082
rect 50042 34040 50089 34082
rect 49703 34000 49712 34040
rect 49874 34000 49876 34040
rect 49916 34000 49918 34040
rect 50080 34000 50089 34040
rect 49703 33958 49750 34000
rect 49874 33958 49918 34000
rect 50042 33958 50089 34000
rect 64823 34040 64870 34082
rect 64994 34040 65038 34082
rect 65162 34040 65209 34082
rect 64823 34000 64832 34040
rect 64994 34000 64996 34040
rect 65036 34000 65038 34040
rect 65200 34000 65209 34040
rect 64823 33958 64870 34000
rect 64994 33958 65038 34000
rect 65162 33958 65209 34000
rect 79943 34040 79990 34082
rect 80114 34040 80158 34082
rect 80282 34040 80329 34082
rect 79943 34000 79952 34040
rect 80114 34000 80116 34040
rect 80156 34000 80158 34040
rect 80320 34000 80329 34040
rect 79943 33958 79990 34000
rect 80114 33958 80158 34000
rect 80282 33958 80329 34000
rect 95063 34040 95110 34082
rect 95234 34040 95278 34082
rect 95402 34040 95449 34082
rect 95063 34000 95072 34040
rect 95234 34000 95236 34040
rect 95276 34000 95278 34040
rect 95440 34000 95449 34040
rect 95063 33958 95110 34000
rect 95234 33958 95278 34000
rect 95402 33958 95449 34000
rect 3103 33284 3150 33326
rect 3274 33284 3318 33326
rect 3442 33284 3489 33326
rect 3103 33244 3112 33284
rect 3274 33244 3276 33284
rect 3316 33244 3318 33284
rect 3480 33244 3489 33284
rect 3103 33202 3150 33244
rect 3274 33202 3318 33244
rect 3442 33202 3489 33244
rect 18223 33284 18270 33326
rect 18394 33284 18438 33326
rect 18562 33284 18609 33326
rect 18223 33244 18232 33284
rect 18394 33244 18396 33284
rect 18436 33244 18438 33284
rect 18600 33244 18609 33284
rect 18223 33202 18270 33244
rect 18394 33202 18438 33244
rect 18562 33202 18609 33244
rect 33343 33284 33390 33326
rect 33514 33284 33558 33326
rect 33682 33284 33729 33326
rect 33343 33244 33352 33284
rect 33514 33244 33516 33284
rect 33556 33244 33558 33284
rect 33720 33244 33729 33284
rect 33343 33202 33390 33244
rect 33514 33202 33558 33244
rect 33682 33202 33729 33244
rect 48463 33284 48510 33326
rect 48634 33284 48678 33326
rect 48802 33284 48849 33326
rect 48463 33244 48472 33284
rect 48634 33244 48636 33284
rect 48676 33244 48678 33284
rect 48840 33244 48849 33284
rect 48463 33202 48510 33244
rect 48634 33202 48678 33244
rect 48802 33202 48849 33244
rect 63583 33284 63630 33326
rect 63754 33284 63798 33326
rect 63922 33284 63969 33326
rect 63583 33244 63592 33284
rect 63754 33244 63756 33284
rect 63796 33244 63798 33284
rect 63960 33244 63969 33284
rect 63583 33202 63630 33244
rect 63754 33202 63798 33244
rect 63922 33202 63969 33244
rect 78703 33284 78750 33326
rect 78874 33284 78918 33326
rect 79042 33284 79089 33326
rect 78703 33244 78712 33284
rect 78874 33244 78876 33284
rect 78916 33244 78918 33284
rect 79080 33244 79089 33284
rect 78703 33202 78750 33244
rect 78874 33202 78918 33244
rect 79042 33202 79089 33244
rect 93823 33284 93870 33326
rect 93994 33284 94038 33326
rect 94162 33284 94209 33326
rect 93823 33244 93832 33284
rect 93994 33244 93996 33284
rect 94036 33244 94038 33284
rect 94200 33244 94209 33284
rect 93823 33202 93870 33244
rect 93994 33202 94038 33244
rect 94162 33202 94209 33244
rect 4343 32528 4390 32570
rect 4514 32528 4558 32570
rect 4682 32528 4729 32570
rect 4343 32488 4352 32528
rect 4514 32488 4516 32528
rect 4556 32488 4558 32528
rect 4720 32488 4729 32528
rect 4343 32446 4390 32488
rect 4514 32446 4558 32488
rect 4682 32446 4729 32488
rect 19463 32528 19510 32570
rect 19634 32528 19678 32570
rect 19802 32528 19849 32570
rect 19463 32488 19472 32528
rect 19634 32488 19636 32528
rect 19676 32488 19678 32528
rect 19840 32488 19849 32528
rect 19463 32446 19510 32488
rect 19634 32446 19678 32488
rect 19802 32446 19849 32488
rect 34583 32528 34630 32570
rect 34754 32528 34798 32570
rect 34922 32528 34969 32570
rect 34583 32488 34592 32528
rect 34754 32488 34756 32528
rect 34796 32488 34798 32528
rect 34960 32488 34969 32528
rect 34583 32446 34630 32488
rect 34754 32446 34798 32488
rect 34922 32446 34969 32488
rect 49703 32528 49750 32570
rect 49874 32528 49918 32570
rect 50042 32528 50089 32570
rect 49703 32488 49712 32528
rect 49874 32488 49876 32528
rect 49916 32488 49918 32528
rect 50080 32488 50089 32528
rect 49703 32446 49750 32488
rect 49874 32446 49918 32488
rect 50042 32446 50089 32488
rect 64823 32528 64870 32570
rect 64994 32528 65038 32570
rect 65162 32528 65209 32570
rect 64823 32488 64832 32528
rect 64994 32488 64996 32528
rect 65036 32488 65038 32528
rect 65200 32488 65209 32528
rect 64823 32446 64870 32488
rect 64994 32446 65038 32488
rect 65162 32446 65209 32488
rect 79943 32528 79990 32570
rect 80114 32528 80158 32570
rect 80282 32528 80329 32570
rect 79943 32488 79952 32528
rect 80114 32488 80116 32528
rect 80156 32488 80158 32528
rect 80320 32488 80329 32528
rect 79943 32446 79990 32488
rect 80114 32446 80158 32488
rect 80282 32446 80329 32488
rect 95063 32528 95110 32570
rect 95234 32528 95278 32570
rect 95402 32528 95449 32570
rect 95063 32488 95072 32528
rect 95234 32488 95236 32528
rect 95276 32488 95278 32528
rect 95440 32488 95449 32528
rect 95063 32446 95110 32488
rect 95234 32446 95278 32488
rect 95402 32446 95449 32488
rect 3103 31772 3150 31814
rect 3274 31772 3318 31814
rect 3442 31772 3489 31814
rect 3103 31732 3112 31772
rect 3274 31732 3276 31772
rect 3316 31732 3318 31772
rect 3480 31732 3489 31772
rect 3103 31690 3150 31732
rect 3274 31690 3318 31732
rect 3442 31690 3489 31732
rect 18223 31772 18270 31814
rect 18394 31772 18438 31814
rect 18562 31772 18609 31814
rect 18223 31732 18232 31772
rect 18394 31732 18396 31772
rect 18436 31732 18438 31772
rect 18600 31732 18609 31772
rect 18223 31690 18270 31732
rect 18394 31690 18438 31732
rect 18562 31690 18609 31732
rect 33343 31772 33390 31814
rect 33514 31772 33558 31814
rect 33682 31772 33729 31814
rect 33343 31732 33352 31772
rect 33514 31732 33516 31772
rect 33556 31732 33558 31772
rect 33720 31732 33729 31772
rect 33343 31690 33390 31732
rect 33514 31690 33558 31732
rect 33682 31690 33729 31732
rect 48463 31772 48510 31814
rect 48634 31772 48678 31814
rect 48802 31772 48849 31814
rect 48463 31732 48472 31772
rect 48634 31732 48636 31772
rect 48676 31732 48678 31772
rect 48840 31732 48849 31772
rect 48463 31690 48510 31732
rect 48634 31690 48678 31732
rect 48802 31690 48849 31732
rect 63583 31772 63630 31814
rect 63754 31772 63798 31814
rect 63922 31772 63969 31814
rect 63583 31732 63592 31772
rect 63754 31732 63756 31772
rect 63796 31732 63798 31772
rect 63960 31732 63969 31772
rect 63583 31690 63630 31732
rect 63754 31690 63798 31732
rect 63922 31690 63969 31732
rect 78703 31772 78750 31814
rect 78874 31772 78918 31814
rect 79042 31772 79089 31814
rect 78703 31732 78712 31772
rect 78874 31732 78876 31772
rect 78916 31732 78918 31772
rect 79080 31732 79089 31772
rect 78703 31690 78750 31732
rect 78874 31690 78918 31732
rect 79042 31690 79089 31732
rect 93823 31772 93870 31814
rect 93994 31772 94038 31814
rect 94162 31772 94209 31814
rect 93823 31732 93832 31772
rect 93994 31732 93996 31772
rect 94036 31732 94038 31772
rect 94200 31732 94209 31772
rect 93823 31690 93870 31732
rect 93994 31690 94038 31732
rect 94162 31690 94209 31732
rect 4343 31016 4390 31058
rect 4514 31016 4558 31058
rect 4682 31016 4729 31058
rect 4343 30976 4352 31016
rect 4514 30976 4516 31016
rect 4556 30976 4558 31016
rect 4720 30976 4729 31016
rect 4343 30934 4390 30976
rect 4514 30934 4558 30976
rect 4682 30934 4729 30976
rect 19463 31016 19510 31058
rect 19634 31016 19678 31058
rect 19802 31016 19849 31058
rect 19463 30976 19472 31016
rect 19634 30976 19636 31016
rect 19676 30976 19678 31016
rect 19840 30976 19849 31016
rect 19463 30934 19510 30976
rect 19634 30934 19678 30976
rect 19802 30934 19849 30976
rect 34583 31016 34630 31058
rect 34754 31016 34798 31058
rect 34922 31016 34969 31058
rect 34583 30976 34592 31016
rect 34754 30976 34756 31016
rect 34796 30976 34798 31016
rect 34960 30976 34969 31016
rect 34583 30934 34630 30976
rect 34754 30934 34798 30976
rect 34922 30934 34969 30976
rect 49703 31016 49750 31058
rect 49874 31016 49918 31058
rect 50042 31016 50089 31058
rect 49703 30976 49712 31016
rect 49874 30976 49876 31016
rect 49916 30976 49918 31016
rect 50080 30976 50089 31016
rect 49703 30934 49750 30976
rect 49874 30934 49918 30976
rect 50042 30934 50089 30976
rect 64823 31016 64870 31058
rect 64994 31016 65038 31058
rect 65162 31016 65209 31058
rect 64823 30976 64832 31016
rect 64994 30976 64996 31016
rect 65036 30976 65038 31016
rect 65200 30976 65209 31016
rect 64823 30934 64870 30976
rect 64994 30934 65038 30976
rect 65162 30934 65209 30976
rect 79943 31016 79990 31058
rect 80114 31016 80158 31058
rect 80282 31016 80329 31058
rect 79943 30976 79952 31016
rect 80114 30976 80116 31016
rect 80156 30976 80158 31016
rect 80320 30976 80329 31016
rect 79943 30934 79990 30976
rect 80114 30934 80158 30976
rect 80282 30934 80329 30976
rect 95063 31016 95110 31058
rect 95234 31016 95278 31058
rect 95402 31016 95449 31058
rect 95063 30976 95072 31016
rect 95234 30976 95236 31016
rect 95276 30976 95278 31016
rect 95440 30976 95449 31016
rect 95063 30934 95110 30976
rect 95234 30934 95278 30976
rect 95402 30934 95449 30976
rect 3103 30260 3150 30302
rect 3274 30260 3318 30302
rect 3442 30260 3489 30302
rect 3103 30220 3112 30260
rect 3274 30220 3276 30260
rect 3316 30220 3318 30260
rect 3480 30220 3489 30260
rect 3103 30178 3150 30220
rect 3274 30178 3318 30220
rect 3442 30178 3489 30220
rect 18223 30260 18270 30302
rect 18394 30260 18438 30302
rect 18562 30260 18609 30302
rect 18223 30220 18232 30260
rect 18394 30220 18396 30260
rect 18436 30220 18438 30260
rect 18600 30220 18609 30260
rect 18223 30178 18270 30220
rect 18394 30178 18438 30220
rect 18562 30178 18609 30220
rect 33343 30260 33390 30302
rect 33514 30260 33558 30302
rect 33682 30260 33729 30302
rect 33343 30220 33352 30260
rect 33514 30220 33516 30260
rect 33556 30220 33558 30260
rect 33720 30220 33729 30260
rect 33343 30178 33390 30220
rect 33514 30178 33558 30220
rect 33682 30178 33729 30220
rect 48463 30260 48510 30302
rect 48634 30260 48678 30302
rect 48802 30260 48849 30302
rect 48463 30220 48472 30260
rect 48634 30220 48636 30260
rect 48676 30220 48678 30260
rect 48840 30220 48849 30260
rect 48463 30178 48510 30220
rect 48634 30178 48678 30220
rect 48802 30178 48849 30220
rect 63583 30260 63630 30302
rect 63754 30260 63798 30302
rect 63922 30260 63969 30302
rect 63583 30220 63592 30260
rect 63754 30220 63756 30260
rect 63796 30220 63798 30260
rect 63960 30220 63969 30260
rect 63583 30178 63630 30220
rect 63754 30178 63798 30220
rect 63922 30178 63969 30220
rect 78703 30260 78750 30302
rect 78874 30260 78918 30302
rect 79042 30260 79089 30302
rect 78703 30220 78712 30260
rect 78874 30220 78876 30260
rect 78916 30220 78918 30260
rect 79080 30220 79089 30260
rect 78703 30178 78750 30220
rect 78874 30178 78918 30220
rect 79042 30178 79089 30220
rect 93823 30260 93870 30302
rect 93994 30260 94038 30302
rect 94162 30260 94209 30302
rect 93823 30220 93832 30260
rect 93994 30220 93996 30260
rect 94036 30220 94038 30260
rect 94200 30220 94209 30260
rect 93823 30178 93870 30220
rect 93994 30178 94038 30220
rect 94162 30178 94209 30220
rect 4343 29504 4390 29546
rect 4514 29504 4558 29546
rect 4682 29504 4729 29546
rect 4343 29464 4352 29504
rect 4514 29464 4516 29504
rect 4556 29464 4558 29504
rect 4720 29464 4729 29504
rect 4343 29422 4390 29464
rect 4514 29422 4558 29464
rect 4682 29422 4729 29464
rect 19463 29504 19510 29546
rect 19634 29504 19678 29546
rect 19802 29504 19849 29546
rect 19463 29464 19472 29504
rect 19634 29464 19636 29504
rect 19676 29464 19678 29504
rect 19840 29464 19849 29504
rect 19463 29422 19510 29464
rect 19634 29422 19678 29464
rect 19802 29422 19849 29464
rect 34583 29504 34630 29546
rect 34754 29504 34798 29546
rect 34922 29504 34969 29546
rect 34583 29464 34592 29504
rect 34754 29464 34756 29504
rect 34796 29464 34798 29504
rect 34960 29464 34969 29504
rect 34583 29422 34630 29464
rect 34754 29422 34798 29464
rect 34922 29422 34969 29464
rect 49703 29504 49750 29546
rect 49874 29504 49918 29546
rect 50042 29504 50089 29546
rect 49703 29464 49712 29504
rect 49874 29464 49876 29504
rect 49916 29464 49918 29504
rect 50080 29464 50089 29504
rect 49703 29422 49750 29464
rect 49874 29422 49918 29464
rect 50042 29422 50089 29464
rect 64823 29504 64870 29546
rect 64994 29504 65038 29546
rect 65162 29504 65209 29546
rect 64823 29464 64832 29504
rect 64994 29464 64996 29504
rect 65036 29464 65038 29504
rect 65200 29464 65209 29504
rect 64823 29422 64870 29464
rect 64994 29422 65038 29464
rect 65162 29422 65209 29464
rect 79943 29504 79990 29546
rect 80114 29504 80158 29546
rect 80282 29504 80329 29546
rect 79943 29464 79952 29504
rect 80114 29464 80116 29504
rect 80156 29464 80158 29504
rect 80320 29464 80329 29504
rect 79943 29422 79990 29464
rect 80114 29422 80158 29464
rect 80282 29422 80329 29464
rect 95063 29504 95110 29546
rect 95234 29504 95278 29546
rect 95402 29504 95449 29546
rect 95063 29464 95072 29504
rect 95234 29464 95236 29504
rect 95276 29464 95278 29504
rect 95440 29464 95449 29504
rect 95063 29422 95110 29464
rect 95234 29422 95278 29464
rect 95402 29422 95449 29464
rect 3103 28748 3150 28790
rect 3274 28748 3318 28790
rect 3442 28748 3489 28790
rect 3103 28708 3112 28748
rect 3274 28708 3276 28748
rect 3316 28708 3318 28748
rect 3480 28708 3489 28748
rect 3103 28666 3150 28708
rect 3274 28666 3318 28708
rect 3442 28666 3489 28708
rect 18223 28748 18270 28790
rect 18394 28748 18438 28790
rect 18562 28748 18609 28790
rect 18223 28708 18232 28748
rect 18394 28708 18396 28748
rect 18436 28708 18438 28748
rect 18600 28708 18609 28748
rect 18223 28666 18270 28708
rect 18394 28666 18438 28708
rect 18562 28666 18609 28708
rect 33343 28748 33390 28790
rect 33514 28748 33558 28790
rect 33682 28748 33729 28790
rect 33343 28708 33352 28748
rect 33514 28708 33516 28748
rect 33556 28708 33558 28748
rect 33720 28708 33729 28748
rect 33343 28666 33390 28708
rect 33514 28666 33558 28708
rect 33682 28666 33729 28708
rect 48463 28748 48510 28790
rect 48634 28748 48678 28790
rect 48802 28748 48849 28790
rect 48463 28708 48472 28748
rect 48634 28708 48636 28748
rect 48676 28708 48678 28748
rect 48840 28708 48849 28748
rect 48463 28666 48510 28708
rect 48634 28666 48678 28708
rect 48802 28666 48849 28708
rect 63583 28748 63630 28790
rect 63754 28748 63798 28790
rect 63922 28748 63969 28790
rect 63583 28708 63592 28748
rect 63754 28708 63756 28748
rect 63796 28708 63798 28748
rect 63960 28708 63969 28748
rect 63583 28666 63630 28708
rect 63754 28666 63798 28708
rect 63922 28666 63969 28708
rect 78703 28748 78750 28790
rect 78874 28748 78918 28790
rect 79042 28748 79089 28790
rect 78703 28708 78712 28748
rect 78874 28708 78876 28748
rect 78916 28708 78918 28748
rect 79080 28708 79089 28748
rect 78703 28666 78750 28708
rect 78874 28666 78918 28708
rect 79042 28666 79089 28708
rect 93823 28748 93870 28790
rect 93994 28748 94038 28790
rect 94162 28748 94209 28790
rect 93823 28708 93832 28748
rect 93994 28708 93996 28748
rect 94036 28708 94038 28748
rect 94200 28708 94209 28748
rect 93823 28666 93870 28708
rect 93994 28666 94038 28708
rect 94162 28666 94209 28708
rect 4343 27992 4390 28034
rect 4514 27992 4558 28034
rect 4682 27992 4729 28034
rect 4343 27952 4352 27992
rect 4514 27952 4516 27992
rect 4556 27952 4558 27992
rect 4720 27952 4729 27992
rect 4343 27910 4390 27952
rect 4514 27910 4558 27952
rect 4682 27910 4729 27952
rect 19463 27992 19510 28034
rect 19634 27992 19678 28034
rect 19802 27992 19849 28034
rect 19463 27952 19472 27992
rect 19634 27952 19636 27992
rect 19676 27952 19678 27992
rect 19840 27952 19849 27992
rect 19463 27910 19510 27952
rect 19634 27910 19678 27952
rect 19802 27910 19849 27952
rect 34583 27992 34630 28034
rect 34754 27992 34798 28034
rect 34922 27992 34969 28034
rect 34583 27952 34592 27992
rect 34754 27952 34756 27992
rect 34796 27952 34798 27992
rect 34960 27952 34969 27992
rect 34583 27910 34630 27952
rect 34754 27910 34798 27952
rect 34922 27910 34969 27952
rect 49703 27992 49750 28034
rect 49874 27992 49918 28034
rect 50042 27992 50089 28034
rect 49703 27952 49712 27992
rect 49874 27952 49876 27992
rect 49916 27952 49918 27992
rect 50080 27952 50089 27992
rect 49703 27910 49750 27952
rect 49874 27910 49918 27952
rect 50042 27910 50089 27952
rect 64823 27992 64870 28034
rect 64994 27992 65038 28034
rect 65162 27992 65209 28034
rect 64823 27952 64832 27992
rect 64994 27952 64996 27992
rect 65036 27952 65038 27992
rect 65200 27952 65209 27992
rect 64823 27910 64870 27952
rect 64994 27910 65038 27952
rect 65162 27910 65209 27952
rect 79943 27992 79990 28034
rect 80114 27992 80158 28034
rect 80282 27992 80329 28034
rect 79943 27952 79952 27992
rect 80114 27952 80116 27992
rect 80156 27952 80158 27992
rect 80320 27952 80329 27992
rect 79943 27910 79990 27952
rect 80114 27910 80158 27952
rect 80282 27910 80329 27952
rect 95063 27992 95110 28034
rect 95234 27992 95278 28034
rect 95402 27992 95449 28034
rect 95063 27952 95072 27992
rect 95234 27952 95236 27992
rect 95276 27952 95278 27992
rect 95440 27952 95449 27992
rect 95063 27910 95110 27952
rect 95234 27910 95278 27952
rect 95402 27910 95449 27952
rect 3103 27236 3150 27278
rect 3274 27236 3318 27278
rect 3442 27236 3489 27278
rect 3103 27196 3112 27236
rect 3274 27196 3276 27236
rect 3316 27196 3318 27236
rect 3480 27196 3489 27236
rect 3103 27154 3150 27196
rect 3274 27154 3318 27196
rect 3442 27154 3489 27196
rect 18223 27236 18270 27278
rect 18394 27236 18438 27278
rect 18562 27236 18609 27278
rect 18223 27196 18232 27236
rect 18394 27196 18396 27236
rect 18436 27196 18438 27236
rect 18600 27196 18609 27236
rect 18223 27154 18270 27196
rect 18394 27154 18438 27196
rect 18562 27154 18609 27196
rect 33343 27236 33390 27278
rect 33514 27236 33558 27278
rect 33682 27236 33729 27278
rect 33343 27196 33352 27236
rect 33514 27196 33516 27236
rect 33556 27196 33558 27236
rect 33720 27196 33729 27236
rect 33343 27154 33390 27196
rect 33514 27154 33558 27196
rect 33682 27154 33729 27196
rect 48463 27236 48510 27278
rect 48634 27236 48678 27278
rect 48802 27236 48849 27278
rect 48463 27196 48472 27236
rect 48634 27196 48636 27236
rect 48676 27196 48678 27236
rect 48840 27196 48849 27236
rect 48463 27154 48510 27196
rect 48634 27154 48678 27196
rect 48802 27154 48849 27196
rect 63583 27236 63630 27278
rect 63754 27236 63798 27278
rect 63922 27236 63969 27278
rect 63583 27196 63592 27236
rect 63754 27196 63756 27236
rect 63796 27196 63798 27236
rect 63960 27196 63969 27236
rect 63583 27154 63630 27196
rect 63754 27154 63798 27196
rect 63922 27154 63969 27196
rect 78703 27236 78750 27278
rect 78874 27236 78918 27278
rect 79042 27236 79089 27278
rect 78703 27196 78712 27236
rect 78874 27196 78876 27236
rect 78916 27196 78918 27236
rect 79080 27196 79089 27236
rect 78703 27154 78750 27196
rect 78874 27154 78918 27196
rect 79042 27154 79089 27196
rect 93823 27236 93870 27278
rect 93994 27236 94038 27278
rect 94162 27236 94209 27278
rect 93823 27196 93832 27236
rect 93994 27196 93996 27236
rect 94036 27196 94038 27236
rect 94200 27196 94209 27236
rect 93823 27154 93870 27196
rect 93994 27154 94038 27196
rect 94162 27154 94209 27196
rect 4343 26480 4390 26522
rect 4514 26480 4558 26522
rect 4682 26480 4729 26522
rect 4343 26440 4352 26480
rect 4514 26440 4516 26480
rect 4556 26440 4558 26480
rect 4720 26440 4729 26480
rect 4343 26398 4390 26440
rect 4514 26398 4558 26440
rect 4682 26398 4729 26440
rect 19463 26480 19510 26522
rect 19634 26480 19678 26522
rect 19802 26480 19849 26522
rect 19463 26440 19472 26480
rect 19634 26440 19636 26480
rect 19676 26440 19678 26480
rect 19840 26440 19849 26480
rect 19463 26398 19510 26440
rect 19634 26398 19678 26440
rect 19802 26398 19849 26440
rect 34583 26480 34630 26522
rect 34754 26480 34798 26522
rect 34922 26480 34969 26522
rect 34583 26440 34592 26480
rect 34754 26440 34756 26480
rect 34796 26440 34798 26480
rect 34960 26440 34969 26480
rect 34583 26398 34630 26440
rect 34754 26398 34798 26440
rect 34922 26398 34969 26440
rect 49703 26480 49750 26522
rect 49874 26480 49918 26522
rect 50042 26480 50089 26522
rect 49703 26440 49712 26480
rect 49874 26440 49876 26480
rect 49916 26440 49918 26480
rect 50080 26440 50089 26480
rect 49703 26398 49750 26440
rect 49874 26398 49918 26440
rect 50042 26398 50089 26440
rect 64823 26480 64870 26522
rect 64994 26480 65038 26522
rect 65162 26480 65209 26522
rect 64823 26440 64832 26480
rect 64994 26440 64996 26480
rect 65036 26440 65038 26480
rect 65200 26440 65209 26480
rect 64823 26398 64870 26440
rect 64994 26398 65038 26440
rect 65162 26398 65209 26440
rect 79943 26480 79990 26522
rect 80114 26480 80158 26522
rect 80282 26480 80329 26522
rect 79943 26440 79952 26480
rect 80114 26440 80116 26480
rect 80156 26440 80158 26480
rect 80320 26440 80329 26480
rect 79943 26398 79990 26440
rect 80114 26398 80158 26440
rect 80282 26398 80329 26440
rect 95063 26480 95110 26522
rect 95234 26480 95278 26522
rect 95402 26480 95449 26522
rect 95063 26440 95072 26480
rect 95234 26440 95236 26480
rect 95276 26440 95278 26480
rect 95440 26440 95449 26480
rect 95063 26398 95110 26440
rect 95234 26398 95278 26440
rect 95402 26398 95449 26440
rect 3103 25724 3150 25766
rect 3274 25724 3318 25766
rect 3442 25724 3489 25766
rect 3103 25684 3112 25724
rect 3274 25684 3276 25724
rect 3316 25684 3318 25724
rect 3480 25684 3489 25724
rect 3103 25642 3150 25684
rect 3274 25642 3318 25684
rect 3442 25642 3489 25684
rect 18223 25724 18270 25766
rect 18394 25724 18438 25766
rect 18562 25724 18609 25766
rect 18223 25684 18232 25724
rect 18394 25684 18396 25724
rect 18436 25684 18438 25724
rect 18600 25684 18609 25724
rect 18223 25642 18270 25684
rect 18394 25642 18438 25684
rect 18562 25642 18609 25684
rect 33343 25724 33390 25766
rect 33514 25724 33558 25766
rect 33682 25724 33729 25766
rect 33343 25684 33352 25724
rect 33514 25684 33516 25724
rect 33556 25684 33558 25724
rect 33720 25684 33729 25724
rect 33343 25642 33390 25684
rect 33514 25642 33558 25684
rect 33682 25642 33729 25684
rect 48463 25724 48510 25766
rect 48634 25724 48678 25766
rect 48802 25724 48849 25766
rect 48463 25684 48472 25724
rect 48634 25684 48636 25724
rect 48676 25684 48678 25724
rect 48840 25684 48849 25724
rect 48463 25642 48510 25684
rect 48634 25642 48678 25684
rect 48802 25642 48849 25684
rect 63583 25724 63630 25766
rect 63754 25724 63798 25766
rect 63922 25724 63969 25766
rect 63583 25684 63592 25724
rect 63754 25684 63756 25724
rect 63796 25684 63798 25724
rect 63960 25684 63969 25724
rect 63583 25642 63630 25684
rect 63754 25642 63798 25684
rect 63922 25642 63969 25684
rect 78703 25724 78750 25766
rect 78874 25724 78918 25766
rect 79042 25724 79089 25766
rect 78703 25684 78712 25724
rect 78874 25684 78876 25724
rect 78916 25684 78918 25724
rect 79080 25684 79089 25724
rect 78703 25642 78750 25684
rect 78874 25642 78918 25684
rect 79042 25642 79089 25684
rect 93823 25724 93870 25766
rect 93994 25724 94038 25766
rect 94162 25724 94209 25766
rect 93823 25684 93832 25724
rect 93994 25684 93996 25724
rect 94036 25684 94038 25724
rect 94200 25684 94209 25724
rect 93823 25642 93870 25684
rect 93994 25642 94038 25684
rect 94162 25642 94209 25684
rect 4343 24968 4390 25010
rect 4514 24968 4558 25010
rect 4682 24968 4729 25010
rect 4343 24928 4352 24968
rect 4514 24928 4516 24968
rect 4556 24928 4558 24968
rect 4720 24928 4729 24968
rect 4343 24886 4390 24928
rect 4514 24886 4558 24928
rect 4682 24886 4729 24928
rect 19463 24968 19510 25010
rect 19634 24968 19678 25010
rect 19802 24968 19849 25010
rect 19463 24928 19472 24968
rect 19634 24928 19636 24968
rect 19676 24928 19678 24968
rect 19840 24928 19849 24968
rect 19463 24886 19510 24928
rect 19634 24886 19678 24928
rect 19802 24886 19849 24928
rect 34583 24968 34630 25010
rect 34754 24968 34798 25010
rect 34922 24968 34969 25010
rect 34583 24928 34592 24968
rect 34754 24928 34756 24968
rect 34796 24928 34798 24968
rect 34960 24928 34969 24968
rect 34583 24886 34630 24928
rect 34754 24886 34798 24928
rect 34922 24886 34969 24928
rect 49703 24968 49750 25010
rect 49874 24968 49918 25010
rect 50042 24968 50089 25010
rect 49703 24928 49712 24968
rect 49874 24928 49876 24968
rect 49916 24928 49918 24968
rect 50080 24928 50089 24968
rect 49703 24886 49750 24928
rect 49874 24886 49918 24928
rect 50042 24886 50089 24928
rect 64823 24968 64870 25010
rect 64994 24968 65038 25010
rect 65162 24968 65209 25010
rect 64823 24928 64832 24968
rect 64994 24928 64996 24968
rect 65036 24928 65038 24968
rect 65200 24928 65209 24968
rect 64823 24886 64870 24928
rect 64994 24886 65038 24928
rect 65162 24886 65209 24928
rect 79943 24968 79990 25010
rect 80114 24968 80158 25010
rect 80282 24968 80329 25010
rect 79943 24928 79952 24968
rect 80114 24928 80116 24968
rect 80156 24928 80158 24968
rect 80320 24928 80329 24968
rect 79943 24886 79990 24928
rect 80114 24886 80158 24928
rect 80282 24886 80329 24928
rect 95063 24968 95110 25010
rect 95234 24968 95278 25010
rect 95402 24968 95449 25010
rect 95063 24928 95072 24968
rect 95234 24928 95236 24968
rect 95276 24928 95278 24968
rect 95440 24928 95449 24968
rect 95063 24886 95110 24928
rect 95234 24886 95278 24928
rect 95402 24886 95449 24928
rect 3103 24212 3150 24254
rect 3274 24212 3318 24254
rect 3442 24212 3489 24254
rect 3103 24172 3112 24212
rect 3274 24172 3276 24212
rect 3316 24172 3318 24212
rect 3480 24172 3489 24212
rect 3103 24130 3150 24172
rect 3274 24130 3318 24172
rect 3442 24130 3489 24172
rect 18223 24212 18270 24254
rect 18394 24212 18438 24254
rect 18562 24212 18609 24254
rect 18223 24172 18232 24212
rect 18394 24172 18396 24212
rect 18436 24172 18438 24212
rect 18600 24172 18609 24212
rect 18223 24130 18270 24172
rect 18394 24130 18438 24172
rect 18562 24130 18609 24172
rect 33343 24212 33390 24254
rect 33514 24212 33558 24254
rect 33682 24212 33729 24254
rect 33343 24172 33352 24212
rect 33514 24172 33516 24212
rect 33556 24172 33558 24212
rect 33720 24172 33729 24212
rect 33343 24130 33390 24172
rect 33514 24130 33558 24172
rect 33682 24130 33729 24172
rect 48463 24212 48510 24254
rect 48634 24212 48678 24254
rect 48802 24212 48849 24254
rect 48463 24172 48472 24212
rect 48634 24172 48636 24212
rect 48676 24172 48678 24212
rect 48840 24172 48849 24212
rect 48463 24130 48510 24172
rect 48634 24130 48678 24172
rect 48802 24130 48849 24172
rect 63583 24212 63630 24254
rect 63754 24212 63798 24254
rect 63922 24212 63969 24254
rect 63583 24172 63592 24212
rect 63754 24172 63756 24212
rect 63796 24172 63798 24212
rect 63960 24172 63969 24212
rect 63583 24130 63630 24172
rect 63754 24130 63798 24172
rect 63922 24130 63969 24172
rect 78703 24212 78750 24254
rect 78874 24212 78918 24254
rect 79042 24212 79089 24254
rect 78703 24172 78712 24212
rect 78874 24172 78876 24212
rect 78916 24172 78918 24212
rect 79080 24172 79089 24212
rect 78703 24130 78750 24172
rect 78874 24130 78918 24172
rect 79042 24130 79089 24172
rect 93823 24212 93870 24254
rect 93994 24212 94038 24254
rect 94162 24212 94209 24254
rect 93823 24172 93832 24212
rect 93994 24172 93996 24212
rect 94036 24172 94038 24212
rect 94200 24172 94209 24212
rect 93823 24130 93870 24172
rect 93994 24130 94038 24172
rect 94162 24130 94209 24172
rect 4343 23456 4390 23498
rect 4514 23456 4558 23498
rect 4682 23456 4729 23498
rect 4343 23416 4352 23456
rect 4514 23416 4516 23456
rect 4556 23416 4558 23456
rect 4720 23416 4729 23456
rect 4343 23374 4390 23416
rect 4514 23374 4558 23416
rect 4682 23374 4729 23416
rect 19463 23456 19510 23498
rect 19634 23456 19678 23498
rect 19802 23456 19849 23498
rect 19463 23416 19472 23456
rect 19634 23416 19636 23456
rect 19676 23416 19678 23456
rect 19840 23416 19849 23456
rect 19463 23374 19510 23416
rect 19634 23374 19678 23416
rect 19802 23374 19849 23416
rect 34583 23456 34630 23498
rect 34754 23456 34798 23498
rect 34922 23456 34969 23498
rect 34583 23416 34592 23456
rect 34754 23416 34756 23456
rect 34796 23416 34798 23456
rect 34960 23416 34969 23456
rect 34583 23374 34630 23416
rect 34754 23374 34798 23416
rect 34922 23374 34969 23416
rect 49703 23456 49750 23498
rect 49874 23456 49918 23498
rect 50042 23456 50089 23498
rect 49703 23416 49712 23456
rect 49874 23416 49876 23456
rect 49916 23416 49918 23456
rect 50080 23416 50089 23456
rect 49703 23374 49750 23416
rect 49874 23374 49918 23416
rect 50042 23374 50089 23416
rect 64823 23456 64870 23498
rect 64994 23456 65038 23498
rect 65162 23456 65209 23498
rect 64823 23416 64832 23456
rect 64994 23416 64996 23456
rect 65036 23416 65038 23456
rect 65200 23416 65209 23456
rect 64823 23374 64870 23416
rect 64994 23374 65038 23416
rect 65162 23374 65209 23416
rect 79943 23456 79990 23498
rect 80114 23456 80158 23498
rect 80282 23456 80329 23498
rect 79943 23416 79952 23456
rect 80114 23416 80116 23456
rect 80156 23416 80158 23456
rect 80320 23416 80329 23456
rect 79943 23374 79990 23416
rect 80114 23374 80158 23416
rect 80282 23374 80329 23416
rect 95063 23456 95110 23498
rect 95234 23456 95278 23498
rect 95402 23456 95449 23498
rect 95063 23416 95072 23456
rect 95234 23416 95236 23456
rect 95276 23416 95278 23456
rect 95440 23416 95449 23456
rect 95063 23374 95110 23416
rect 95234 23374 95278 23416
rect 95402 23374 95449 23416
rect 3103 22700 3150 22742
rect 3274 22700 3318 22742
rect 3442 22700 3489 22742
rect 3103 22660 3112 22700
rect 3274 22660 3276 22700
rect 3316 22660 3318 22700
rect 3480 22660 3489 22700
rect 3103 22618 3150 22660
rect 3274 22618 3318 22660
rect 3442 22618 3489 22660
rect 18223 22700 18270 22742
rect 18394 22700 18438 22742
rect 18562 22700 18609 22742
rect 18223 22660 18232 22700
rect 18394 22660 18396 22700
rect 18436 22660 18438 22700
rect 18600 22660 18609 22700
rect 18223 22618 18270 22660
rect 18394 22618 18438 22660
rect 18562 22618 18609 22660
rect 33343 22700 33390 22742
rect 33514 22700 33558 22742
rect 33682 22700 33729 22742
rect 33343 22660 33352 22700
rect 33514 22660 33516 22700
rect 33556 22660 33558 22700
rect 33720 22660 33729 22700
rect 33343 22618 33390 22660
rect 33514 22618 33558 22660
rect 33682 22618 33729 22660
rect 48463 22700 48510 22742
rect 48634 22700 48678 22742
rect 48802 22700 48849 22742
rect 48463 22660 48472 22700
rect 48634 22660 48636 22700
rect 48676 22660 48678 22700
rect 48840 22660 48849 22700
rect 48463 22618 48510 22660
rect 48634 22618 48678 22660
rect 48802 22618 48849 22660
rect 63583 22700 63630 22742
rect 63754 22700 63798 22742
rect 63922 22700 63969 22742
rect 63583 22660 63592 22700
rect 63754 22660 63756 22700
rect 63796 22660 63798 22700
rect 63960 22660 63969 22700
rect 63583 22618 63630 22660
rect 63754 22618 63798 22660
rect 63922 22618 63969 22660
rect 78703 22700 78750 22742
rect 78874 22700 78918 22742
rect 79042 22700 79089 22742
rect 78703 22660 78712 22700
rect 78874 22660 78876 22700
rect 78916 22660 78918 22700
rect 79080 22660 79089 22700
rect 78703 22618 78750 22660
rect 78874 22618 78918 22660
rect 79042 22618 79089 22660
rect 93823 22700 93870 22742
rect 93994 22700 94038 22742
rect 94162 22700 94209 22742
rect 93823 22660 93832 22700
rect 93994 22660 93996 22700
rect 94036 22660 94038 22700
rect 94200 22660 94209 22700
rect 93823 22618 93870 22660
rect 93994 22618 94038 22660
rect 94162 22618 94209 22660
rect 4343 21944 4390 21986
rect 4514 21944 4558 21986
rect 4682 21944 4729 21986
rect 4343 21904 4352 21944
rect 4514 21904 4516 21944
rect 4556 21904 4558 21944
rect 4720 21904 4729 21944
rect 4343 21862 4390 21904
rect 4514 21862 4558 21904
rect 4682 21862 4729 21904
rect 19463 21944 19510 21986
rect 19634 21944 19678 21986
rect 19802 21944 19849 21986
rect 19463 21904 19472 21944
rect 19634 21904 19636 21944
rect 19676 21904 19678 21944
rect 19840 21904 19849 21944
rect 19463 21862 19510 21904
rect 19634 21862 19678 21904
rect 19802 21862 19849 21904
rect 34583 21944 34630 21986
rect 34754 21944 34798 21986
rect 34922 21944 34969 21986
rect 34583 21904 34592 21944
rect 34754 21904 34756 21944
rect 34796 21904 34798 21944
rect 34960 21904 34969 21944
rect 34583 21862 34630 21904
rect 34754 21862 34798 21904
rect 34922 21862 34969 21904
rect 49703 21944 49750 21986
rect 49874 21944 49918 21986
rect 50042 21944 50089 21986
rect 49703 21904 49712 21944
rect 49874 21904 49876 21944
rect 49916 21904 49918 21944
rect 50080 21904 50089 21944
rect 49703 21862 49750 21904
rect 49874 21862 49918 21904
rect 50042 21862 50089 21904
rect 64823 21944 64870 21986
rect 64994 21944 65038 21986
rect 65162 21944 65209 21986
rect 64823 21904 64832 21944
rect 64994 21904 64996 21944
rect 65036 21904 65038 21944
rect 65200 21904 65209 21944
rect 64823 21862 64870 21904
rect 64994 21862 65038 21904
rect 65162 21862 65209 21904
rect 79943 21944 79990 21986
rect 80114 21944 80158 21986
rect 80282 21944 80329 21986
rect 79943 21904 79952 21944
rect 80114 21904 80116 21944
rect 80156 21904 80158 21944
rect 80320 21904 80329 21944
rect 79943 21862 79990 21904
rect 80114 21862 80158 21904
rect 80282 21862 80329 21904
rect 95063 21944 95110 21986
rect 95234 21944 95278 21986
rect 95402 21944 95449 21986
rect 95063 21904 95072 21944
rect 95234 21904 95236 21944
rect 95276 21904 95278 21944
rect 95440 21904 95449 21944
rect 95063 21862 95110 21904
rect 95234 21862 95278 21904
rect 95402 21862 95449 21904
rect 3103 21188 3150 21230
rect 3274 21188 3318 21230
rect 3442 21188 3489 21230
rect 3103 21148 3112 21188
rect 3274 21148 3276 21188
rect 3316 21148 3318 21188
rect 3480 21148 3489 21188
rect 3103 21106 3150 21148
rect 3274 21106 3318 21148
rect 3442 21106 3489 21148
rect 18223 21188 18270 21230
rect 18394 21188 18438 21230
rect 18562 21188 18609 21230
rect 18223 21148 18232 21188
rect 18394 21148 18396 21188
rect 18436 21148 18438 21188
rect 18600 21148 18609 21188
rect 18223 21106 18270 21148
rect 18394 21106 18438 21148
rect 18562 21106 18609 21148
rect 33343 21188 33390 21230
rect 33514 21188 33558 21230
rect 33682 21188 33729 21230
rect 33343 21148 33352 21188
rect 33514 21148 33516 21188
rect 33556 21148 33558 21188
rect 33720 21148 33729 21188
rect 33343 21106 33390 21148
rect 33514 21106 33558 21148
rect 33682 21106 33729 21148
rect 48463 21188 48510 21230
rect 48634 21188 48678 21230
rect 48802 21188 48849 21230
rect 48463 21148 48472 21188
rect 48634 21148 48636 21188
rect 48676 21148 48678 21188
rect 48840 21148 48849 21188
rect 48463 21106 48510 21148
rect 48634 21106 48678 21148
rect 48802 21106 48849 21148
rect 63583 21188 63630 21230
rect 63754 21188 63798 21230
rect 63922 21188 63969 21230
rect 63583 21148 63592 21188
rect 63754 21148 63756 21188
rect 63796 21148 63798 21188
rect 63960 21148 63969 21188
rect 63583 21106 63630 21148
rect 63754 21106 63798 21148
rect 63922 21106 63969 21148
rect 78703 21188 78750 21230
rect 78874 21188 78918 21230
rect 79042 21188 79089 21230
rect 78703 21148 78712 21188
rect 78874 21148 78876 21188
rect 78916 21148 78918 21188
rect 79080 21148 79089 21188
rect 78703 21106 78750 21148
rect 78874 21106 78918 21148
rect 79042 21106 79089 21148
rect 93823 21188 93870 21230
rect 93994 21188 94038 21230
rect 94162 21188 94209 21230
rect 93823 21148 93832 21188
rect 93994 21148 93996 21188
rect 94036 21148 94038 21188
rect 94200 21148 94209 21188
rect 93823 21106 93870 21148
rect 93994 21106 94038 21148
rect 94162 21106 94209 21148
rect 4343 20432 4390 20474
rect 4514 20432 4558 20474
rect 4682 20432 4729 20474
rect 4343 20392 4352 20432
rect 4514 20392 4516 20432
rect 4556 20392 4558 20432
rect 4720 20392 4729 20432
rect 4343 20350 4390 20392
rect 4514 20350 4558 20392
rect 4682 20350 4729 20392
rect 19463 20432 19510 20474
rect 19634 20432 19678 20474
rect 19802 20432 19849 20474
rect 19463 20392 19472 20432
rect 19634 20392 19636 20432
rect 19676 20392 19678 20432
rect 19840 20392 19849 20432
rect 19463 20350 19510 20392
rect 19634 20350 19678 20392
rect 19802 20350 19849 20392
rect 34583 20432 34630 20474
rect 34754 20432 34798 20474
rect 34922 20432 34969 20474
rect 34583 20392 34592 20432
rect 34754 20392 34756 20432
rect 34796 20392 34798 20432
rect 34960 20392 34969 20432
rect 34583 20350 34630 20392
rect 34754 20350 34798 20392
rect 34922 20350 34969 20392
rect 49703 20432 49750 20474
rect 49874 20432 49918 20474
rect 50042 20432 50089 20474
rect 49703 20392 49712 20432
rect 49874 20392 49876 20432
rect 49916 20392 49918 20432
rect 50080 20392 50089 20432
rect 49703 20350 49750 20392
rect 49874 20350 49918 20392
rect 50042 20350 50089 20392
rect 64823 20432 64870 20474
rect 64994 20432 65038 20474
rect 65162 20432 65209 20474
rect 64823 20392 64832 20432
rect 64994 20392 64996 20432
rect 65036 20392 65038 20432
rect 65200 20392 65209 20432
rect 64823 20350 64870 20392
rect 64994 20350 65038 20392
rect 65162 20350 65209 20392
rect 79943 20432 79990 20474
rect 80114 20432 80158 20474
rect 80282 20432 80329 20474
rect 79943 20392 79952 20432
rect 80114 20392 80116 20432
rect 80156 20392 80158 20432
rect 80320 20392 80329 20432
rect 79943 20350 79990 20392
rect 80114 20350 80158 20392
rect 80282 20350 80329 20392
rect 95063 20432 95110 20474
rect 95234 20432 95278 20474
rect 95402 20432 95449 20474
rect 95063 20392 95072 20432
rect 95234 20392 95236 20432
rect 95276 20392 95278 20432
rect 95440 20392 95449 20432
rect 95063 20350 95110 20392
rect 95234 20350 95278 20392
rect 95402 20350 95449 20392
rect 3103 19676 3150 19718
rect 3274 19676 3318 19718
rect 3442 19676 3489 19718
rect 3103 19636 3112 19676
rect 3274 19636 3276 19676
rect 3316 19636 3318 19676
rect 3480 19636 3489 19676
rect 3103 19594 3150 19636
rect 3274 19594 3318 19636
rect 3442 19594 3489 19636
rect 18223 19676 18270 19718
rect 18394 19676 18438 19718
rect 18562 19676 18609 19718
rect 18223 19636 18232 19676
rect 18394 19636 18396 19676
rect 18436 19636 18438 19676
rect 18600 19636 18609 19676
rect 18223 19594 18270 19636
rect 18394 19594 18438 19636
rect 18562 19594 18609 19636
rect 33343 19676 33390 19718
rect 33514 19676 33558 19718
rect 33682 19676 33729 19718
rect 33343 19636 33352 19676
rect 33514 19636 33516 19676
rect 33556 19636 33558 19676
rect 33720 19636 33729 19676
rect 33343 19594 33390 19636
rect 33514 19594 33558 19636
rect 33682 19594 33729 19636
rect 48463 19676 48510 19718
rect 48634 19676 48678 19718
rect 48802 19676 48849 19718
rect 48463 19636 48472 19676
rect 48634 19636 48636 19676
rect 48676 19636 48678 19676
rect 48840 19636 48849 19676
rect 48463 19594 48510 19636
rect 48634 19594 48678 19636
rect 48802 19594 48849 19636
rect 63583 19676 63630 19718
rect 63754 19676 63798 19718
rect 63922 19676 63969 19718
rect 63583 19636 63592 19676
rect 63754 19636 63756 19676
rect 63796 19636 63798 19676
rect 63960 19636 63969 19676
rect 63583 19594 63630 19636
rect 63754 19594 63798 19636
rect 63922 19594 63969 19636
rect 78703 19676 78750 19718
rect 78874 19676 78918 19718
rect 79042 19676 79089 19718
rect 78703 19636 78712 19676
rect 78874 19636 78876 19676
rect 78916 19636 78918 19676
rect 79080 19636 79089 19676
rect 78703 19594 78750 19636
rect 78874 19594 78918 19636
rect 79042 19594 79089 19636
rect 93823 19676 93870 19718
rect 93994 19676 94038 19718
rect 94162 19676 94209 19718
rect 93823 19636 93832 19676
rect 93994 19636 93996 19676
rect 94036 19636 94038 19676
rect 94200 19636 94209 19676
rect 93823 19594 93870 19636
rect 93994 19594 94038 19636
rect 94162 19594 94209 19636
rect 4343 18920 4390 18962
rect 4514 18920 4558 18962
rect 4682 18920 4729 18962
rect 4343 18880 4352 18920
rect 4514 18880 4516 18920
rect 4556 18880 4558 18920
rect 4720 18880 4729 18920
rect 4343 18838 4390 18880
rect 4514 18838 4558 18880
rect 4682 18838 4729 18880
rect 19463 18920 19510 18962
rect 19634 18920 19678 18962
rect 19802 18920 19849 18962
rect 19463 18880 19472 18920
rect 19634 18880 19636 18920
rect 19676 18880 19678 18920
rect 19840 18880 19849 18920
rect 19463 18838 19510 18880
rect 19634 18838 19678 18880
rect 19802 18838 19849 18880
rect 34583 18920 34630 18962
rect 34754 18920 34798 18962
rect 34922 18920 34969 18962
rect 34583 18880 34592 18920
rect 34754 18880 34756 18920
rect 34796 18880 34798 18920
rect 34960 18880 34969 18920
rect 34583 18838 34630 18880
rect 34754 18838 34798 18880
rect 34922 18838 34969 18880
rect 49703 18920 49750 18962
rect 49874 18920 49918 18962
rect 50042 18920 50089 18962
rect 49703 18880 49712 18920
rect 49874 18880 49876 18920
rect 49916 18880 49918 18920
rect 50080 18880 50089 18920
rect 49703 18838 49750 18880
rect 49874 18838 49918 18880
rect 50042 18838 50089 18880
rect 64823 18920 64870 18962
rect 64994 18920 65038 18962
rect 65162 18920 65209 18962
rect 64823 18880 64832 18920
rect 64994 18880 64996 18920
rect 65036 18880 65038 18920
rect 65200 18880 65209 18920
rect 64823 18838 64870 18880
rect 64994 18838 65038 18880
rect 65162 18838 65209 18880
rect 79943 18920 79990 18962
rect 80114 18920 80158 18962
rect 80282 18920 80329 18962
rect 79943 18880 79952 18920
rect 80114 18880 80116 18920
rect 80156 18880 80158 18920
rect 80320 18880 80329 18920
rect 79943 18838 79990 18880
rect 80114 18838 80158 18880
rect 80282 18838 80329 18880
rect 95063 18920 95110 18962
rect 95234 18920 95278 18962
rect 95402 18920 95449 18962
rect 95063 18880 95072 18920
rect 95234 18880 95236 18920
rect 95276 18880 95278 18920
rect 95440 18880 95449 18920
rect 95063 18838 95110 18880
rect 95234 18838 95278 18880
rect 95402 18838 95449 18880
rect 3103 18164 3150 18206
rect 3274 18164 3318 18206
rect 3442 18164 3489 18206
rect 3103 18124 3112 18164
rect 3274 18124 3276 18164
rect 3316 18124 3318 18164
rect 3480 18124 3489 18164
rect 3103 18082 3150 18124
rect 3274 18082 3318 18124
rect 3442 18082 3489 18124
rect 18223 18164 18270 18206
rect 18394 18164 18438 18206
rect 18562 18164 18609 18206
rect 18223 18124 18232 18164
rect 18394 18124 18396 18164
rect 18436 18124 18438 18164
rect 18600 18124 18609 18164
rect 18223 18082 18270 18124
rect 18394 18082 18438 18124
rect 18562 18082 18609 18124
rect 33343 18164 33390 18206
rect 33514 18164 33558 18206
rect 33682 18164 33729 18206
rect 33343 18124 33352 18164
rect 33514 18124 33516 18164
rect 33556 18124 33558 18164
rect 33720 18124 33729 18164
rect 33343 18082 33390 18124
rect 33514 18082 33558 18124
rect 33682 18082 33729 18124
rect 48463 18164 48510 18206
rect 48634 18164 48678 18206
rect 48802 18164 48849 18206
rect 48463 18124 48472 18164
rect 48634 18124 48636 18164
rect 48676 18124 48678 18164
rect 48840 18124 48849 18164
rect 48463 18082 48510 18124
rect 48634 18082 48678 18124
rect 48802 18082 48849 18124
rect 63583 18164 63630 18206
rect 63754 18164 63798 18206
rect 63922 18164 63969 18206
rect 63583 18124 63592 18164
rect 63754 18124 63756 18164
rect 63796 18124 63798 18164
rect 63960 18124 63969 18164
rect 63583 18082 63630 18124
rect 63754 18082 63798 18124
rect 63922 18082 63969 18124
rect 78703 18164 78750 18206
rect 78874 18164 78918 18206
rect 79042 18164 79089 18206
rect 78703 18124 78712 18164
rect 78874 18124 78876 18164
rect 78916 18124 78918 18164
rect 79080 18124 79089 18164
rect 78703 18082 78750 18124
rect 78874 18082 78918 18124
rect 79042 18082 79089 18124
rect 93823 18164 93870 18206
rect 93994 18164 94038 18206
rect 94162 18164 94209 18206
rect 93823 18124 93832 18164
rect 93994 18124 93996 18164
rect 94036 18124 94038 18164
rect 94200 18124 94209 18164
rect 93823 18082 93870 18124
rect 93994 18082 94038 18124
rect 94162 18082 94209 18124
rect 4343 17408 4390 17450
rect 4514 17408 4558 17450
rect 4682 17408 4729 17450
rect 4343 17368 4352 17408
rect 4514 17368 4516 17408
rect 4556 17368 4558 17408
rect 4720 17368 4729 17408
rect 4343 17326 4390 17368
rect 4514 17326 4558 17368
rect 4682 17326 4729 17368
rect 19463 17408 19510 17450
rect 19634 17408 19678 17450
rect 19802 17408 19849 17450
rect 19463 17368 19472 17408
rect 19634 17368 19636 17408
rect 19676 17368 19678 17408
rect 19840 17368 19849 17408
rect 19463 17326 19510 17368
rect 19634 17326 19678 17368
rect 19802 17326 19849 17368
rect 34583 17408 34630 17450
rect 34754 17408 34798 17450
rect 34922 17408 34969 17450
rect 34583 17368 34592 17408
rect 34754 17368 34756 17408
rect 34796 17368 34798 17408
rect 34960 17368 34969 17408
rect 34583 17326 34630 17368
rect 34754 17326 34798 17368
rect 34922 17326 34969 17368
rect 49703 17408 49750 17450
rect 49874 17408 49918 17450
rect 50042 17408 50089 17450
rect 49703 17368 49712 17408
rect 49874 17368 49876 17408
rect 49916 17368 49918 17408
rect 50080 17368 50089 17408
rect 49703 17326 49750 17368
rect 49874 17326 49918 17368
rect 50042 17326 50089 17368
rect 64823 17408 64870 17450
rect 64994 17408 65038 17450
rect 65162 17408 65209 17450
rect 64823 17368 64832 17408
rect 64994 17368 64996 17408
rect 65036 17368 65038 17408
rect 65200 17368 65209 17408
rect 64823 17326 64870 17368
rect 64994 17326 65038 17368
rect 65162 17326 65209 17368
rect 79943 17408 79990 17450
rect 80114 17408 80158 17450
rect 80282 17408 80329 17450
rect 79943 17368 79952 17408
rect 80114 17368 80116 17408
rect 80156 17368 80158 17408
rect 80320 17368 80329 17408
rect 79943 17326 79990 17368
rect 80114 17326 80158 17368
rect 80282 17326 80329 17368
rect 95063 17408 95110 17450
rect 95234 17408 95278 17450
rect 95402 17408 95449 17450
rect 95063 17368 95072 17408
rect 95234 17368 95236 17408
rect 95276 17368 95278 17408
rect 95440 17368 95449 17408
rect 95063 17326 95110 17368
rect 95234 17326 95278 17368
rect 95402 17326 95449 17368
rect 3103 16652 3150 16694
rect 3274 16652 3318 16694
rect 3442 16652 3489 16694
rect 3103 16612 3112 16652
rect 3274 16612 3276 16652
rect 3316 16612 3318 16652
rect 3480 16612 3489 16652
rect 3103 16570 3150 16612
rect 3274 16570 3318 16612
rect 3442 16570 3489 16612
rect 18223 16652 18270 16694
rect 18394 16652 18438 16694
rect 18562 16652 18609 16694
rect 18223 16612 18232 16652
rect 18394 16612 18396 16652
rect 18436 16612 18438 16652
rect 18600 16612 18609 16652
rect 18223 16570 18270 16612
rect 18394 16570 18438 16612
rect 18562 16570 18609 16612
rect 33343 16652 33390 16694
rect 33514 16652 33558 16694
rect 33682 16652 33729 16694
rect 33343 16612 33352 16652
rect 33514 16612 33516 16652
rect 33556 16612 33558 16652
rect 33720 16612 33729 16652
rect 33343 16570 33390 16612
rect 33514 16570 33558 16612
rect 33682 16570 33729 16612
rect 48463 16652 48510 16694
rect 48634 16652 48678 16694
rect 48802 16652 48849 16694
rect 48463 16612 48472 16652
rect 48634 16612 48636 16652
rect 48676 16612 48678 16652
rect 48840 16612 48849 16652
rect 48463 16570 48510 16612
rect 48634 16570 48678 16612
rect 48802 16570 48849 16612
rect 63583 16652 63630 16694
rect 63754 16652 63798 16694
rect 63922 16652 63969 16694
rect 63583 16612 63592 16652
rect 63754 16612 63756 16652
rect 63796 16612 63798 16652
rect 63960 16612 63969 16652
rect 63583 16570 63630 16612
rect 63754 16570 63798 16612
rect 63922 16570 63969 16612
rect 78703 16652 78750 16694
rect 78874 16652 78918 16694
rect 79042 16652 79089 16694
rect 78703 16612 78712 16652
rect 78874 16612 78876 16652
rect 78916 16612 78918 16652
rect 79080 16612 79089 16652
rect 78703 16570 78750 16612
rect 78874 16570 78918 16612
rect 79042 16570 79089 16612
rect 93823 16652 93870 16694
rect 93994 16652 94038 16694
rect 94162 16652 94209 16694
rect 93823 16612 93832 16652
rect 93994 16612 93996 16652
rect 94036 16612 94038 16652
rect 94200 16612 94209 16652
rect 93823 16570 93870 16612
rect 93994 16570 94038 16612
rect 94162 16570 94209 16612
rect 4343 15896 4390 15938
rect 4514 15896 4558 15938
rect 4682 15896 4729 15938
rect 4343 15856 4352 15896
rect 4514 15856 4516 15896
rect 4556 15856 4558 15896
rect 4720 15856 4729 15896
rect 4343 15814 4390 15856
rect 4514 15814 4558 15856
rect 4682 15814 4729 15856
rect 19463 15896 19510 15938
rect 19634 15896 19678 15938
rect 19802 15896 19849 15938
rect 19463 15856 19472 15896
rect 19634 15856 19636 15896
rect 19676 15856 19678 15896
rect 19840 15856 19849 15896
rect 19463 15814 19510 15856
rect 19634 15814 19678 15856
rect 19802 15814 19849 15856
rect 34583 15896 34630 15938
rect 34754 15896 34798 15938
rect 34922 15896 34969 15938
rect 34583 15856 34592 15896
rect 34754 15856 34756 15896
rect 34796 15856 34798 15896
rect 34960 15856 34969 15896
rect 34583 15814 34630 15856
rect 34754 15814 34798 15856
rect 34922 15814 34969 15856
rect 49703 15896 49750 15938
rect 49874 15896 49918 15938
rect 50042 15896 50089 15938
rect 49703 15856 49712 15896
rect 49874 15856 49876 15896
rect 49916 15856 49918 15896
rect 50080 15856 50089 15896
rect 49703 15814 49750 15856
rect 49874 15814 49918 15856
rect 50042 15814 50089 15856
rect 64823 15896 64870 15938
rect 64994 15896 65038 15938
rect 65162 15896 65209 15938
rect 64823 15856 64832 15896
rect 64994 15856 64996 15896
rect 65036 15856 65038 15896
rect 65200 15856 65209 15896
rect 64823 15814 64870 15856
rect 64994 15814 65038 15856
rect 65162 15814 65209 15856
rect 79943 15896 79990 15938
rect 80114 15896 80158 15938
rect 80282 15896 80329 15938
rect 79943 15856 79952 15896
rect 80114 15856 80116 15896
rect 80156 15856 80158 15896
rect 80320 15856 80329 15896
rect 79943 15814 79990 15856
rect 80114 15814 80158 15856
rect 80282 15814 80329 15856
rect 95063 15896 95110 15938
rect 95234 15896 95278 15938
rect 95402 15896 95449 15938
rect 95063 15856 95072 15896
rect 95234 15856 95236 15896
rect 95276 15856 95278 15896
rect 95440 15856 95449 15896
rect 95063 15814 95110 15856
rect 95234 15814 95278 15856
rect 95402 15814 95449 15856
rect 3103 15140 3150 15182
rect 3274 15140 3318 15182
rect 3442 15140 3489 15182
rect 3103 15100 3112 15140
rect 3274 15100 3276 15140
rect 3316 15100 3318 15140
rect 3480 15100 3489 15140
rect 3103 15058 3150 15100
rect 3274 15058 3318 15100
rect 3442 15058 3489 15100
rect 18223 15140 18270 15182
rect 18394 15140 18438 15182
rect 18562 15140 18609 15182
rect 18223 15100 18232 15140
rect 18394 15100 18396 15140
rect 18436 15100 18438 15140
rect 18600 15100 18609 15140
rect 18223 15058 18270 15100
rect 18394 15058 18438 15100
rect 18562 15058 18609 15100
rect 33343 15140 33390 15182
rect 33514 15140 33558 15182
rect 33682 15140 33729 15182
rect 33343 15100 33352 15140
rect 33514 15100 33516 15140
rect 33556 15100 33558 15140
rect 33720 15100 33729 15140
rect 33343 15058 33390 15100
rect 33514 15058 33558 15100
rect 33682 15058 33729 15100
rect 48463 15140 48510 15182
rect 48634 15140 48678 15182
rect 48802 15140 48849 15182
rect 48463 15100 48472 15140
rect 48634 15100 48636 15140
rect 48676 15100 48678 15140
rect 48840 15100 48849 15140
rect 48463 15058 48510 15100
rect 48634 15058 48678 15100
rect 48802 15058 48849 15100
rect 63583 15140 63630 15182
rect 63754 15140 63798 15182
rect 63922 15140 63969 15182
rect 63583 15100 63592 15140
rect 63754 15100 63756 15140
rect 63796 15100 63798 15140
rect 63960 15100 63969 15140
rect 63583 15058 63630 15100
rect 63754 15058 63798 15100
rect 63922 15058 63969 15100
rect 78703 15140 78750 15182
rect 78874 15140 78918 15182
rect 79042 15140 79089 15182
rect 78703 15100 78712 15140
rect 78874 15100 78876 15140
rect 78916 15100 78918 15140
rect 79080 15100 79089 15140
rect 78703 15058 78750 15100
rect 78874 15058 78918 15100
rect 79042 15058 79089 15100
rect 93823 15140 93870 15182
rect 93994 15140 94038 15182
rect 94162 15140 94209 15182
rect 93823 15100 93832 15140
rect 93994 15100 93996 15140
rect 94036 15100 94038 15140
rect 94200 15100 94209 15140
rect 93823 15058 93870 15100
rect 93994 15058 94038 15100
rect 94162 15058 94209 15100
rect 4343 14384 4390 14426
rect 4514 14384 4558 14426
rect 4682 14384 4729 14426
rect 4343 14344 4352 14384
rect 4514 14344 4516 14384
rect 4556 14344 4558 14384
rect 4720 14344 4729 14384
rect 4343 14302 4390 14344
rect 4514 14302 4558 14344
rect 4682 14302 4729 14344
rect 19463 14384 19510 14426
rect 19634 14384 19678 14426
rect 19802 14384 19849 14426
rect 19463 14344 19472 14384
rect 19634 14344 19636 14384
rect 19676 14344 19678 14384
rect 19840 14344 19849 14384
rect 19463 14302 19510 14344
rect 19634 14302 19678 14344
rect 19802 14302 19849 14344
rect 34583 14384 34630 14426
rect 34754 14384 34798 14426
rect 34922 14384 34969 14426
rect 34583 14344 34592 14384
rect 34754 14344 34756 14384
rect 34796 14344 34798 14384
rect 34960 14344 34969 14384
rect 34583 14302 34630 14344
rect 34754 14302 34798 14344
rect 34922 14302 34969 14344
rect 49703 14384 49750 14426
rect 49874 14384 49918 14426
rect 50042 14384 50089 14426
rect 49703 14344 49712 14384
rect 49874 14344 49876 14384
rect 49916 14344 49918 14384
rect 50080 14344 50089 14384
rect 49703 14302 49750 14344
rect 49874 14302 49918 14344
rect 50042 14302 50089 14344
rect 64823 14384 64870 14426
rect 64994 14384 65038 14426
rect 65162 14384 65209 14426
rect 64823 14344 64832 14384
rect 64994 14344 64996 14384
rect 65036 14344 65038 14384
rect 65200 14344 65209 14384
rect 64823 14302 64870 14344
rect 64994 14302 65038 14344
rect 65162 14302 65209 14344
rect 79943 14384 79990 14426
rect 80114 14384 80158 14426
rect 80282 14384 80329 14426
rect 79943 14344 79952 14384
rect 80114 14344 80116 14384
rect 80156 14344 80158 14384
rect 80320 14344 80329 14384
rect 79943 14302 79990 14344
rect 80114 14302 80158 14344
rect 80282 14302 80329 14344
rect 95063 14384 95110 14426
rect 95234 14384 95278 14426
rect 95402 14384 95449 14426
rect 95063 14344 95072 14384
rect 95234 14344 95236 14384
rect 95276 14344 95278 14384
rect 95440 14344 95449 14384
rect 95063 14302 95110 14344
rect 95234 14302 95278 14344
rect 95402 14302 95449 14344
rect 3103 13628 3150 13670
rect 3274 13628 3318 13670
rect 3442 13628 3489 13670
rect 3103 13588 3112 13628
rect 3274 13588 3276 13628
rect 3316 13588 3318 13628
rect 3480 13588 3489 13628
rect 3103 13546 3150 13588
rect 3274 13546 3318 13588
rect 3442 13546 3489 13588
rect 18223 13628 18270 13670
rect 18394 13628 18438 13670
rect 18562 13628 18609 13670
rect 18223 13588 18232 13628
rect 18394 13588 18396 13628
rect 18436 13588 18438 13628
rect 18600 13588 18609 13628
rect 18223 13546 18270 13588
rect 18394 13546 18438 13588
rect 18562 13546 18609 13588
rect 33343 13628 33390 13670
rect 33514 13628 33558 13670
rect 33682 13628 33729 13670
rect 33343 13588 33352 13628
rect 33514 13588 33516 13628
rect 33556 13588 33558 13628
rect 33720 13588 33729 13628
rect 33343 13546 33390 13588
rect 33514 13546 33558 13588
rect 33682 13546 33729 13588
rect 48463 13628 48510 13670
rect 48634 13628 48678 13670
rect 48802 13628 48849 13670
rect 48463 13588 48472 13628
rect 48634 13588 48636 13628
rect 48676 13588 48678 13628
rect 48840 13588 48849 13628
rect 48463 13546 48510 13588
rect 48634 13546 48678 13588
rect 48802 13546 48849 13588
rect 63583 13628 63630 13670
rect 63754 13628 63798 13670
rect 63922 13628 63969 13670
rect 63583 13588 63592 13628
rect 63754 13588 63756 13628
rect 63796 13588 63798 13628
rect 63960 13588 63969 13628
rect 63583 13546 63630 13588
rect 63754 13546 63798 13588
rect 63922 13546 63969 13588
rect 78703 13628 78750 13670
rect 78874 13628 78918 13670
rect 79042 13628 79089 13670
rect 78703 13588 78712 13628
rect 78874 13588 78876 13628
rect 78916 13588 78918 13628
rect 79080 13588 79089 13628
rect 78703 13546 78750 13588
rect 78874 13546 78918 13588
rect 79042 13546 79089 13588
rect 93823 13628 93870 13670
rect 93994 13628 94038 13670
rect 94162 13628 94209 13670
rect 93823 13588 93832 13628
rect 93994 13588 93996 13628
rect 94036 13588 94038 13628
rect 94200 13588 94209 13628
rect 93823 13546 93870 13588
rect 93994 13546 94038 13588
rect 94162 13546 94209 13588
rect 4343 12872 4390 12914
rect 4514 12872 4558 12914
rect 4682 12872 4729 12914
rect 4343 12832 4352 12872
rect 4514 12832 4516 12872
rect 4556 12832 4558 12872
rect 4720 12832 4729 12872
rect 4343 12790 4390 12832
rect 4514 12790 4558 12832
rect 4682 12790 4729 12832
rect 19463 12872 19510 12914
rect 19634 12872 19678 12914
rect 19802 12872 19849 12914
rect 19463 12832 19472 12872
rect 19634 12832 19636 12872
rect 19676 12832 19678 12872
rect 19840 12832 19849 12872
rect 19463 12790 19510 12832
rect 19634 12790 19678 12832
rect 19802 12790 19849 12832
rect 34583 12872 34630 12914
rect 34754 12872 34798 12914
rect 34922 12872 34969 12914
rect 34583 12832 34592 12872
rect 34754 12832 34756 12872
rect 34796 12832 34798 12872
rect 34960 12832 34969 12872
rect 34583 12790 34630 12832
rect 34754 12790 34798 12832
rect 34922 12790 34969 12832
rect 49703 12872 49750 12914
rect 49874 12872 49918 12914
rect 50042 12872 50089 12914
rect 49703 12832 49712 12872
rect 49874 12832 49876 12872
rect 49916 12832 49918 12872
rect 50080 12832 50089 12872
rect 49703 12790 49750 12832
rect 49874 12790 49918 12832
rect 50042 12790 50089 12832
rect 64823 12872 64870 12914
rect 64994 12872 65038 12914
rect 65162 12872 65209 12914
rect 64823 12832 64832 12872
rect 64994 12832 64996 12872
rect 65036 12832 65038 12872
rect 65200 12832 65209 12872
rect 64823 12790 64870 12832
rect 64994 12790 65038 12832
rect 65162 12790 65209 12832
rect 79943 12872 79990 12914
rect 80114 12872 80158 12914
rect 80282 12872 80329 12914
rect 79943 12832 79952 12872
rect 80114 12832 80116 12872
rect 80156 12832 80158 12872
rect 80320 12832 80329 12872
rect 79943 12790 79990 12832
rect 80114 12790 80158 12832
rect 80282 12790 80329 12832
rect 95063 12872 95110 12914
rect 95234 12872 95278 12914
rect 95402 12872 95449 12914
rect 95063 12832 95072 12872
rect 95234 12832 95236 12872
rect 95276 12832 95278 12872
rect 95440 12832 95449 12872
rect 95063 12790 95110 12832
rect 95234 12790 95278 12832
rect 95402 12790 95449 12832
rect 3103 12116 3150 12158
rect 3274 12116 3318 12158
rect 3442 12116 3489 12158
rect 3103 12076 3112 12116
rect 3274 12076 3276 12116
rect 3316 12076 3318 12116
rect 3480 12076 3489 12116
rect 3103 12034 3150 12076
rect 3274 12034 3318 12076
rect 3442 12034 3489 12076
rect 18223 12116 18270 12158
rect 18394 12116 18438 12158
rect 18562 12116 18609 12158
rect 18223 12076 18232 12116
rect 18394 12076 18396 12116
rect 18436 12076 18438 12116
rect 18600 12076 18609 12116
rect 18223 12034 18270 12076
rect 18394 12034 18438 12076
rect 18562 12034 18609 12076
rect 33343 12116 33390 12158
rect 33514 12116 33558 12158
rect 33682 12116 33729 12158
rect 33343 12076 33352 12116
rect 33514 12076 33516 12116
rect 33556 12076 33558 12116
rect 33720 12076 33729 12116
rect 33343 12034 33390 12076
rect 33514 12034 33558 12076
rect 33682 12034 33729 12076
rect 48463 12116 48510 12158
rect 48634 12116 48678 12158
rect 48802 12116 48849 12158
rect 48463 12076 48472 12116
rect 48634 12076 48636 12116
rect 48676 12076 48678 12116
rect 48840 12076 48849 12116
rect 48463 12034 48510 12076
rect 48634 12034 48678 12076
rect 48802 12034 48849 12076
rect 63583 12116 63630 12158
rect 63754 12116 63798 12158
rect 63922 12116 63969 12158
rect 63583 12076 63592 12116
rect 63754 12076 63756 12116
rect 63796 12076 63798 12116
rect 63960 12076 63969 12116
rect 63583 12034 63630 12076
rect 63754 12034 63798 12076
rect 63922 12034 63969 12076
rect 78703 12116 78750 12158
rect 78874 12116 78918 12158
rect 79042 12116 79089 12158
rect 78703 12076 78712 12116
rect 78874 12076 78876 12116
rect 78916 12076 78918 12116
rect 79080 12076 79089 12116
rect 78703 12034 78750 12076
rect 78874 12034 78918 12076
rect 79042 12034 79089 12076
rect 93823 12116 93870 12158
rect 93994 12116 94038 12158
rect 94162 12116 94209 12158
rect 93823 12076 93832 12116
rect 93994 12076 93996 12116
rect 94036 12076 94038 12116
rect 94200 12076 94209 12116
rect 93823 12034 93870 12076
rect 93994 12034 94038 12076
rect 94162 12034 94209 12076
rect 4343 11360 4390 11402
rect 4514 11360 4558 11402
rect 4682 11360 4729 11402
rect 4343 11320 4352 11360
rect 4514 11320 4516 11360
rect 4556 11320 4558 11360
rect 4720 11320 4729 11360
rect 4343 11278 4390 11320
rect 4514 11278 4558 11320
rect 4682 11278 4729 11320
rect 19463 11360 19510 11402
rect 19634 11360 19678 11402
rect 19802 11360 19849 11402
rect 19463 11320 19472 11360
rect 19634 11320 19636 11360
rect 19676 11320 19678 11360
rect 19840 11320 19849 11360
rect 19463 11278 19510 11320
rect 19634 11278 19678 11320
rect 19802 11278 19849 11320
rect 34583 11360 34630 11402
rect 34754 11360 34798 11402
rect 34922 11360 34969 11402
rect 34583 11320 34592 11360
rect 34754 11320 34756 11360
rect 34796 11320 34798 11360
rect 34960 11320 34969 11360
rect 34583 11278 34630 11320
rect 34754 11278 34798 11320
rect 34922 11278 34969 11320
rect 49703 11360 49750 11402
rect 49874 11360 49918 11402
rect 50042 11360 50089 11402
rect 49703 11320 49712 11360
rect 49874 11320 49876 11360
rect 49916 11320 49918 11360
rect 50080 11320 50089 11360
rect 49703 11278 49750 11320
rect 49874 11278 49918 11320
rect 50042 11278 50089 11320
rect 64823 11360 64870 11402
rect 64994 11360 65038 11402
rect 65162 11360 65209 11402
rect 64823 11320 64832 11360
rect 64994 11320 64996 11360
rect 65036 11320 65038 11360
rect 65200 11320 65209 11360
rect 64823 11278 64870 11320
rect 64994 11278 65038 11320
rect 65162 11278 65209 11320
rect 79943 11360 79990 11402
rect 80114 11360 80158 11402
rect 80282 11360 80329 11402
rect 79943 11320 79952 11360
rect 80114 11320 80116 11360
rect 80156 11320 80158 11360
rect 80320 11320 80329 11360
rect 79943 11278 79990 11320
rect 80114 11278 80158 11320
rect 80282 11278 80329 11320
rect 95063 11360 95110 11402
rect 95234 11360 95278 11402
rect 95402 11360 95449 11402
rect 95063 11320 95072 11360
rect 95234 11320 95236 11360
rect 95276 11320 95278 11360
rect 95440 11320 95449 11360
rect 95063 11278 95110 11320
rect 95234 11278 95278 11320
rect 95402 11278 95449 11320
rect 3103 10604 3150 10646
rect 3274 10604 3318 10646
rect 3442 10604 3489 10646
rect 3103 10564 3112 10604
rect 3274 10564 3276 10604
rect 3316 10564 3318 10604
rect 3480 10564 3489 10604
rect 3103 10522 3150 10564
rect 3274 10522 3318 10564
rect 3442 10522 3489 10564
rect 18223 10604 18270 10646
rect 18394 10604 18438 10646
rect 18562 10604 18609 10646
rect 18223 10564 18232 10604
rect 18394 10564 18396 10604
rect 18436 10564 18438 10604
rect 18600 10564 18609 10604
rect 18223 10522 18270 10564
rect 18394 10522 18438 10564
rect 18562 10522 18609 10564
rect 33343 10604 33390 10646
rect 33514 10604 33558 10646
rect 33682 10604 33729 10646
rect 33343 10564 33352 10604
rect 33514 10564 33516 10604
rect 33556 10564 33558 10604
rect 33720 10564 33729 10604
rect 33343 10522 33390 10564
rect 33514 10522 33558 10564
rect 33682 10522 33729 10564
rect 48463 10604 48510 10646
rect 48634 10604 48678 10646
rect 48802 10604 48849 10646
rect 48463 10564 48472 10604
rect 48634 10564 48636 10604
rect 48676 10564 48678 10604
rect 48840 10564 48849 10604
rect 48463 10522 48510 10564
rect 48634 10522 48678 10564
rect 48802 10522 48849 10564
rect 63583 10604 63630 10646
rect 63754 10604 63798 10646
rect 63922 10604 63969 10646
rect 63583 10564 63592 10604
rect 63754 10564 63756 10604
rect 63796 10564 63798 10604
rect 63960 10564 63969 10604
rect 63583 10522 63630 10564
rect 63754 10522 63798 10564
rect 63922 10522 63969 10564
rect 78703 10604 78750 10646
rect 78874 10604 78918 10646
rect 79042 10604 79089 10646
rect 78703 10564 78712 10604
rect 78874 10564 78876 10604
rect 78916 10564 78918 10604
rect 79080 10564 79089 10604
rect 78703 10522 78750 10564
rect 78874 10522 78918 10564
rect 79042 10522 79089 10564
rect 93823 10604 93870 10646
rect 93994 10604 94038 10646
rect 94162 10604 94209 10646
rect 93823 10564 93832 10604
rect 93994 10564 93996 10604
rect 94036 10564 94038 10604
rect 94200 10564 94209 10604
rect 93823 10522 93870 10564
rect 93994 10522 94038 10564
rect 94162 10522 94209 10564
rect 4343 9848 4390 9890
rect 4514 9848 4558 9890
rect 4682 9848 4729 9890
rect 4343 9808 4352 9848
rect 4514 9808 4516 9848
rect 4556 9808 4558 9848
rect 4720 9808 4729 9848
rect 4343 9766 4390 9808
rect 4514 9766 4558 9808
rect 4682 9766 4729 9808
rect 19463 9848 19510 9890
rect 19634 9848 19678 9890
rect 19802 9848 19849 9890
rect 19463 9808 19472 9848
rect 19634 9808 19636 9848
rect 19676 9808 19678 9848
rect 19840 9808 19849 9848
rect 19463 9766 19510 9808
rect 19634 9766 19678 9808
rect 19802 9766 19849 9808
rect 34583 9848 34630 9890
rect 34754 9848 34798 9890
rect 34922 9848 34969 9890
rect 34583 9808 34592 9848
rect 34754 9808 34756 9848
rect 34796 9808 34798 9848
rect 34960 9808 34969 9848
rect 34583 9766 34630 9808
rect 34754 9766 34798 9808
rect 34922 9766 34969 9808
rect 49703 9848 49750 9890
rect 49874 9848 49918 9890
rect 50042 9848 50089 9890
rect 49703 9808 49712 9848
rect 49874 9808 49876 9848
rect 49916 9808 49918 9848
rect 50080 9808 50089 9848
rect 49703 9766 49750 9808
rect 49874 9766 49918 9808
rect 50042 9766 50089 9808
rect 64823 9848 64870 9890
rect 64994 9848 65038 9890
rect 65162 9848 65209 9890
rect 64823 9808 64832 9848
rect 64994 9808 64996 9848
rect 65036 9808 65038 9848
rect 65200 9808 65209 9848
rect 64823 9766 64870 9808
rect 64994 9766 65038 9808
rect 65162 9766 65209 9808
rect 79943 9848 79990 9890
rect 80114 9848 80158 9890
rect 80282 9848 80329 9890
rect 79943 9808 79952 9848
rect 80114 9808 80116 9848
rect 80156 9808 80158 9848
rect 80320 9808 80329 9848
rect 79943 9766 79990 9808
rect 80114 9766 80158 9808
rect 80282 9766 80329 9808
rect 95063 9848 95110 9890
rect 95234 9848 95278 9890
rect 95402 9848 95449 9890
rect 95063 9808 95072 9848
rect 95234 9808 95236 9848
rect 95276 9808 95278 9848
rect 95440 9808 95449 9848
rect 95063 9766 95110 9808
rect 95234 9766 95278 9808
rect 95402 9766 95449 9808
rect 3103 9092 3150 9134
rect 3274 9092 3318 9134
rect 3442 9092 3489 9134
rect 3103 9052 3112 9092
rect 3274 9052 3276 9092
rect 3316 9052 3318 9092
rect 3480 9052 3489 9092
rect 3103 9010 3150 9052
rect 3274 9010 3318 9052
rect 3442 9010 3489 9052
rect 18223 9092 18270 9134
rect 18394 9092 18438 9134
rect 18562 9092 18609 9134
rect 18223 9052 18232 9092
rect 18394 9052 18396 9092
rect 18436 9052 18438 9092
rect 18600 9052 18609 9092
rect 18223 9010 18270 9052
rect 18394 9010 18438 9052
rect 18562 9010 18609 9052
rect 33343 9092 33390 9134
rect 33514 9092 33558 9134
rect 33682 9092 33729 9134
rect 33343 9052 33352 9092
rect 33514 9052 33516 9092
rect 33556 9052 33558 9092
rect 33720 9052 33729 9092
rect 33343 9010 33390 9052
rect 33514 9010 33558 9052
rect 33682 9010 33729 9052
rect 48463 9092 48510 9134
rect 48634 9092 48678 9134
rect 48802 9092 48849 9134
rect 48463 9052 48472 9092
rect 48634 9052 48636 9092
rect 48676 9052 48678 9092
rect 48840 9052 48849 9092
rect 48463 9010 48510 9052
rect 48634 9010 48678 9052
rect 48802 9010 48849 9052
rect 63583 9092 63630 9134
rect 63754 9092 63798 9134
rect 63922 9092 63969 9134
rect 63583 9052 63592 9092
rect 63754 9052 63756 9092
rect 63796 9052 63798 9092
rect 63960 9052 63969 9092
rect 63583 9010 63630 9052
rect 63754 9010 63798 9052
rect 63922 9010 63969 9052
rect 78703 9092 78750 9134
rect 78874 9092 78918 9134
rect 79042 9092 79089 9134
rect 78703 9052 78712 9092
rect 78874 9052 78876 9092
rect 78916 9052 78918 9092
rect 79080 9052 79089 9092
rect 78703 9010 78750 9052
rect 78874 9010 78918 9052
rect 79042 9010 79089 9052
rect 93823 9092 93870 9134
rect 93994 9092 94038 9134
rect 94162 9092 94209 9134
rect 93823 9052 93832 9092
rect 93994 9052 93996 9092
rect 94036 9052 94038 9092
rect 94200 9052 94209 9092
rect 93823 9010 93870 9052
rect 93994 9010 94038 9052
rect 94162 9010 94209 9052
rect 4343 8336 4390 8378
rect 4514 8336 4558 8378
rect 4682 8336 4729 8378
rect 4343 8296 4352 8336
rect 4514 8296 4516 8336
rect 4556 8296 4558 8336
rect 4720 8296 4729 8336
rect 4343 8254 4390 8296
rect 4514 8254 4558 8296
rect 4682 8254 4729 8296
rect 19463 8336 19510 8378
rect 19634 8336 19678 8378
rect 19802 8336 19849 8378
rect 19463 8296 19472 8336
rect 19634 8296 19636 8336
rect 19676 8296 19678 8336
rect 19840 8296 19849 8336
rect 19463 8254 19510 8296
rect 19634 8254 19678 8296
rect 19802 8254 19849 8296
rect 34583 8336 34630 8378
rect 34754 8336 34798 8378
rect 34922 8336 34969 8378
rect 34583 8296 34592 8336
rect 34754 8296 34756 8336
rect 34796 8296 34798 8336
rect 34960 8296 34969 8336
rect 34583 8254 34630 8296
rect 34754 8254 34798 8296
rect 34922 8254 34969 8296
rect 49703 8336 49750 8378
rect 49874 8336 49918 8378
rect 50042 8336 50089 8378
rect 49703 8296 49712 8336
rect 49874 8296 49876 8336
rect 49916 8296 49918 8336
rect 50080 8296 50089 8336
rect 49703 8254 49750 8296
rect 49874 8254 49918 8296
rect 50042 8254 50089 8296
rect 64823 8336 64870 8378
rect 64994 8336 65038 8378
rect 65162 8336 65209 8378
rect 64823 8296 64832 8336
rect 64994 8296 64996 8336
rect 65036 8296 65038 8336
rect 65200 8296 65209 8336
rect 64823 8254 64870 8296
rect 64994 8254 65038 8296
rect 65162 8254 65209 8296
rect 79943 8336 79990 8378
rect 80114 8336 80158 8378
rect 80282 8336 80329 8378
rect 79943 8296 79952 8336
rect 80114 8296 80116 8336
rect 80156 8296 80158 8336
rect 80320 8296 80329 8336
rect 79943 8254 79990 8296
rect 80114 8254 80158 8296
rect 80282 8254 80329 8296
rect 95063 8336 95110 8378
rect 95234 8336 95278 8378
rect 95402 8336 95449 8378
rect 95063 8296 95072 8336
rect 95234 8296 95236 8336
rect 95276 8296 95278 8336
rect 95440 8296 95449 8336
rect 95063 8254 95110 8296
rect 95234 8254 95278 8296
rect 95402 8254 95449 8296
rect 3103 7580 3150 7622
rect 3274 7580 3318 7622
rect 3442 7580 3489 7622
rect 3103 7540 3112 7580
rect 3274 7540 3276 7580
rect 3316 7540 3318 7580
rect 3480 7540 3489 7580
rect 3103 7498 3150 7540
rect 3274 7498 3318 7540
rect 3442 7498 3489 7540
rect 18223 7580 18270 7622
rect 18394 7580 18438 7622
rect 18562 7580 18609 7622
rect 18223 7540 18232 7580
rect 18394 7540 18396 7580
rect 18436 7540 18438 7580
rect 18600 7540 18609 7580
rect 18223 7498 18270 7540
rect 18394 7498 18438 7540
rect 18562 7498 18609 7540
rect 33343 7580 33390 7622
rect 33514 7580 33558 7622
rect 33682 7580 33729 7622
rect 33343 7540 33352 7580
rect 33514 7540 33516 7580
rect 33556 7540 33558 7580
rect 33720 7540 33729 7580
rect 33343 7498 33390 7540
rect 33514 7498 33558 7540
rect 33682 7498 33729 7540
rect 48463 7580 48510 7622
rect 48634 7580 48678 7622
rect 48802 7580 48849 7622
rect 48463 7540 48472 7580
rect 48634 7540 48636 7580
rect 48676 7540 48678 7580
rect 48840 7540 48849 7580
rect 48463 7498 48510 7540
rect 48634 7498 48678 7540
rect 48802 7498 48849 7540
rect 63583 7580 63630 7622
rect 63754 7580 63798 7622
rect 63922 7580 63969 7622
rect 63583 7540 63592 7580
rect 63754 7540 63756 7580
rect 63796 7540 63798 7580
rect 63960 7540 63969 7580
rect 63583 7498 63630 7540
rect 63754 7498 63798 7540
rect 63922 7498 63969 7540
rect 78703 7580 78750 7622
rect 78874 7580 78918 7622
rect 79042 7580 79089 7622
rect 78703 7540 78712 7580
rect 78874 7540 78876 7580
rect 78916 7540 78918 7580
rect 79080 7540 79089 7580
rect 78703 7498 78750 7540
rect 78874 7498 78918 7540
rect 79042 7498 79089 7540
rect 93823 7580 93870 7622
rect 93994 7580 94038 7622
rect 94162 7580 94209 7622
rect 93823 7540 93832 7580
rect 93994 7540 93996 7580
rect 94036 7540 94038 7580
rect 94200 7540 94209 7580
rect 93823 7498 93870 7540
rect 93994 7498 94038 7540
rect 94162 7498 94209 7540
rect 4343 6824 4390 6866
rect 4514 6824 4558 6866
rect 4682 6824 4729 6866
rect 4343 6784 4352 6824
rect 4514 6784 4516 6824
rect 4556 6784 4558 6824
rect 4720 6784 4729 6824
rect 4343 6742 4390 6784
rect 4514 6742 4558 6784
rect 4682 6742 4729 6784
rect 19463 6824 19510 6866
rect 19634 6824 19678 6866
rect 19802 6824 19849 6866
rect 19463 6784 19472 6824
rect 19634 6784 19636 6824
rect 19676 6784 19678 6824
rect 19840 6784 19849 6824
rect 19463 6742 19510 6784
rect 19634 6742 19678 6784
rect 19802 6742 19849 6784
rect 34583 6824 34630 6866
rect 34754 6824 34798 6866
rect 34922 6824 34969 6866
rect 34583 6784 34592 6824
rect 34754 6784 34756 6824
rect 34796 6784 34798 6824
rect 34960 6784 34969 6824
rect 34583 6742 34630 6784
rect 34754 6742 34798 6784
rect 34922 6742 34969 6784
rect 49703 6824 49750 6866
rect 49874 6824 49918 6866
rect 50042 6824 50089 6866
rect 49703 6784 49712 6824
rect 49874 6784 49876 6824
rect 49916 6784 49918 6824
rect 50080 6784 50089 6824
rect 49703 6742 49750 6784
rect 49874 6742 49918 6784
rect 50042 6742 50089 6784
rect 64823 6824 64870 6866
rect 64994 6824 65038 6866
rect 65162 6824 65209 6866
rect 64823 6784 64832 6824
rect 64994 6784 64996 6824
rect 65036 6784 65038 6824
rect 65200 6784 65209 6824
rect 64823 6742 64870 6784
rect 64994 6742 65038 6784
rect 65162 6742 65209 6784
rect 79943 6824 79990 6866
rect 80114 6824 80158 6866
rect 80282 6824 80329 6866
rect 79943 6784 79952 6824
rect 80114 6784 80116 6824
rect 80156 6784 80158 6824
rect 80320 6784 80329 6824
rect 79943 6742 79990 6784
rect 80114 6742 80158 6784
rect 80282 6742 80329 6784
rect 95063 6824 95110 6866
rect 95234 6824 95278 6866
rect 95402 6824 95449 6866
rect 95063 6784 95072 6824
rect 95234 6784 95236 6824
rect 95276 6784 95278 6824
rect 95440 6784 95449 6824
rect 95063 6742 95110 6784
rect 95234 6742 95278 6784
rect 95402 6742 95449 6784
rect 3103 6068 3150 6110
rect 3274 6068 3318 6110
rect 3442 6068 3489 6110
rect 3103 6028 3112 6068
rect 3274 6028 3276 6068
rect 3316 6028 3318 6068
rect 3480 6028 3489 6068
rect 3103 5986 3150 6028
rect 3274 5986 3318 6028
rect 3442 5986 3489 6028
rect 18223 6068 18270 6110
rect 18394 6068 18438 6110
rect 18562 6068 18609 6110
rect 18223 6028 18232 6068
rect 18394 6028 18396 6068
rect 18436 6028 18438 6068
rect 18600 6028 18609 6068
rect 18223 5986 18270 6028
rect 18394 5986 18438 6028
rect 18562 5986 18609 6028
rect 33343 6068 33390 6110
rect 33514 6068 33558 6110
rect 33682 6068 33729 6110
rect 33343 6028 33352 6068
rect 33514 6028 33516 6068
rect 33556 6028 33558 6068
rect 33720 6028 33729 6068
rect 33343 5986 33390 6028
rect 33514 5986 33558 6028
rect 33682 5986 33729 6028
rect 48463 6068 48510 6110
rect 48634 6068 48678 6110
rect 48802 6068 48849 6110
rect 48463 6028 48472 6068
rect 48634 6028 48636 6068
rect 48676 6028 48678 6068
rect 48840 6028 48849 6068
rect 48463 5986 48510 6028
rect 48634 5986 48678 6028
rect 48802 5986 48849 6028
rect 63583 6068 63630 6110
rect 63754 6068 63798 6110
rect 63922 6068 63969 6110
rect 63583 6028 63592 6068
rect 63754 6028 63756 6068
rect 63796 6028 63798 6068
rect 63960 6028 63969 6068
rect 63583 5986 63630 6028
rect 63754 5986 63798 6028
rect 63922 5986 63969 6028
rect 78703 6068 78750 6110
rect 78874 6068 78918 6110
rect 79042 6068 79089 6110
rect 78703 6028 78712 6068
rect 78874 6028 78876 6068
rect 78916 6028 78918 6068
rect 79080 6028 79089 6068
rect 78703 5986 78750 6028
rect 78874 5986 78918 6028
rect 79042 5986 79089 6028
rect 93823 6068 93870 6110
rect 93994 6068 94038 6110
rect 94162 6068 94209 6110
rect 93823 6028 93832 6068
rect 93994 6028 93996 6068
rect 94036 6028 94038 6068
rect 94200 6028 94209 6068
rect 93823 5986 93870 6028
rect 93994 5986 94038 6028
rect 94162 5986 94209 6028
rect 4343 5312 4390 5354
rect 4514 5312 4558 5354
rect 4682 5312 4729 5354
rect 4343 5272 4352 5312
rect 4514 5272 4516 5312
rect 4556 5272 4558 5312
rect 4720 5272 4729 5312
rect 4343 5230 4390 5272
rect 4514 5230 4558 5272
rect 4682 5230 4729 5272
rect 19463 5312 19510 5354
rect 19634 5312 19678 5354
rect 19802 5312 19849 5354
rect 19463 5272 19472 5312
rect 19634 5272 19636 5312
rect 19676 5272 19678 5312
rect 19840 5272 19849 5312
rect 19463 5230 19510 5272
rect 19634 5230 19678 5272
rect 19802 5230 19849 5272
rect 34583 5312 34630 5354
rect 34754 5312 34798 5354
rect 34922 5312 34969 5354
rect 34583 5272 34592 5312
rect 34754 5272 34756 5312
rect 34796 5272 34798 5312
rect 34960 5272 34969 5312
rect 34583 5230 34630 5272
rect 34754 5230 34798 5272
rect 34922 5230 34969 5272
rect 49703 5312 49750 5354
rect 49874 5312 49918 5354
rect 50042 5312 50089 5354
rect 49703 5272 49712 5312
rect 49874 5272 49876 5312
rect 49916 5272 49918 5312
rect 50080 5272 50089 5312
rect 49703 5230 49750 5272
rect 49874 5230 49918 5272
rect 50042 5230 50089 5272
rect 64823 5312 64870 5354
rect 64994 5312 65038 5354
rect 65162 5312 65209 5354
rect 64823 5272 64832 5312
rect 64994 5272 64996 5312
rect 65036 5272 65038 5312
rect 65200 5272 65209 5312
rect 64823 5230 64870 5272
rect 64994 5230 65038 5272
rect 65162 5230 65209 5272
rect 79943 5312 79990 5354
rect 80114 5312 80158 5354
rect 80282 5312 80329 5354
rect 79943 5272 79952 5312
rect 80114 5272 80116 5312
rect 80156 5272 80158 5312
rect 80320 5272 80329 5312
rect 79943 5230 79990 5272
rect 80114 5230 80158 5272
rect 80282 5230 80329 5272
rect 95063 5312 95110 5354
rect 95234 5312 95278 5354
rect 95402 5312 95449 5354
rect 95063 5272 95072 5312
rect 95234 5272 95236 5312
rect 95276 5272 95278 5312
rect 95440 5272 95449 5312
rect 95063 5230 95110 5272
rect 95234 5230 95278 5272
rect 95402 5230 95449 5272
rect 3103 4556 3150 4598
rect 3274 4556 3318 4598
rect 3442 4556 3489 4598
rect 3103 4516 3112 4556
rect 3274 4516 3276 4556
rect 3316 4516 3318 4556
rect 3480 4516 3489 4556
rect 3103 4474 3150 4516
rect 3274 4474 3318 4516
rect 3442 4474 3489 4516
rect 18223 4556 18270 4598
rect 18394 4556 18438 4598
rect 18562 4556 18609 4598
rect 18223 4516 18232 4556
rect 18394 4516 18396 4556
rect 18436 4516 18438 4556
rect 18600 4516 18609 4556
rect 18223 4474 18270 4516
rect 18394 4474 18438 4516
rect 18562 4474 18609 4516
rect 33343 4556 33390 4598
rect 33514 4556 33558 4598
rect 33682 4556 33729 4598
rect 33343 4516 33352 4556
rect 33514 4516 33516 4556
rect 33556 4516 33558 4556
rect 33720 4516 33729 4556
rect 33343 4474 33390 4516
rect 33514 4474 33558 4516
rect 33682 4474 33729 4516
rect 48463 4556 48510 4598
rect 48634 4556 48678 4598
rect 48802 4556 48849 4598
rect 48463 4516 48472 4556
rect 48634 4516 48636 4556
rect 48676 4516 48678 4556
rect 48840 4516 48849 4556
rect 48463 4474 48510 4516
rect 48634 4474 48678 4516
rect 48802 4474 48849 4516
rect 63583 4556 63630 4598
rect 63754 4556 63798 4598
rect 63922 4556 63969 4598
rect 63583 4516 63592 4556
rect 63754 4516 63756 4556
rect 63796 4516 63798 4556
rect 63960 4516 63969 4556
rect 63583 4474 63630 4516
rect 63754 4474 63798 4516
rect 63922 4474 63969 4516
rect 78703 4556 78750 4598
rect 78874 4556 78918 4598
rect 79042 4556 79089 4598
rect 78703 4516 78712 4556
rect 78874 4516 78876 4556
rect 78916 4516 78918 4556
rect 79080 4516 79089 4556
rect 78703 4474 78750 4516
rect 78874 4474 78918 4516
rect 79042 4474 79089 4516
rect 93823 4556 93870 4598
rect 93994 4556 94038 4598
rect 94162 4556 94209 4598
rect 93823 4516 93832 4556
rect 93994 4516 93996 4556
rect 94036 4516 94038 4556
rect 94200 4516 94209 4556
rect 93823 4474 93870 4516
rect 93994 4474 94038 4516
rect 94162 4474 94209 4516
rect 4343 3800 4390 3842
rect 4514 3800 4558 3842
rect 4682 3800 4729 3842
rect 4343 3760 4352 3800
rect 4514 3760 4516 3800
rect 4556 3760 4558 3800
rect 4720 3760 4729 3800
rect 4343 3718 4390 3760
rect 4514 3718 4558 3760
rect 4682 3718 4729 3760
rect 19463 3800 19510 3842
rect 19634 3800 19678 3842
rect 19802 3800 19849 3842
rect 19463 3760 19472 3800
rect 19634 3760 19636 3800
rect 19676 3760 19678 3800
rect 19840 3760 19849 3800
rect 19463 3718 19510 3760
rect 19634 3718 19678 3760
rect 19802 3718 19849 3760
rect 34583 3800 34630 3842
rect 34754 3800 34798 3842
rect 34922 3800 34969 3842
rect 34583 3760 34592 3800
rect 34754 3760 34756 3800
rect 34796 3760 34798 3800
rect 34960 3760 34969 3800
rect 34583 3718 34630 3760
rect 34754 3718 34798 3760
rect 34922 3718 34969 3760
rect 49703 3800 49750 3842
rect 49874 3800 49918 3842
rect 50042 3800 50089 3842
rect 49703 3760 49712 3800
rect 49874 3760 49876 3800
rect 49916 3760 49918 3800
rect 50080 3760 50089 3800
rect 49703 3718 49750 3760
rect 49874 3718 49918 3760
rect 50042 3718 50089 3760
rect 64823 3800 64870 3842
rect 64994 3800 65038 3842
rect 65162 3800 65209 3842
rect 64823 3760 64832 3800
rect 64994 3760 64996 3800
rect 65036 3760 65038 3800
rect 65200 3760 65209 3800
rect 64823 3718 64870 3760
rect 64994 3718 65038 3760
rect 65162 3718 65209 3760
rect 79943 3800 79990 3842
rect 80114 3800 80158 3842
rect 80282 3800 80329 3842
rect 79943 3760 79952 3800
rect 80114 3760 80116 3800
rect 80156 3760 80158 3800
rect 80320 3760 80329 3800
rect 79943 3718 79990 3760
rect 80114 3718 80158 3760
rect 80282 3718 80329 3760
rect 95063 3800 95110 3842
rect 95234 3800 95278 3842
rect 95402 3800 95449 3842
rect 95063 3760 95072 3800
rect 95234 3760 95236 3800
rect 95276 3760 95278 3800
rect 95440 3760 95449 3800
rect 95063 3718 95110 3760
rect 95234 3718 95278 3760
rect 95402 3718 95449 3760
rect 3103 3044 3150 3086
rect 3274 3044 3318 3086
rect 3442 3044 3489 3086
rect 3103 3004 3112 3044
rect 3274 3004 3276 3044
rect 3316 3004 3318 3044
rect 3480 3004 3489 3044
rect 3103 2962 3150 3004
rect 3274 2962 3318 3004
rect 3442 2962 3489 3004
rect 18223 3044 18270 3086
rect 18394 3044 18438 3086
rect 18562 3044 18609 3086
rect 18223 3004 18232 3044
rect 18394 3004 18396 3044
rect 18436 3004 18438 3044
rect 18600 3004 18609 3044
rect 18223 2962 18270 3004
rect 18394 2962 18438 3004
rect 18562 2962 18609 3004
rect 33343 3044 33390 3086
rect 33514 3044 33558 3086
rect 33682 3044 33729 3086
rect 33343 3004 33352 3044
rect 33514 3004 33516 3044
rect 33556 3004 33558 3044
rect 33720 3004 33729 3044
rect 33343 2962 33390 3004
rect 33514 2962 33558 3004
rect 33682 2962 33729 3004
rect 48463 3044 48510 3086
rect 48634 3044 48678 3086
rect 48802 3044 48849 3086
rect 48463 3004 48472 3044
rect 48634 3004 48636 3044
rect 48676 3004 48678 3044
rect 48840 3004 48849 3044
rect 48463 2962 48510 3004
rect 48634 2962 48678 3004
rect 48802 2962 48849 3004
rect 63583 3044 63630 3086
rect 63754 3044 63798 3086
rect 63922 3044 63969 3086
rect 63583 3004 63592 3044
rect 63754 3004 63756 3044
rect 63796 3004 63798 3044
rect 63960 3004 63969 3044
rect 63583 2962 63630 3004
rect 63754 2962 63798 3004
rect 63922 2962 63969 3004
rect 78703 3044 78750 3086
rect 78874 3044 78918 3086
rect 79042 3044 79089 3086
rect 78703 3004 78712 3044
rect 78874 3004 78876 3044
rect 78916 3004 78918 3044
rect 79080 3004 79089 3044
rect 78703 2962 78750 3004
rect 78874 2962 78918 3004
rect 79042 2962 79089 3004
rect 93823 3044 93870 3086
rect 93994 3044 94038 3086
rect 94162 3044 94209 3086
rect 93823 3004 93832 3044
rect 93994 3004 93996 3044
rect 94036 3004 94038 3044
rect 94200 3004 94209 3044
rect 93823 2962 93870 3004
rect 93994 2962 94038 3004
rect 94162 2962 94209 3004
rect 4343 2288 4390 2330
rect 4514 2288 4558 2330
rect 4682 2288 4729 2330
rect 4343 2248 4352 2288
rect 4514 2248 4516 2288
rect 4556 2248 4558 2288
rect 4720 2248 4729 2288
rect 4343 2206 4390 2248
rect 4514 2206 4558 2248
rect 4682 2206 4729 2248
rect 19463 2288 19510 2330
rect 19634 2288 19678 2330
rect 19802 2288 19849 2330
rect 19463 2248 19472 2288
rect 19634 2248 19636 2288
rect 19676 2248 19678 2288
rect 19840 2248 19849 2288
rect 19463 2206 19510 2248
rect 19634 2206 19678 2248
rect 19802 2206 19849 2248
rect 34583 2288 34630 2330
rect 34754 2288 34798 2330
rect 34922 2288 34969 2330
rect 34583 2248 34592 2288
rect 34754 2248 34756 2288
rect 34796 2248 34798 2288
rect 34960 2248 34969 2288
rect 34583 2206 34630 2248
rect 34754 2206 34798 2248
rect 34922 2206 34969 2248
rect 49703 2288 49750 2330
rect 49874 2288 49918 2330
rect 50042 2288 50089 2330
rect 49703 2248 49712 2288
rect 49874 2248 49876 2288
rect 49916 2248 49918 2288
rect 50080 2248 50089 2288
rect 49703 2206 49750 2248
rect 49874 2206 49918 2248
rect 50042 2206 50089 2248
rect 64823 2288 64870 2330
rect 64994 2288 65038 2330
rect 65162 2288 65209 2330
rect 64823 2248 64832 2288
rect 64994 2248 64996 2288
rect 65036 2248 65038 2288
rect 65200 2248 65209 2288
rect 64823 2206 64870 2248
rect 64994 2206 65038 2248
rect 65162 2206 65209 2248
rect 79943 2288 79990 2330
rect 80114 2288 80158 2330
rect 80282 2288 80329 2330
rect 79943 2248 79952 2288
rect 80114 2248 80116 2288
rect 80156 2248 80158 2288
rect 80320 2248 80329 2288
rect 79943 2206 79990 2248
rect 80114 2206 80158 2248
rect 80282 2206 80329 2248
rect 95063 2288 95110 2330
rect 95234 2288 95278 2330
rect 95402 2288 95449 2330
rect 95063 2248 95072 2288
rect 95234 2248 95236 2288
rect 95276 2248 95278 2288
rect 95440 2248 95449 2288
rect 95063 2206 95110 2248
rect 95234 2206 95278 2248
rect 95402 2206 95449 2248
rect 3103 1532 3150 1574
rect 3274 1532 3318 1574
rect 3442 1532 3489 1574
rect 3103 1492 3112 1532
rect 3274 1492 3276 1532
rect 3316 1492 3318 1532
rect 3480 1492 3489 1532
rect 3103 1450 3150 1492
rect 3274 1450 3318 1492
rect 3442 1450 3489 1492
rect 18223 1532 18270 1574
rect 18394 1532 18438 1574
rect 18562 1532 18609 1574
rect 18223 1492 18232 1532
rect 18394 1492 18396 1532
rect 18436 1492 18438 1532
rect 18600 1492 18609 1532
rect 18223 1450 18270 1492
rect 18394 1450 18438 1492
rect 18562 1450 18609 1492
rect 33343 1532 33390 1574
rect 33514 1532 33558 1574
rect 33682 1532 33729 1574
rect 33343 1492 33352 1532
rect 33514 1492 33516 1532
rect 33556 1492 33558 1532
rect 33720 1492 33729 1532
rect 33343 1450 33390 1492
rect 33514 1450 33558 1492
rect 33682 1450 33729 1492
rect 48463 1532 48510 1574
rect 48634 1532 48678 1574
rect 48802 1532 48849 1574
rect 48463 1492 48472 1532
rect 48634 1492 48636 1532
rect 48676 1492 48678 1532
rect 48840 1492 48849 1532
rect 48463 1450 48510 1492
rect 48634 1450 48678 1492
rect 48802 1450 48849 1492
rect 63583 1532 63630 1574
rect 63754 1532 63798 1574
rect 63922 1532 63969 1574
rect 63583 1492 63592 1532
rect 63754 1492 63756 1532
rect 63796 1492 63798 1532
rect 63960 1492 63969 1532
rect 63583 1450 63630 1492
rect 63754 1450 63798 1492
rect 63922 1450 63969 1492
rect 78703 1532 78750 1574
rect 78874 1532 78918 1574
rect 79042 1532 79089 1574
rect 78703 1492 78712 1532
rect 78874 1492 78876 1532
rect 78916 1492 78918 1532
rect 79080 1492 79089 1532
rect 78703 1450 78750 1492
rect 78874 1450 78918 1492
rect 79042 1450 79089 1492
rect 93823 1532 93870 1574
rect 93994 1532 94038 1574
rect 94162 1532 94209 1574
rect 93823 1492 93832 1532
rect 93994 1492 93996 1532
rect 94036 1492 94038 1532
rect 94200 1492 94209 1532
rect 93823 1450 93870 1492
rect 93994 1450 94038 1492
rect 94162 1450 94209 1492
rect 4343 776 4390 818
rect 4514 776 4558 818
rect 4682 776 4729 818
rect 4343 736 4352 776
rect 4514 736 4516 776
rect 4556 736 4558 776
rect 4720 736 4729 776
rect 4343 694 4390 736
rect 4514 694 4558 736
rect 4682 694 4729 736
rect 19463 776 19510 818
rect 19634 776 19678 818
rect 19802 776 19849 818
rect 19463 736 19472 776
rect 19634 736 19636 776
rect 19676 736 19678 776
rect 19840 736 19849 776
rect 19463 694 19510 736
rect 19634 694 19678 736
rect 19802 694 19849 736
rect 34583 776 34630 818
rect 34754 776 34798 818
rect 34922 776 34969 818
rect 34583 736 34592 776
rect 34754 736 34756 776
rect 34796 736 34798 776
rect 34960 736 34969 776
rect 34583 694 34630 736
rect 34754 694 34798 736
rect 34922 694 34969 736
rect 49703 776 49750 818
rect 49874 776 49918 818
rect 50042 776 50089 818
rect 49703 736 49712 776
rect 49874 736 49876 776
rect 49916 736 49918 776
rect 50080 736 50089 776
rect 49703 694 49750 736
rect 49874 694 49918 736
rect 50042 694 50089 736
rect 64823 776 64870 818
rect 64994 776 65038 818
rect 65162 776 65209 818
rect 64823 736 64832 776
rect 64994 736 64996 776
rect 65036 736 65038 776
rect 65200 736 65209 776
rect 64823 694 64870 736
rect 64994 694 65038 736
rect 65162 694 65209 736
rect 79943 776 79990 818
rect 80114 776 80158 818
rect 80282 776 80329 818
rect 79943 736 79952 776
rect 80114 736 80116 776
rect 80156 736 80158 776
rect 80320 736 80329 776
rect 79943 694 79990 736
rect 80114 694 80158 736
rect 80282 694 80329 736
rect 95063 776 95110 818
rect 95234 776 95278 818
rect 95402 776 95449 818
rect 95063 736 95072 776
rect 95234 736 95236 776
rect 95276 736 95278 776
rect 95440 736 95449 776
rect 95063 694 95110 736
rect 95234 694 95278 736
rect 95402 694 95449 736
<< via5 >>
rect 4390 38576 4514 38618
rect 4558 38576 4682 38618
rect 4390 38536 4392 38576
rect 4392 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4514 38576
rect 4558 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4680 38576
rect 4680 38536 4682 38576
rect 4390 38494 4514 38536
rect 4558 38494 4682 38536
rect 19510 38576 19634 38618
rect 19678 38576 19802 38618
rect 19510 38536 19512 38576
rect 19512 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19634 38576
rect 19678 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19800 38576
rect 19800 38536 19802 38576
rect 19510 38494 19634 38536
rect 19678 38494 19802 38536
rect 34630 38576 34754 38618
rect 34798 38576 34922 38618
rect 34630 38536 34632 38576
rect 34632 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34754 38576
rect 34798 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34920 38576
rect 34920 38536 34922 38576
rect 34630 38494 34754 38536
rect 34798 38494 34922 38536
rect 49750 38576 49874 38618
rect 49918 38576 50042 38618
rect 49750 38536 49752 38576
rect 49752 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49874 38576
rect 49918 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50040 38576
rect 50040 38536 50042 38576
rect 49750 38494 49874 38536
rect 49918 38494 50042 38536
rect 64870 38576 64994 38618
rect 65038 38576 65162 38618
rect 64870 38536 64872 38576
rect 64872 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64994 38576
rect 65038 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65160 38576
rect 65160 38536 65162 38576
rect 64870 38494 64994 38536
rect 65038 38494 65162 38536
rect 79990 38576 80114 38618
rect 80158 38576 80282 38618
rect 79990 38536 79992 38576
rect 79992 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80114 38576
rect 80158 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80280 38576
rect 80280 38536 80282 38576
rect 79990 38494 80114 38536
rect 80158 38494 80282 38536
rect 95110 38576 95234 38618
rect 95278 38576 95402 38618
rect 95110 38536 95112 38576
rect 95112 38536 95154 38576
rect 95154 38536 95194 38576
rect 95194 38536 95234 38576
rect 95278 38536 95318 38576
rect 95318 38536 95358 38576
rect 95358 38536 95400 38576
rect 95400 38536 95402 38576
rect 95110 38494 95234 38536
rect 95278 38494 95402 38536
rect 3150 37820 3274 37862
rect 3318 37820 3442 37862
rect 3150 37780 3152 37820
rect 3152 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3274 37820
rect 3318 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3440 37820
rect 3440 37780 3442 37820
rect 3150 37738 3274 37780
rect 3318 37738 3442 37780
rect 18270 37820 18394 37862
rect 18438 37820 18562 37862
rect 18270 37780 18272 37820
rect 18272 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18394 37820
rect 18438 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18560 37820
rect 18560 37780 18562 37820
rect 18270 37738 18394 37780
rect 18438 37738 18562 37780
rect 33390 37820 33514 37862
rect 33558 37820 33682 37862
rect 33390 37780 33392 37820
rect 33392 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33514 37820
rect 33558 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33680 37820
rect 33680 37780 33682 37820
rect 33390 37738 33514 37780
rect 33558 37738 33682 37780
rect 48510 37820 48634 37862
rect 48678 37820 48802 37862
rect 48510 37780 48512 37820
rect 48512 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48634 37820
rect 48678 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48800 37820
rect 48800 37780 48802 37820
rect 48510 37738 48634 37780
rect 48678 37738 48802 37780
rect 63630 37820 63754 37862
rect 63798 37820 63922 37862
rect 63630 37780 63632 37820
rect 63632 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63754 37820
rect 63798 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63920 37820
rect 63920 37780 63922 37820
rect 63630 37738 63754 37780
rect 63798 37738 63922 37780
rect 78750 37820 78874 37862
rect 78918 37820 79042 37862
rect 78750 37780 78752 37820
rect 78752 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78874 37820
rect 78918 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79040 37820
rect 79040 37780 79042 37820
rect 78750 37738 78874 37780
rect 78918 37738 79042 37780
rect 93870 37820 93994 37862
rect 94038 37820 94162 37862
rect 93870 37780 93872 37820
rect 93872 37780 93914 37820
rect 93914 37780 93954 37820
rect 93954 37780 93994 37820
rect 94038 37780 94078 37820
rect 94078 37780 94118 37820
rect 94118 37780 94160 37820
rect 94160 37780 94162 37820
rect 93870 37738 93994 37780
rect 94038 37738 94162 37780
rect 4390 37064 4514 37106
rect 4558 37064 4682 37106
rect 4390 37024 4392 37064
rect 4392 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4514 37064
rect 4558 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4680 37064
rect 4680 37024 4682 37064
rect 4390 36982 4514 37024
rect 4558 36982 4682 37024
rect 19510 37064 19634 37106
rect 19678 37064 19802 37106
rect 19510 37024 19512 37064
rect 19512 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19634 37064
rect 19678 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19800 37064
rect 19800 37024 19802 37064
rect 19510 36982 19634 37024
rect 19678 36982 19802 37024
rect 34630 37064 34754 37106
rect 34798 37064 34922 37106
rect 34630 37024 34632 37064
rect 34632 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34754 37064
rect 34798 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34920 37064
rect 34920 37024 34922 37064
rect 34630 36982 34754 37024
rect 34798 36982 34922 37024
rect 49750 37064 49874 37106
rect 49918 37064 50042 37106
rect 49750 37024 49752 37064
rect 49752 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49874 37064
rect 49918 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50040 37064
rect 50040 37024 50042 37064
rect 49750 36982 49874 37024
rect 49918 36982 50042 37024
rect 64870 37064 64994 37106
rect 65038 37064 65162 37106
rect 64870 37024 64872 37064
rect 64872 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64994 37064
rect 65038 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65160 37064
rect 65160 37024 65162 37064
rect 64870 36982 64994 37024
rect 65038 36982 65162 37024
rect 79990 37064 80114 37106
rect 80158 37064 80282 37106
rect 79990 37024 79992 37064
rect 79992 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80114 37064
rect 80158 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80280 37064
rect 80280 37024 80282 37064
rect 79990 36982 80114 37024
rect 80158 36982 80282 37024
rect 95110 37064 95234 37106
rect 95278 37064 95402 37106
rect 95110 37024 95112 37064
rect 95112 37024 95154 37064
rect 95154 37024 95194 37064
rect 95194 37024 95234 37064
rect 95278 37024 95318 37064
rect 95318 37024 95358 37064
rect 95358 37024 95400 37064
rect 95400 37024 95402 37064
rect 95110 36982 95234 37024
rect 95278 36982 95402 37024
rect 3150 36308 3274 36350
rect 3318 36308 3442 36350
rect 3150 36268 3152 36308
rect 3152 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3274 36308
rect 3318 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3440 36308
rect 3440 36268 3442 36308
rect 3150 36226 3274 36268
rect 3318 36226 3442 36268
rect 18270 36308 18394 36350
rect 18438 36308 18562 36350
rect 18270 36268 18272 36308
rect 18272 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18394 36308
rect 18438 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18560 36308
rect 18560 36268 18562 36308
rect 18270 36226 18394 36268
rect 18438 36226 18562 36268
rect 33390 36308 33514 36350
rect 33558 36308 33682 36350
rect 33390 36268 33392 36308
rect 33392 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33514 36308
rect 33558 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33680 36308
rect 33680 36268 33682 36308
rect 33390 36226 33514 36268
rect 33558 36226 33682 36268
rect 48510 36308 48634 36350
rect 48678 36308 48802 36350
rect 48510 36268 48512 36308
rect 48512 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48634 36308
rect 48678 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48800 36308
rect 48800 36268 48802 36308
rect 48510 36226 48634 36268
rect 48678 36226 48802 36268
rect 63630 36308 63754 36350
rect 63798 36308 63922 36350
rect 63630 36268 63632 36308
rect 63632 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63754 36308
rect 63798 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63920 36308
rect 63920 36268 63922 36308
rect 63630 36226 63754 36268
rect 63798 36226 63922 36268
rect 78750 36308 78874 36350
rect 78918 36308 79042 36350
rect 78750 36268 78752 36308
rect 78752 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78874 36308
rect 78918 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79040 36308
rect 79040 36268 79042 36308
rect 78750 36226 78874 36268
rect 78918 36226 79042 36268
rect 93870 36308 93994 36350
rect 94038 36308 94162 36350
rect 93870 36268 93872 36308
rect 93872 36268 93914 36308
rect 93914 36268 93954 36308
rect 93954 36268 93994 36308
rect 94038 36268 94078 36308
rect 94078 36268 94118 36308
rect 94118 36268 94160 36308
rect 94160 36268 94162 36308
rect 93870 36226 93994 36268
rect 94038 36226 94162 36268
rect 4390 35552 4514 35594
rect 4558 35552 4682 35594
rect 4390 35512 4392 35552
rect 4392 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4514 35552
rect 4558 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4680 35552
rect 4680 35512 4682 35552
rect 4390 35470 4514 35512
rect 4558 35470 4682 35512
rect 19510 35552 19634 35594
rect 19678 35552 19802 35594
rect 19510 35512 19512 35552
rect 19512 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19634 35552
rect 19678 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19800 35552
rect 19800 35512 19802 35552
rect 19510 35470 19634 35512
rect 19678 35470 19802 35512
rect 34630 35552 34754 35594
rect 34798 35552 34922 35594
rect 34630 35512 34632 35552
rect 34632 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34754 35552
rect 34798 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34920 35552
rect 34920 35512 34922 35552
rect 34630 35470 34754 35512
rect 34798 35470 34922 35512
rect 49750 35552 49874 35594
rect 49918 35552 50042 35594
rect 49750 35512 49752 35552
rect 49752 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49874 35552
rect 49918 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50040 35552
rect 50040 35512 50042 35552
rect 49750 35470 49874 35512
rect 49918 35470 50042 35512
rect 64870 35552 64994 35594
rect 65038 35552 65162 35594
rect 64870 35512 64872 35552
rect 64872 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64994 35552
rect 65038 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65160 35552
rect 65160 35512 65162 35552
rect 64870 35470 64994 35512
rect 65038 35470 65162 35512
rect 79990 35552 80114 35594
rect 80158 35552 80282 35594
rect 79990 35512 79992 35552
rect 79992 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80114 35552
rect 80158 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80280 35552
rect 80280 35512 80282 35552
rect 79990 35470 80114 35512
rect 80158 35470 80282 35512
rect 95110 35552 95234 35594
rect 95278 35552 95402 35594
rect 95110 35512 95112 35552
rect 95112 35512 95154 35552
rect 95154 35512 95194 35552
rect 95194 35512 95234 35552
rect 95278 35512 95318 35552
rect 95318 35512 95358 35552
rect 95358 35512 95400 35552
rect 95400 35512 95402 35552
rect 95110 35470 95234 35512
rect 95278 35470 95402 35512
rect 3150 34796 3274 34838
rect 3318 34796 3442 34838
rect 3150 34756 3152 34796
rect 3152 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3274 34796
rect 3318 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3440 34796
rect 3440 34756 3442 34796
rect 3150 34714 3274 34756
rect 3318 34714 3442 34756
rect 18270 34796 18394 34838
rect 18438 34796 18562 34838
rect 18270 34756 18272 34796
rect 18272 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18394 34796
rect 18438 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18560 34796
rect 18560 34756 18562 34796
rect 18270 34714 18394 34756
rect 18438 34714 18562 34756
rect 33390 34796 33514 34838
rect 33558 34796 33682 34838
rect 33390 34756 33392 34796
rect 33392 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33514 34796
rect 33558 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33680 34796
rect 33680 34756 33682 34796
rect 33390 34714 33514 34756
rect 33558 34714 33682 34756
rect 48510 34796 48634 34838
rect 48678 34796 48802 34838
rect 48510 34756 48512 34796
rect 48512 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48634 34796
rect 48678 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48800 34796
rect 48800 34756 48802 34796
rect 48510 34714 48634 34756
rect 48678 34714 48802 34756
rect 63630 34796 63754 34838
rect 63798 34796 63922 34838
rect 63630 34756 63632 34796
rect 63632 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63754 34796
rect 63798 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63920 34796
rect 63920 34756 63922 34796
rect 63630 34714 63754 34756
rect 63798 34714 63922 34756
rect 78750 34796 78874 34838
rect 78918 34796 79042 34838
rect 78750 34756 78752 34796
rect 78752 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78874 34796
rect 78918 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79040 34796
rect 79040 34756 79042 34796
rect 78750 34714 78874 34756
rect 78918 34714 79042 34756
rect 93870 34796 93994 34838
rect 94038 34796 94162 34838
rect 93870 34756 93872 34796
rect 93872 34756 93914 34796
rect 93914 34756 93954 34796
rect 93954 34756 93994 34796
rect 94038 34756 94078 34796
rect 94078 34756 94118 34796
rect 94118 34756 94160 34796
rect 94160 34756 94162 34796
rect 93870 34714 93994 34756
rect 94038 34714 94162 34756
rect 4390 34040 4514 34082
rect 4558 34040 4682 34082
rect 4390 34000 4392 34040
rect 4392 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4514 34040
rect 4558 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4680 34040
rect 4680 34000 4682 34040
rect 4390 33958 4514 34000
rect 4558 33958 4682 34000
rect 19510 34040 19634 34082
rect 19678 34040 19802 34082
rect 19510 34000 19512 34040
rect 19512 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19634 34040
rect 19678 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19800 34040
rect 19800 34000 19802 34040
rect 19510 33958 19634 34000
rect 19678 33958 19802 34000
rect 34630 34040 34754 34082
rect 34798 34040 34922 34082
rect 34630 34000 34632 34040
rect 34632 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34754 34040
rect 34798 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34920 34040
rect 34920 34000 34922 34040
rect 34630 33958 34754 34000
rect 34798 33958 34922 34000
rect 49750 34040 49874 34082
rect 49918 34040 50042 34082
rect 49750 34000 49752 34040
rect 49752 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49874 34040
rect 49918 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50040 34040
rect 50040 34000 50042 34040
rect 49750 33958 49874 34000
rect 49918 33958 50042 34000
rect 64870 34040 64994 34082
rect 65038 34040 65162 34082
rect 64870 34000 64872 34040
rect 64872 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64994 34040
rect 65038 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65160 34040
rect 65160 34000 65162 34040
rect 64870 33958 64994 34000
rect 65038 33958 65162 34000
rect 79990 34040 80114 34082
rect 80158 34040 80282 34082
rect 79990 34000 79992 34040
rect 79992 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80114 34040
rect 80158 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80280 34040
rect 80280 34000 80282 34040
rect 79990 33958 80114 34000
rect 80158 33958 80282 34000
rect 95110 34040 95234 34082
rect 95278 34040 95402 34082
rect 95110 34000 95112 34040
rect 95112 34000 95154 34040
rect 95154 34000 95194 34040
rect 95194 34000 95234 34040
rect 95278 34000 95318 34040
rect 95318 34000 95358 34040
rect 95358 34000 95400 34040
rect 95400 34000 95402 34040
rect 95110 33958 95234 34000
rect 95278 33958 95402 34000
rect 3150 33284 3274 33326
rect 3318 33284 3442 33326
rect 3150 33244 3152 33284
rect 3152 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3274 33284
rect 3318 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3440 33284
rect 3440 33244 3442 33284
rect 3150 33202 3274 33244
rect 3318 33202 3442 33244
rect 18270 33284 18394 33326
rect 18438 33284 18562 33326
rect 18270 33244 18272 33284
rect 18272 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18394 33284
rect 18438 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18560 33284
rect 18560 33244 18562 33284
rect 18270 33202 18394 33244
rect 18438 33202 18562 33244
rect 33390 33284 33514 33326
rect 33558 33284 33682 33326
rect 33390 33244 33392 33284
rect 33392 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33514 33284
rect 33558 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33680 33284
rect 33680 33244 33682 33284
rect 33390 33202 33514 33244
rect 33558 33202 33682 33244
rect 48510 33284 48634 33326
rect 48678 33284 48802 33326
rect 48510 33244 48512 33284
rect 48512 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48634 33284
rect 48678 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48800 33284
rect 48800 33244 48802 33284
rect 48510 33202 48634 33244
rect 48678 33202 48802 33244
rect 63630 33284 63754 33326
rect 63798 33284 63922 33326
rect 63630 33244 63632 33284
rect 63632 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63754 33284
rect 63798 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63920 33284
rect 63920 33244 63922 33284
rect 63630 33202 63754 33244
rect 63798 33202 63922 33244
rect 78750 33284 78874 33326
rect 78918 33284 79042 33326
rect 78750 33244 78752 33284
rect 78752 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78874 33284
rect 78918 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79040 33284
rect 79040 33244 79042 33284
rect 78750 33202 78874 33244
rect 78918 33202 79042 33244
rect 93870 33284 93994 33326
rect 94038 33284 94162 33326
rect 93870 33244 93872 33284
rect 93872 33244 93914 33284
rect 93914 33244 93954 33284
rect 93954 33244 93994 33284
rect 94038 33244 94078 33284
rect 94078 33244 94118 33284
rect 94118 33244 94160 33284
rect 94160 33244 94162 33284
rect 93870 33202 93994 33244
rect 94038 33202 94162 33244
rect 4390 32528 4514 32570
rect 4558 32528 4682 32570
rect 4390 32488 4392 32528
rect 4392 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4514 32528
rect 4558 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4680 32528
rect 4680 32488 4682 32528
rect 4390 32446 4514 32488
rect 4558 32446 4682 32488
rect 19510 32528 19634 32570
rect 19678 32528 19802 32570
rect 19510 32488 19512 32528
rect 19512 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19634 32528
rect 19678 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19800 32528
rect 19800 32488 19802 32528
rect 19510 32446 19634 32488
rect 19678 32446 19802 32488
rect 34630 32528 34754 32570
rect 34798 32528 34922 32570
rect 34630 32488 34632 32528
rect 34632 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34754 32528
rect 34798 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34920 32528
rect 34920 32488 34922 32528
rect 34630 32446 34754 32488
rect 34798 32446 34922 32488
rect 49750 32528 49874 32570
rect 49918 32528 50042 32570
rect 49750 32488 49752 32528
rect 49752 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49874 32528
rect 49918 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50040 32528
rect 50040 32488 50042 32528
rect 49750 32446 49874 32488
rect 49918 32446 50042 32488
rect 64870 32528 64994 32570
rect 65038 32528 65162 32570
rect 64870 32488 64872 32528
rect 64872 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64994 32528
rect 65038 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65160 32528
rect 65160 32488 65162 32528
rect 64870 32446 64994 32488
rect 65038 32446 65162 32488
rect 79990 32528 80114 32570
rect 80158 32528 80282 32570
rect 79990 32488 79992 32528
rect 79992 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80114 32528
rect 80158 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80280 32528
rect 80280 32488 80282 32528
rect 79990 32446 80114 32488
rect 80158 32446 80282 32488
rect 95110 32528 95234 32570
rect 95278 32528 95402 32570
rect 95110 32488 95112 32528
rect 95112 32488 95154 32528
rect 95154 32488 95194 32528
rect 95194 32488 95234 32528
rect 95278 32488 95318 32528
rect 95318 32488 95358 32528
rect 95358 32488 95400 32528
rect 95400 32488 95402 32528
rect 95110 32446 95234 32488
rect 95278 32446 95402 32488
rect 3150 31772 3274 31814
rect 3318 31772 3442 31814
rect 3150 31732 3152 31772
rect 3152 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3274 31772
rect 3318 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3440 31772
rect 3440 31732 3442 31772
rect 3150 31690 3274 31732
rect 3318 31690 3442 31732
rect 18270 31772 18394 31814
rect 18438 31772 18562 31814
rect 18270 31732 18272 31772
rect 18272 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18394 31772
rect 18438 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18560 31772
rect 18560 31732 18562 31772
rect 18270 31690 18394 31732
rect 18438 31690 18562 31732
rect 33390 31772 33514 31814
rect 33558 31772 33682 31814
rect 33390 31732 33392 31772
rect 33392 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33514 31772
rect 33558 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33680 31772
rect 33680 31732 33682 31772
rect 33390 31690 33514 31732
rect 33558 31690 33682 31732
rect 48510 31772 48634 31814
rect 48678 31772 48802 31814
rect 48510 31732 48512 31772
rect 48512 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48634 31772
rect 48678 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48800 31772
rect 48800 31732 48802 31772
rect 48510 31690 48634 31732
rect 48678 31690 48802 31732
rect 63630 31772 63754 31814
rect 63798 31772 63922 31814
rect 63630 31732 63632 31772
rect 63632 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63754 31772
rect 63798 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63920 31772
rect 63920 31732 63922 31772
rect 63630 31690 63754 31732
rect 63798 31690 63922 31732
rect 78750 31772 78874 31814
rect 78918 31772 79042 31814
rect 78750 31732 78752 31772
rect 78752 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78874 31772
rect 78918 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79040 31772
rect 79040 31732 79042 31772
rect 78750 31690 78874 31732
rect 78918 31690 79042 31732
rect 93870 31772 93994 31814
rect 94038 31772 94162 31814
rect 93870 31732 93872 31772
rect 93872 31732 93914 31772
rect 93914 31732 93954 31772
rect 93954 31732 93994 31772
rect 94038 31732 94078 31772
rect 94078 31732 94118 31772
rect 94118 31732 94160 31772
rect 94160 31732 94162 31772
rect 93870 31690 93994 31732
rect 94038 31690 94162 31732
rect 4390 31016 4514 31058
rect 4558 31016 4682 31058
rect 4390 30976 4392 31016
rect 4392 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4514 31016
rect 4558 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4680 31016
rect 4680 30976 4682 31016
rect 4390 30934 4514 30976
rect 4558 30934 4682 30976
rect 19510 31016 19634 31058
rect 19678 31016 19802 31058
rect 19510 30976 19512 31016
rect 19512 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19634 31016
rect 19678 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19800 31016
rect 19800 30976 19802 31016
rect 19510 30934 19634 30976
rect 19678 30934 19802 30976
rect 34630 31016 34754 31058
rect 34798 31016 34922 31058
rect 34630 30976 34632 31016
rect 34632 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34754 31016
rect 34798 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34920 31016
rect 34920 30976 34922 31016
rect 34630 30934 34754 30976
rect 34798 30934 34922 30976
rect 49750 31016 49874 31058
rect 49918 31016 50042 31058
rect 49750 30976 49752 31016
rect 49752 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49874 31016
rect 49918 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50040 31016
rect 50040 30976 50042 31016
rect 49750 30934 49874 30976
rect 49918 30934 50042 30976
rect 64870 31016 64994 31058
rect 65038 31016 65162 31058
rect 64870 30976 64872 31016
rect 64872 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64994 31016
rect 65038 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65160 31016
rect 65160 30976 65162 31016
rect 64870 30934 64994 30976
rect 65038 30934 65162 30976
rect 79990 31016 80114 31058
rect 80158 31016 80282 31058
rect 79990 30976 79992 31016
rect 79992 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80114 31016
rect 80158 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80280 31016
rect 80280 30976 80282 31016
rect 79990 30934 80114 30976
rect 80158 30934 80282 30976
rect 95110 31016 95234 31058
rect 95278 31016 95402 31058
rect 95110 30976 95112 31016
rect 95112 30976 95154 31016
rect 95154 30976 95194 31016
rect 95194 30976 95234 31016
rect 95278 30976 95318 31016
rect 95318 30976 95358 31016
rect 95358 30976 95400 31016
rect 95400 30976 95402 31016
rect 95110 30934 95234 30976
rect 95278 30934 95402 30976
rect 3150 30260 3274 30302
rect 3318 30260 3442 30302
rect 3150 30220 3152 30260
rect 3152 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3274 30260
rect 3318 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3440 30260
rect 3440 30220 3442 30260
rect 3150 30178 3274 30220
rect 3318 30178 3442 30220
rect 18270 30260 18394 30302
rect 18438 30260 18562 30302
rect 18270 30220 18272 30260
rect 18272 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18394 30260
rect 18438 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18560 30260
rect 18560 30220 18562 30260
rect 18270 30178 18394 30220
rect 18438 30178 18562 30220
rect 33390 30260 33514 30302
rect 33558 30260 33682 30302
rect 33390 30220 33392 30260
rect 33392 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33514 30260
rect 33558 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33680 30260
rect 33680 30220 33682 30260
rect 33390 30178 33514 30220
rect 33558 30178 33682 30220
rect 48510 30260 48634 30302
rect 48678 30260 48802 30302
rect 48510 30220 48512 30260
rect 48512 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48634 30260
rect 48678 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48800 30260
rect 48800 30220 48802 30260
rect 48510 30178 48634 30220
rect 48678 30178 48802 30220
rect 63630 30260 63754 30302
rect 63798 30260 63922 30302
rect 63630 30220 63632 30260
rect 63632 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63754 30260
rect 63798 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63920 30260
rect 63920 30220 63922 30260
rect 63630 30178 63754 30220
rect 63798 30178 63922 30220
rect 78750 30260 78874 30302
rect 78918 30260 79042 30302
rect 78750 30220 78752 30260
rect 78752 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78874 30260
rect 78918 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79040 30260
rect 79040 30220 79042 30260
rect 78750 30178 78874 30220
rect 78918 30178 79042 30220
rect 93870 30260 93994 30302
rect 94038 30260 94162 30302
rect 93870 30220 93872 30260
rect 93872 30220 93914 30260
rect 93914 30220 93954 30260
rect 93954 30220 93994 30260
rect 94038 30220 94078 30260
rect 94078 30220 94118 30260
rect 94118 30220 94160 30260
rect 94160 30220 94162 30260
rect 93870 30178 93994 30220
rect 94038 30178 94162 30220
rect 4390 29504 4514 29546
rect 4558 29504 4682 29546
rect 4390 29464 4392 29504
rect 4392 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4514 29504
rect 4558 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4680 29504
rect 4680 29464 4682 29504
rect 4390 29422 4514 29464
rect 4558 29422 4682 29464
rect 19510 29504 19634 29546
rect 19678 29504 19802 29546
rect 19510 29464 19512 29504
rect 19512 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19634 29504
rect 19678 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19800 29504
rect 19800 29464 19802 29504
rect 19510 29422 19634 29464
rect 19678 29422 19802 29464
rect 34630 29504 34754 29546
rect 34798 29504 34922 29546
rect 34630 29464 34632 29504
rect 34632 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34754 29504
rect 34798 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34920 29504
rect 34920 29464 34922 29504
rect 34630 29422 34754 29464
rect 34798 29422 34922 29464
rect 49750 29504 49874 29546
rect 49918 29504 50042 29546
rect 49750 29464 49752 29504
rect 49752 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49874 29504
rect 49918 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50040 29504
rect 50040 29464 50042 29504
rect 49750 29422 49874 29464
rect 49918 29422 50042 29464
rect 64870 29504 64994 29546
rect 65038 29504 65162 29546
rect 64870 29464 64872 29504
rect 64872 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64994 29504
rect 65038 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65160 29504
rect 65160 29464 65162 29504
rect 64870 29422 64994 29464
rect 65038 29422 65162 29464
rect 79990 29504 80114 29546
rect 80158 29504 80282 29546
rect 79990 29464 79992 29504
rect 79992 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80114 29504
rect 80158 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80280 29504
rect 80280 29464 80282 29504
rect 79990 29422 80114 29464
rect 80158 29422 80282 29464
rect 95110 29504 95234 29546
rect 95278 29504 95402 29546
rect 95110 29464 95112 29504
rect 95112 29464 95154 29504
rect 95154 29464 95194 29504
rect 95194 29464 95234 29504
rect 95278 29464 95318 29504
rect 95318 29464 95358 29504
rect 95358 29464 95400 29504
rect 95400 29464 95402 29504
rect 95110 29422 95234 29464
rect 95278 29422 95402 29464
rect 3150 28748 3274 28790
rect 3318 28748 3442 28790
rect 3150 28708 3152 28748
rect 3152 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3274 28748
rect 3318 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3440 28748
rect 3440 28708 3442 28748
rect 3150 28666 3274 28708
rect 3318 28666 3442 28708
rect 18270 28748 18394 28790
rect 18438 28748 18562 28790
rect 18270 28708 18272 28748
rect 18272 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18394 28748
rect 18438 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18560 28748
rect 18560 28708 18562 28748
rect 18270 28666 18394 28708
rect 18438 28666 18562 28708
rect 33390 28748 33514 28790
rect 33558 28748 33682 28790
rect 33390 28708 33392 28748
rect 33392 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33514 28748
rect 33558 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33680 28748
rect 33680 28708 33682 28748
rect 33390 28666 33514 28708
rect 33558 28666 33682 28708
rect 48510 28748 48634 28790
rect 48678 28748 48802 28790
rect 48510 28708 48512 28748
rect 48512 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48634 28748
rect 48678 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48800 28748
rect 48800 28708 48802 28748
rect 48510 28666 48634 28708
rect 48678 28666 48802 28708
rect 63630 28748 63754 28790
rect 63798 28748 63922 28790
rect 63630 28708 63632 28748
rect 63632 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63754 28748
rect 63798 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63920 28748
rect 63920 28708 63922 28748
rect 63630 28666 63754 28708
rect 63798 28666 63922 28708
rect 78750 28748 78874 28790
rect 78918 28748 79042 28790
rect 78750 28708 78752 28748
rect 78752 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78874 28748
rect 78918 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79040 28748
rect 79040 28708 79042 28748
rect 78750 28666 78874 28708
rect 78918 28666 79042 28708
rect 93870 28748 93994 28790
rect 94038 28748 94162 28790
rect 93870 28708 93872 28748
rect 93872 28708 93914 28748
rect 93914 28708 93954 28748
rect 93954 28708 93994 28748
rect 94038 28708 94078 28748
rect 94078 28708 94118 28748
rect 94118 28708 94160 28748
rect 94160 28708 94162 28748
rect 93870 28666 93994 28708
rect 94038 28666 94162 28708
rect 4390 27992 4514 28034
rect 4558 27992 4682 28034
rect 4390 27952 4392 27992
rect 4392 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4514 27992
rect 4558 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4680 27992
rect 4680 27952 4682 27992
rect 4390 27910 4514 27952
rect 4558 27910 4682 27952
rect 19510 27992 19634 28034
rect 19678 27992 19802 28034
rect 19510 27952 19512 27992
rect 19512 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19634 27992
rect 19678 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19800 27992
rect 19800 27952 19802 27992
rect 19510 27910 19634 27952
rect 19678 27910 19802 27952
rect 34630 27992 34754 28034
rect 34798 27992 34922 28034
rect 34630 27952 34632 27992
rect 34632 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34754 27992
rect 34798 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34920 27992
rect 34920 27952 34922 27992
rect 34630 27910 34754 27952
rect 34798 27910 34922 27952
rect 49750 27992 49874 28034
rect 49918 27992 50042 28034
rect 49750 27952 49752 27992
rect 49752 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49874 27992
rect 49918 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50040 27992
rect 50040 27952 50042 27992
rect 49750 27910 49874 27952
rect 49918 27910 50042 27952
rect 64870 27992 64994 28034
rect 65038 27992 65162 28034
rect 64870 27952 64872 27992
rect 64872 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64994 27992
rect 65038 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65160 27992
rect 65160 27952 65162 27992
rect 64870 27910 64994 27952
rect 65038 27910 65162 27952
rect 79990 27992 80114 28034
rect 80158 27992 80282 28034
rect 79990 27952 79992 27992
rect 79992 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80114 27992
rect 80158 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80280 27992
rect 80280 27952 80282 27992
rect 79990 27910 80114 27952
rect 80158 27910 80282 27952
rect 95110 27992 95234 28034
rect 95278 27992 95402 28034
rect 95110 27952 95112 27992
rect 95112 27952 95154 27992
rect 95154 27952 95194 27992
rect 95194 27952 95234 27992
rect 95278 27952 95318 27992
rect 95318 27952 95358 27992
rect 95358 27952 95400 27992
rect 95400 27952 95402 27992
rect 95110 27910 95234 27952
rect 95278 27910 95402 27952
rect 3150 27236 3274 27278
rect 3318 27236 3442 27278
rect 3150 27196 3152 27236
rect 3152 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3274 27236
rect 3318 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3440 27236
rect 3440 27196 3442 27236
rect 3150 27154 3274 27196
rect 3318 27154 3442 27196
rect 18270 27236 18394 27278
rect 18438 27236 18562 27278
rect 18270 27196 18272 27236
rect 18272 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18394 27236
rect 18438 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18560 27236
rect 18560 27196 18562 27236
rect 18270 27154 18394 27196
rect 18438 27154 18562 27196
rect 33390 27236 33514 27278
rect 33558 27236 33682 27278
rect 33390 27196 33392 27236
rect 33392 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33514 27236
rect 33558 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33680 27236
rect 33680 27196 33682 27236
rect 33390 27154 33514 27196
rect 33558 27154 33682 27196
rect 48510 27236 48634 27278
rect 48678 27236 48802 27278
rect 48510 27196 48512 27236
rect 48512 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48634 27236
rect 48678 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48800 27236
rect 48800 27196 48802 27236
rect 48510 27154 48634 27196
rect 48678 27154 48802 27196
rect 63630 27236 63754 27278
rect 63798 27236 63922 27278
rect 63630 27196 63632 27236
rect 63632 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63754 27236
rect 63798 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63920 27236
rect 63920 27196 63922 27236
rect 63630 27154 63754 27196
rect 63798 27154 63922 27196
rect 78750 27236 78874 27278
rect 78918 27236 79042 27278
rect 78750 27196 78752 27236
rect 78752 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78874 27236
rect 78918 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79040 27236
rect 79040 27196 79042 27236
rect 78750 27154 78874 27196
rect 78918 27154 79042 27196
rect 93870 27236 93994 27278
rect 94038 27236 94162 27278
rect 93870 27196 93872 27236
rect 93872 27196 93914 27236
rect 93914 27196 93954 27236
rect 93954 27196 93994 27236
rect 94038 27196 94078 27236
rect 94078 27196 94118 27236
rect 94118 27196 94160 27236
rect 94160 27196 94162 27236
rect 93870 27154 93994 27196
rect 94038 27154 94162 27196
rect 4390 26480 4514 26522
rect 4558 26480 4682 26522
rect 4390 26440 4392 26480
rect 4392 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4514 26480
rect 4558 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4680 26480
rect 4680 26440 4682 26480
rect 4390 26398 4514 26440
rect 4558 26398 4682 26440
rect 19510 26480 19634 26522
rect 19678 26480 19802 26522
rect 19510 26440 19512 26480
rect 19512 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19634 26480
rect 19678 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19800 26480
rect 19800 26440 19802 26480
rect 19510 26398 19634 26440
rect 19678 26398 19802 26440
rect 34630 26480 34754 26522
rect 34798 26480 34922 26522
rect 34630 26440 34632 26480
rect 34632 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34754 26480
rect 34798 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34920 26480
rect 34920 26440 34922 26480
rect 34630 26398 34754 26440
rect 34798 26398 34922 26440
rect 49750 26480 49874 26522
rect 49918 26480 50042 26522
rect 49750 26440 49752 26480
rect 49752 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49874 26480
rect 49918 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50040 26480
rect 50040 26440 50042 26480
rect 49750 26398 49874 26440
rect 49918 26398 50042 26440
rect 64870 26480 64994 26522
rect 65038 26480 65162 26522
rect 64870 26440 64872 26480
rect 64872 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64994 26480
rect 65038 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65160 26480
rect 65160 26440 65162 26480
rect 64870 26398 64994 26440
rect 65038 26398 65162 26440
rect 79990 26480 80114 26522
rect 80158 26480 80282 26522
rect 79990 26440 79992 26480
rect 79992 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80114 26480
rect 80158 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80280 26480
rect 80280 26440 80282 26480
rect 79990 26398 80114 26440
rect 80158 26398 80282 26440
rect 95110 26480 95234 26522
rect 95278 26480 95402 26522
rect 95110 26440 95112 26480
rect 95112 26440 95154 26480
rect 95154 26440 95194 26480
rect 95194 26440 95234 26480
rect 95278 26440 95318 26480
rect 95318 26440 95358 26480
rect 95358 26440 95400 26480
rect 95400 26440 95402 26480
rect 95110 26398 95234 26440
rect 95278 26398 95402 26440
rect 3150 25724 3274 25766
rect 3318 25724 3442 25766
rect 3150 25684 3152 25724
rect 3152 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3274 25724
rect 3318 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3440 25724
rect 3440 25684 3442 25724
rect 3150 25642 3274 25684
rect 3318 25642 3442 25684
rect 18270 25724 18394 25766
rect 18438 25724 18562 25766
rect 18270 25684 18272 25724
rect 18272 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18394 25724
rect 18438 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18560 25724
rect 18560 25684 18562 25724
rect 18270 25642 18394 25684
rect 18438 25642 18562 25684
rect 33390 25724 33514 25766
rect 33558 25724 33682 25766
rect 33390 25684 33392 25724
rect 33392 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33514 25724
rect 33558 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33680 25724
rect 33680 25684 33682 25724
rect 33390 25642 33514 25684
rect 33558 25642 33682 25684
rect 48510 25724 48634 25766
rect 48678 25724 48802 25766
rect 48510 25684 48512 25724
rect 48512 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48634 25724
rect 48678 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48800 25724
rect 48800 25684 48802 25724
rect 48510 25642 48634 25684
rect 48678 25642 48802 25684
rect 63630 25724 63754 25766
rect 63798 25724 63922 25766
rect 63630 25684 63632 25724
rect 63632 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63754 25724
rect 63798 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63920 25724
rect 63920 25684 63922 25724
rect 63630 25642 63754 25684
rect 63798 25642 63922 25684
rect 78750 25724 78874 25766
rect 78918 25724 79042 25766
rect 78750 25684 78752 25724
rect 78752 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78874 25724
rect 78918 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79040 25724
rect 79040 25684 79042 25724
rect 78750 25642 78874 25684
rect 78918 25642 79042 25684
rect 93870 25724 93994 25766
rect 94038 25724 94162 25766
rect 93870 25684 93872 25724
rect 93872 25684 93914 25724
rect 93914 25684 93954 25724
rect 93954 25684 93994 25724
rect 94038 25684 94078 25724
rect 94078 25684 94118 25724
rect 94118 25684 94160 25724
rect 94160 25684 94162 25724
rect 93870 25642 93994 25684
rect 94038 25642 94162 25684
rect 4390 24968 4514 25010
rect 4558 24968 4682 25010
rect 4390 24928 4392 24968
rect 4392 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4514 24968
rect 4558 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4680 24968
rect 4680 24928 4682 24968
rect 4390 24886 4514 24928
rect 4558 24886 4682 24928
rect 19510 24968 19634 25010
rect 19678 24968 19802 25010
rect 19510 24928 19512 24968
rect 19512 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19634 24968
rect 19678 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19800 24968
rect 19800 24928 19802 24968
rect 19510 24886 19634 24928
rect 19678 24886 19802 24928
rect 34630 24968 34754 25010
rect 34798 24968 34922 25010
rect 34630 24928 34632 24968
rect 34632 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34754 24968
rect 34798 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34920 24968
rect 34920 24928 34922 24968
rect 34630 24886 34754 24928
rect 34798 24886 34922 24928
rect 49750 24968 49874 25010
rect 49918 24968 50042 25010
rect 49750 24928 49752 24968
rect 49752 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49874 24968
rect 49918 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50040 24968
rect 50040 24928 50042 24968
rect 49750 24886 49874 24928
rect 49918 24886 50042 24928
rect 64870 24968 64994 25010
rect 65038 24968 65162 25010
rect 64870 24928 64872 24968
rect 64872 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64994 24968
rect 65038 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65160 24968
rect 65160 24928 65162 24968
rect 64870 24886 64994 24928
rect 65038 24886 65162 24928
rect 79990 24968 80114 25010
rect 80158 24968 80282 25010
rect 79990 24928 79992 24968
rect 79992 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80114 24968
rect 80158 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80280 24968
rect 80280 24928 80282 24968
rect 79990 24886 80114 24928
rect 80158 24886 80282 24928
rect 95110 24968 95234 25010
rect 95278 24968 95402 25010
rect 95110 24928 95112 24968
rect 95112 24928 95154 24968
rect 95154 24928 95194 24968
rect 95194 24928 95234 24968
rect 95278 24928 95318 24968
rect 95318 24928 95358 24968
rect 95358 24928 95400 24968
rect 95400 24928 95402 24968
rect 95110 24886 95234 24928
rect 95278 24886 95402 24928
rect 3150 24212 3274 24254
rect 3318 24212 3442 24254
rect 3150 24172 3152 24212
rect 3152 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3274 24212
rect 3318 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3440 24212
rect 3440 24172 3442 24212
rect 3150 24130 3274 24172
rect 3318 24130 3442 24172
rect 18270 24212 18394 24254
rect 18438 24212 18562 24254
rect 18270 24172 18272 24212
rect 18272 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18394 24212
rect 18438 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18560 24212
rect 18560 24172 18562 24212
rect 18270 24130 18394 24172
rect 18438 24130 18562 24172
rect 33390 24212 33514 24254
rect 33558 24212 33682 24254
rect 33390 24172 33392 24212
rect 33392 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33514 24212
rect 33558 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33680 24212
rect 33680 24172 33682 24212
rect 33390 24130 33514 24172
rect 33558 24130 33682 24172
rect 48510 24212 48634 24254
rect 48678 24212 48802 24254
rect 48510 24172 48512 24212
rect 48512 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48634 24212
rect 48678 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48800 24212
rect 48800 24172 48802 24212
rect 48510 24130 48634 24172
rect 48678 24130 48802 24172
rect 63630 24212 63754 24254
rect 63798 24212 63922 24254
rect 63630 24172 63632 24212
rect 63632 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63754 24212
rect 63798 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63920 24212
rect 63920 24172 63922 24212
rect 63630 24130 63754 24172
rect 63798 24130 63922 24172
rect 78750 24212 78874 24254
rect 78918 24212 79042 24254
rect 78750 24172 78752 24212
rect 78752 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78874 24212
rect 78918 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79040 24212
rect 79040 24172 79042 24212
rect 78750 24130 78874 24172
rect 78918 24130 79042 24172
rect 93870 24212 93994 24254
rect 94038 24212 94162 24254
rect 93870 24172 93872 24212
rect 93872 24172 93914 24212
rect 93914 24172 93954 24212
rect 93954 24172 93994 24212
rect 94038 24172 94078 24212
rect 94078 24172 94118 24212
rect 94118 24172 94160 24212
rect 94160 24172 94162 24212
rect 93870 24130 93994 24172
rect 94038 24130 94162 24172
rect 4390 23456 4514 23498
rect 4558 23456 4682 23498
rect 4390 23416 4392 23456
rect 4392 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4514 23456
rect 4558 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4680 23456
rect 4680 23416 4682 23456
rect 4390 23374 4514 23416
rect 4558 23374 4682 23416
rect 19510 23456 19634 23498
rect 19678 23456 19802 23498
rect 19510 23416 19512 23456
rect 19512 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19634 23456
rect 19678 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19800 23456
rect 19800 23416 19802 23456
rect 19510 23374 19634 23416
rect 19678 23374 19802 23416
rect 34630 23456 34754 23498
rect 34798 23456 34922 23498
rect 34630 23416 34632 23456
rect 34632 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34754 23456
rect 34798 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34920 23456
rect 34920 23416 34922 23456
rect 34630 23374 34754 23416
rect 34798 23374 34922 23416
rect 49750 23456 49874 23498
rect 49918 23456 50042 23498
rect 49750 23416 49752 23456
rect 49752 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49874 23456
rect 49918 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50040 23456
rect 50040 23416 50042 23456
rect 49750 23374 49874 23416
rect 49918 23374 50042 23416
rect 64870 23456 64994 23498
rect 65038 23456 65162 23498
rect 64870 23416 64872 23456
rect 64872 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64994 23456
rect 65038 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65160 23456
rect 65160 23416 65162 23456
rect 64870 23374 64994 23416
rect 65038 23374 65162 23416
rect 79990 23456 80114 23498
rect 80158 23456 80282 23498
rect 79990 23416 79992 23456
rect 79992 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80114 23456
rect 80158 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80280 23456
rect 80280 23416 80282 23456
rect 79990 23374 80114 23416
rect 80158 23374 80282 23416
rect 95110 23456 95234 23498
rect 95278 23456 95402 23498
rect 95110 23416 95112 23456
rect 95112 23416 95154 23456
rect 95154 23416 95194 23456
rect 95194 23416 95234 23456
rect 95278 23416 95318 23456
rect 95318 23416 95358 23456
rect 95358 23416 95400 23456
rect 95400 23416 95402 23456
rect 95110 23374 95234 23416
rect 95278 23374 95402 23416
rect 3150 22700 3274 22742
rect 3318 22700 3442 22742
rect 3150 22660 3152 22700
rect 3152 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3274 22700
rect 3318 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3440 22700
rect 3440 22660 3442 22700
rect 3150 22618 3274 22660
rect 3318 22618 3442 22660
rect 18270 22700 18394 22742
rect 18438 22700 18562 22742
rect 18270 22660 18272 22700
rect 18272 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18394 22700
rect 18438 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18560 22700
rect 18560 22660 18562 22700
rect 18270 22618 18394 22660
rect 18438 22618 18562 22660
rect 33390 22700 33514 22742
rect 33558 22700 33682 22742
rect 33390 22660 33392 22700
rect 33392 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33514 22700
rect 33558 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33680 22700
rect 33680 22660 33682 22700
rect 33390 22618 33514 22660
rect 33558 22618 33682 22660
rect 48510 22700 48634 22742
rect 48678 22700 48802 22742
rect 48510 22660 48512 22700
rect 48512 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48634 22700
rect 48678 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48800 22700
rect 48800 22660 48802 22700
rect 48510 22618 48634 22660
rect 48678 22618 48802 22660
rect 63630 22700 63754 22742
rect 63798 22700 63922 22742
rect 63630 22660 63632 22700
rect 63632 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63754 22700
rect 63798 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63920 22700
rect 63920 22660 63922 22700
rect 63630 22618 63754 22660
rect 63798 22618 63922 22660
rect 78750 22700 78874 22742
rect 78918 22700 79042 22742
rect 78750 22660 78752 22700
rect 78752 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78874 22700
rect 78918 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79040 22700
rect 79040 22660 79042 22700
rect 78750 22618 78874 22660
rect 78918 22618 79042 22660
rect 93870 22700 93994 22742
rect 94038 22700 94162 22742
rect 93870 22660 93872 22700
rect 93872 22660 93914 22700
rect 93914 22660 93954 22700
rect 93954 22660 93994 22700
rect 94038 22660 94078 22700
rect 94078 22660 94118 22700
rect 94118 22660 94160 22700
rect 94160 22660 94162 22700
rect 93870 22618 93994 22660
rect 94038 22618 94162 22660
rect 4390 21944 4514 21986
rect 4558 21944 4682 21986
rect 4390 21904 4392 21944
rect 4392 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4514 21944
rect 4558 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4680 21944
rect 4680 21904 4682 21944
rect 4390 21862 4514 21904
rect 4558 21862 4682 21904
rect 19510 21944 19634 21986
rect 19678 21944 19802 21986
rect 19510 21904 19512 21944
rect 19512 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19634 21944
rect 19678 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19800 21944
rect 19800 21904 19802 21944
rect 19510 21862 19634 21904
rect 19678 21862 19802 21904
rect 34630 21944 34754 21986
rect 34798 21944 34922 21986
rect 34630 21904 34632 21944
rect 34632 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34754 21944
rect 34798 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34920 21944
rect 34920 21904 34922 21944
rect 34630 21862 34754 21904
rect 34798 21862 34922 21904
rect 49750 21944 49874 21986
rect 49918 21944 50042 21986
rect 49750 21904 49752 21944
rect 49752 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49874 21944
rect 49918 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50040 21944
rect 50040 21904 50042 21944
rect 49750 21862 49874 21904
rect 49918 21862 50042 21904
rect 64870 21944 64994 21986
rect 65038 21944 65162 21986
rect 64870 21904 64872 21944
rect 64872 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64994 21944
rect 65038 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65160 21944
rect 65160 21904 65162 21944
rect 64870 21862 64994 21904
rect 65038 21862 65162 21904
rect 79990 21944 80114 21986
rect 80158 21944 80282 21986
rect 79990 21904 79992 21944
rect 79992 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80114 21944
rect 80158 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80280 21944
rect 80280 21904 80282 21944
rect 79990 21862 80114 21904
rect 80158 21862 80282 21904
rect 95110 21944 95234 21986
rect 95278 21944 95402 21986
rect 95110 21904 95112 21944
rect 95112 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95234 21944
rect 95278 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95400 21944
rect 95400 21904 95402 21944
rect 95110 21862 95234 21904
rect 95278 21862 95402 21904
rect 3150 21188 3274 21230
rect 3318 21188 3442 21230
rect 3150 21148 3152 21188
rect 3152 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3274 21188
rect 3318 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3440 21188
rect 3440 21148 3442 21188
rect 3150 21106 3274 21148
rect 3318 21106 3442 21148
rect 18270 21188 18394 21230
rect 18438 21188 18562 21230
rect 18270 21148 18272 21188
rect 18272 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18394 21188
rect 18438 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18560 21188
rect 18560 21148 18562 21188
rect 18270 21106 18394 21148
rect 18438 21106 18562 21148
rect 33390 21188 33514 21230
rect 33558 21188 33682 21230
rect 33390 21148 33392 21188
rect 33392 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33514 21188
rect 33558 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33680 21188
rect 33680 21148 33682 21188
rect 33390 21106 33514 21148
rect 33558 21106 33682 21148
rect 48510 21188 48634 21230
rect 48678 21188 48802 21230
rect 48510 21148 48512 21188
rect 48512 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48634 21188
rect 48678 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48800 21188
rect 48800 21148 48802 21188
rect 48510 21106 48634 21148
rect 48678 21106 48802 21148
rect 63630 21188 63754 21230
rect 63798 21188 63922 21230
rect 63630 21148 63632 21188
rect 63632 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63754 21188
rect 63798 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63920 21188
rect 63920 21148 63922 21188
rect 63630 21106 63754 21148
rect 63798 21106 63922 21148
rect 78750 21188 78874 21230
rect 78918 21188 79042 21230
rect 78750 21148 78752 21188
rect 78752 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78874 21188
rect 78918 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79040 21188
rect 79040 21148 79042 21188
rect 78750 21106 78874 21148
rect 78918 21106 79042 21148
rect 93870 21188 93994 21230
rect 94038 21188 94162 21230
rect 93870 21148 93872 21188
rect 93872 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93994 21188
rect 94038 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94160 21188
rect 94160 21148 94162 21188
rect 93870 21106 93994 21148
rect 94038 21106 94162 21148
rect 4390 20432 4514 20474
rect 4558 20432 4682 20474
rect 4390 20392 4392 20432
rect 4392 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4514 20432
rect 4558 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4680 20432
rect 4680 20392 4682 20432
rect 4390 20350 4514 20392
rect 4558 20350 4682 20392
rect 19510 20432 19634 20474
rect 19678 20432 19802 20474
rect 19510 20392 19512 20432
rect 19512 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19634 20432
rect 19678 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19800 20432
rect 19800 20392 19802 20432
rect 19510 20350 19634 20392
rect 19678 20350 19802 20392
rect 34630 20432 34754 20474
rect 34798 20432 34922 20474
rect 34630 20392 34632 20432
rect 34632 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34754 20432
rect 34798 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34920 20432
rect 34920 20392 34922 20432
rect 34630 20350 34754 20392
rect 34798 20350 34922 20392
rect 49750 20432 49874 20474
rect 49918 20432 50042 20474
rect 49750 20392 49752 20432
rect 49752 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49874 20432
rect 49918 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50040 20432
rect 50040 20392 50042 20432
rect 49750 20350 49874 20392
rect 49918 20350 50042 20392
rect 64870 20432 64994 20474
rect 65038 20432 65162 20474
rect 64870 20392 64872 20432
rect 64872 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64994 20432
rect 65038 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65160 20432
rect 65160 20392 65162 20432
rect 64870 20350 64994 20392
rect 65038 20350 65162 20392
rect 79990 20432 80114 20474
rect 80158 20432 80282 20474
rect 79990 20392 79992 20432
rect 79992 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80114 20432
rect 80158 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80280 20432
rect 80280 20392 80282 20432
rect 79990 20350 80114 20392
rect 80158 20350 80282 20392
rect 95110 20432 95234 20474
rect 95278 20432 95402 20474
rect 95110 20392 95112 20432
rect 95112 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95234 20432
rect 95278 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95400 20432
rect 95400 20392 95402 20432
rect 95110 20350 95234 20392
rect 95278 20350 95402 20392
rect 3150 19676 3274 19718
rect 3318 19676 3442 19718
rect 3150 19636 3152 19676
rect 3152 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3274 19676
rect 3318 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3440 19676
rect 3440 19636 3442 19676
rect 3150 19594 3274 19636
rect 3318 19594 3442 19636
rect 18270 19676 18394 19718
rect 18438 19676 18562 19718
rect 18270 19636 18272 19676
rect 18272 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18394 19676
rect 18438 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18560 19676
rect 18560 19636 18562 19676
rect 18270 19594 18394 19636
rect 18438 19594 18562 19636
rect 33390 19676 33514 19718
rect 33558 19676 33682 19718
rect 33390 19636 33392 19676
rect 33392 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33514 19676
rect 33558 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33680 19676
rect 33680 19636 33682 19676
rect 33390 19594 33514 19636
rect 33558 19594 33682 19636
rect 48510 19676 48634 19718
rect 48678 19676 48802 19718
rect 48510 19636 48512 19676
rect 48512 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48634 19676
rect 48678 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48800 19676
rect 48800 19636 48802 19676
rect 48510 19594 48634 19636
rect 48678 19594 48802 19636
rect 63630 19676 63754 19718
rect 63798 19676 63922 19718
rect 63630 19636 63632 19676
rect 63632 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63754 19676
rect 63798 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63920 19676
rect 63920 19636 63922 19676
rect 63630 19594 63754 19636
rect 63798 19594 63922 19636
rect 78750 19676 78874 19718
rect 78918 19676 79042 19718
rect 78750 19636 78752 19676
rect 78752 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78874 19676
rect 78918 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79040 19676
rect 79040 19636 79042 19676
rect 78750 19594 78874 19636
rect 78918 19594 79042 19636
rect 93870 19676 93994 19718
rect 94038 19676 94162 19718
rect 93870 19636 93872 19676
rect 93872 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93994 19676
rect 94038 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94160 19676
rect 94160 19636 94162 19676
rect 93870 19594 93994 19636
rect 94038 19594 94162 19636
rect 4390 18920 4514 18962
rect 4558 18920 4682 18962
rect 4390 18880 4392 18920
rect 4392 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4514 18920
rect 4558 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4680 18920
rect 4680 18880 4682 18920
rect 4390 18838 4514 18880
rect 4558 18838 4682 18880
rect 19510 18920 19634 18962
rect 19678 18920 19802 18962
rect 19510 18880 19512 18920
rect 19512 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19634 18920
rect 19678 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19800 18920
rect 19800 18880 19802 18920
rect 19510 18838 19634 18880
rect 19678 18838 19802 18880
rect 34630 18920 34754 18962
rect 34798 18920 34922 18962
rect 34630 18880 34632 18920
rect 34632 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34754 18920
rect 34798 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34920 18920
rect 34920 18880 34922 18920
rect 34630 18838 34754 18880
rect 34798 18838 34922 18880
rect 49750 18920 49874 18962
rect 49918 18920 50042 18962
rect 49750 18880 49752 18920
rect 49752 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49874 18920
rect 49918 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50040 18920
rect 50040 18880 50042 18920
rect 49750 18838 49874 18880
rect 49918 18838 50042 18880
rect 64870 18920 64994 18962
rect 65038 18920 65162 18962
rect 64870 18880 64872 18920
rect 64872 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64994 18920
rect 65038 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65160 18920
rect 65160 18880 65162 18920
rect 64870 18838 64994 18880
rect 65038 18838 65162 18880
rect 79990 18920 80114 18962
rect 80158 18920 80282 18962
rect 79990 18880 79992 18920
rect 79992 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80114 18920
rect 80158 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80280 18920
rect 80280 18880 80282 18920
rect 79990 18838 80114 18880
rect 80158 18838 80282 18880
rect 95110 18920 95234 18962
rect 95278 18920 95402 18962
rect 95110 18880 95112 18920
rect 95112 18880 95154 18920
rect 95154 18880 95194 18920
rect 95194 18880 95234 18920
rect 95278 18880 95318 18920
rect 95318 18880 95358 18920
rect 95358 18880 95400 18920
rect 95400 18880 95402 18920
rect 95110 18838 95234 18880
rect 95278 18838 95402 18880
rect 3150 18164 3274 18206
rect 3318 18164 3442 18206
rect 3150 18124 3152 18164
rect 3152 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3274 18164
rect 3318 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3440 18164
rect 3440 18124 3442 18164
rect 3150 18082 3274 18124
rect 3318 18082 3442 18124
rect 18270 18164 18394 18206
rect 18438 18164 18562 18206
rect 18270 18124 18272 18164
rect 18272 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18394 18164
rect 18438 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18560 18164
rect 18560 18124 18562 18164
rect 18270 18082 18394 18124
rect 18438 18082 18562 18124
rect 33390 18164 33514 18206
rect 33558 18164 33682 18206
rect 33390 18124 33392 18164
rect 33392 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33514 18164
rect 33558 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33680 18164
rect 33680 18124 33682 18164
rect 33390 18082 33514 18124
rect 33558 18082 33682 18124
rect 48510 18164 48634 18206
rect 48678 18164 48802 18206
rect 48510 18124 48512 18164
rect 48512 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48634 18164
rect 48678 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48800 18164
rect 48800 18124 48802 18164
rect 48510 18082 48634 18124
rect 48678 18082 48802 18124
rect 63630 18164 63754 18206
rect 63798 18164 63922 18206
rect 63630 18124 63632 18164
rect 63632 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63754 18164
rect 63798 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63920 18164
rect 63920 18124 63922 18164
rect 63630 18082 63754 18124
rect 63798 18082 63922 18124
rect 78750 18164 78874 18206
rect 78918 18164 79042 18206
rect 78750 18124 78752 18164
rect 78752 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78874 18164
rect 78918 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79040 18164
rect 79040 18124 79042 18164
rect 78750 18082 78874 18124
rect 78918 18082 79042 18124
rect 93870 18164 93994 18206
rect 94038 18164 94162 18206
rect 93870 18124 93872 18164
rect 93872 18124 93914 18164
rect 93914 18124 93954 18164
rect 93954 18124 93994 18164
rect 94038 18124 94078 18164
rect 94078 18124 94118 18164
rect 94118 18124 94160 18164
rect 94160 18124 94162 18164
rect 93870 18082 93994 18124
rect 94038 18082 94162 18124
rect 4390 17408 4514 17450
rect 4558 17408 4682 17450
rect 4390 17368 4392 17408
rect 4392 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4514 17408
rect 4558 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4680 17408
rect 4680 17368 4682 17408
rect 4390 17326 4514 17368
rect 4558 17326 4682 17368
rect 19510 17408 19634 17450
rect 19678 17408 19802 17450
rect 19510 17368 19512 17408
rect 19512 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19634 17408
rect 19678 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19800 17408
rect 19800 17368 19802 17408
rect 19510 17326 19634 17368
rect 19678 17326 19802 17368
rect 34630 17408 34754 17450
rect 34798 17408 34922 17450
rect 34630 17368 34632 17408
rect 34632 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34754 17408
rect 34798 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34920 17408
rect 34920 17368 34922 17408
rect 34630 17326 34754 17368
rect 34798 17326 34922 17368
rect 49750 17408 49874 17450
rect 49918 17408 50042 17450
rect 49750 17368 49752 17408
rect 49752 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49874 17408
rect 49918 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50040 17408
rect 50040 17368 50042 17408
rect 49750 17326 49874 17368
rect 49918 17326 50042 17368
rect 64870 17408 64994 17450
rect 65038 17408 65162 17450
rect 64870 17368 64872 17408
rect 64872 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64994 17408
rect 65038 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65160 17408
rect 65160 17368 65162 17408
rect 64870 17326 64994 17368
rect 65038 17326 65162 17368
rect 79990 17408 80114 17450
rect 80158 17408 80282 17450
rect 79990 17368 79992 17408
rect 79992 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80114 17408
rect 80158 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80280 17408
rect 80280 17368 80282 17408
rect 79990 17326 80114 17368
rect 80158 17326 80282 17368
rect 95110 17408 95234 17450
rect 95278 17408 95402 17450
rect 95110 17368 95112 17408
rect 95112 17368 95154 17408
rect 95154 17368 95194 17408
rect 95194 17368 95234 17408
rect 95278 17368 95318 17408
rect 95318 17368 95358 17408
rect 95358 17368 95400 17408
rect 95400 17368 95402 17408
rect 95110 17326 95234 17368
rect 95278 17326 95402 17368
rect 3150 16652 3274 16694
rect 3318 16652 3442 16694
rect 3150 16612 3152 16652
rect 3152 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3274 16652
rect 3318 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3440 16652
rect 3440 16612 3442 16652
rect 3150 16570 3274 16612
rect 3318 16570 3442 16612
rect 18270 16652 18394 16694
rect 18438 16652 18562 16694
rect 18270 16612 18272 16652
rect 18272 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18394 16652
rect 18438 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18560 16652
rect 18560 16612 18562 16652
rect 18270 16570 18394 16612
rect 18438 16570 18562 16612
rect 33390 16652 33514 16694
rect 33558 16652 33682 16694
rect 33390 16612 33392 16652
rect 33392 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33514 16652
rect 33558 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33680 16652
rect 33680 16612 33682 16652
rect 33390 16570 33514 16612
rect 33558 16570 33682 16612
rect 48510 16652 48634 16694
rect 48678 16652 48802 16694
rect 48510 16612 48512 16652
rect 48512 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48634 16652
rect 48678 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48800 16652
rect 48800 16612 48802 16652
rect 48510 16570 48634 16612
rect 48678 16570 48802 16612
rect 63630 16652 63754 16694
rect 63798 16652 63922 16694
rect 63630 16612 63632 16652
rect 63632 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63754 16652
rect 63798 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63920 16652
rect 63920 16612 63922 16652
rect 63630 16570 63754 16612
rect 63798 16570 63922 16612
rect 78750 16652 78874 16694
rect 78918 16652 79042 16694
rect 78750 16612 78752 16652
rect 78752 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78874 16652
rect 78918 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79040 16652
rect 79040 16612 79042 16652
rect 78750 16570 78874 16612
rect 78918 16570 79042 16612
rect 93870 16652 93994 16694
rect 94038 16652 94162 16694
rect 93870 16612 93872 16652
rect 93872 16612 93914 16652
rect 93914 16612 93954 16652
rect 93954 16612 93994 16652
rect 94038 16612 94078 16652
rect 94078 16612 94118 16652
rect 94118 16612 94160 16652
rect 94160 16612 94162 16652
rect 93870 16570 93994 16612
rect 94038 16570 94162 16612
rect 4390 15896 4514 15938
rect 4558 15896 4682 15938
rect 4390 15856 4392 15896
rect 4392 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4514 15896
rect 4558 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4680 15896
rect 4680 15856 4682 15896
rect 4390 15814 4514 15856
rect 4558 15814 4682 15856
rect 19510 15896 19634 15938
rect 19678 15896 19802 15938
rect 19510 15856 19512 15896
rect 19512 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19634 15896
rect 19678 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19800 15896
rect 19800 15856 19802 15896
rect 19510 15814 19634 15856
rect 19678 15814 19802 15856
rect 34630 15896 34754 15938
rect 34798 15896 34922 15938
rect 34630 15856 34632 15896
rect 34632 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34754 15896
rect 34798 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34920 15896
rect 34920 15856 34922 15896
rect 34630 15814 34754 15856
rect 34798 15814 34922 15856
rect 49750 15896 49874 15938
rect 49918 15896 50042 15938
rect 49750 15856 49752 15896
rect 49752 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49874 15896
rect 49918 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50040 15896
rect 50040 15856 50042 15896
rect 49750 15814 49874 15856
rect 49918 15814 50042 15856
rect 64870 15896 64994 15938
rect 65038 15896 65162 15938
rect 64870 15856 64872 15896
rect 64872 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64994 15896
rect 65038 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65160 15896
rect 65160 15856 65162 15896
rect 64870 15814 64994 15856
rect 65038 15814 65162 15856
rect 79990 15896 80114 15938
rect 80158 15896 80282 15938
rect 79990 15856 79992 15896
rect 79992 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80114 15896
rect 80158 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80280 15896
rect 80280 15856 80282 15896
rect 79990 15814 80114 15856
rect 80158 15814 80282 15856
rect 95110 15896 95234 15938
rect 95278 15896 95402 15938
rect 95110 15856 95112 15896
rect 95112 15856 95154 15896
rect 95154 15856 95194 15896
rect 95194 15856 95234 15896
rect 95278 15856 95318 15896
rect 95318 15856 95358 15896
rect 95358 15856 95400 15896
rect 95400 15856 95402 15896
rect 95110 15814 95234 15856
rect 95278 15814 95402 15856
rect 3150 15140 3274 15182
rect 3318 15140 3442 15182
rect 3150 15100 3152 15140
rect 3152 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3274 15140
rect 3318 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3440 15140
rect 3440 15100 3442 15140
rect 3150 15058 3274 15100
rect 3318 15058 3442 15100
rect 18270 15140 18394 15182
rect 18438 15140 18562 15182
rect 18270 15100 18272 15140
rect 18272 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18394 15140
rect 18438 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18560 15140
rect 18560 15100 18562 15140
rect 18270 15058 18394 15100
rect 18438 15058 18562 15100
rect 33390 15140 33514 15182
rect 33558 15140 33682 15182
rect 33390 15100 33392 15140
rect 33392 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33514 15140
rect 33558 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33680 15140
rect 33680 15100 33682 15140
rect 33390 15058 33514 15100
rect 33558 15058 33682 15100
rect 48510 15140 48634 15182
rect 48678 15140 48802 15182
rect 48510 15100 48512 15140
rect 48512 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48634 15140
rect 48678 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48800 15140
rect 48800 15100 48802 15140
rect 48510 15058 48634 15100
rect 48678 15058 48802 15100
rect 63630 15140 63754 15182
rect 63798 15140 63922 15182
rect 63630 15100 63632 15140
rect 63632 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63754 15140
rect 63798 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63920 15140
rect 63920 15100 63922 15140
rect 63630 15058 63754 15100
rect 63798 15058 63922 15100
rect 78750 15140 78874 15182
rect 78918 15140 79042 15182
rect 78750 15100 78752 15140
rect 78752 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78874 15140
rect 78918 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79040 15140
rect 79040 15100 79042 15140
rect 78750 15058 78874 15100
rect 78918 15058 79042 15100
rect 93870 15140 93994 15182
rect 94038 15140 94162 15182
rect 93870 15100 93872 15140
rect 93872 15100 93914 15140
rect 93914 15100 93954 15140
rect 93954 15100 93994 15140
rect 94038 15100 94078 15140
rect 94078 15100 94118 15140
rect 94118 15100 94160 15140
rect 94160 15100 94162 15140
rect 93870 15058 93994 15100
rect 94038 15058 94162 15100
rect 4390 14384 4514 14426
rect 4558 14384 4682 14426
rect 4390 14344 4392 14384
rect 4392 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4514 14384
rect 4558 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4680 14384
rect 4680 14344 4682 14384
rect 4390 14302 4514 14344
rect 4558 14302 4682 14344
rect 19510 14384 19634 14426
rect 19678 14384 19802 14426
rect 19510 14344 19512 14384
rect 19512 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19634 14384
rect 19678 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19800 14384
rect 19800 14344 19802 14384
rect 19510 14302 19634 14344
rect 19678 14302 19802 14344
rect 34630 14384 34754 14426
rect 34798 14384 34922 14426
rect 34630 14344 34632 14384
rect 34632 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34754 14384
rect 34798 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34920 14384
rect 34920 14344 34922 14384
rect 34630 14302 34754 14344
rect 34798 14302 34922 14344
rect 49750 14384 49874 14426
rect 49918 14384 50042 14426
rect 49750 14344 49752 14384
rect 49752 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49874 14384
rect 49918 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50040 14384
rect 50040 14344 50042 14384
rect 49750 14302 49874 14344
rect 49918 14302 50042 14344
rect 64870 14384 64994 14426
rect 65038 14384 65162 14426
rect 64870 14344 64872 14384
rect 64872 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64994 14384
rect 65038 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65160 14384
rect 65160 14344 65162 14384
rect 64870 14302 64994 14344
rect 65038 14302 65162 14344
rect 79990 14384 80114 14426
rect 80158 14384 80282 14426
rect 79990 14344 79992 14384
rect 79992 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80114 14384
rect 80158 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80280 14384
rect 80280 14344 80282 14384
rect 79990 14302 80114 14344
rect 80158 14302 80282 14344
rect 95110 14384 95234 14426
rect 95278 14384 95402 14426
rect 95110 14344 95112 14384
rect 95112 14344 95154 14384
rect 95154 14344 95194 14384
rect 95194 14344 95234 14384
rect 95278 14344 95318 14384
rect 95318 14344 95358 14384
rect 95358 14344 95400 14384
rect 95400 14344 95402 14384
rect 95110 14302 95234 14344
rect 95278 14302 95402 14344
rect 3150 13628 3274 13670
rect 3318 13628 3442 13670
rect 3150 13588 3152 13628
rect 3152 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3274 13628
rect 3318 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3440 13628
rect 3440 13588 3442 13628
rect 3150 13546 3274 13588
rect 3318 13546 3442 13588
rect 18270 13628 18394 13670
rect 18438 13628 18562 13670
rect 18270 13588 18272 13628
rect 18272 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18394 13628
rect 18438 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18560 13628
rect 18560 13588 18562 13628
rect 18270 13546 18394 13588
rect 18438 13546 18562 13588
rect 33390 13628 33514 13670
rect 33558 13628 33682 13670
rect 33390 13588 33392 13628
rect 33392 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33514 13628
rect 33558 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33680 13628
rect 33680 13588 33682 13628
rect 33390 13546 33514 13588
rect 33558 13546 33682 13588
rect 48510 13628 48634 13670
rect 48678 13628 48802 13670
rect 48510 13588 48512 13628
rect 48512 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48634 13628
rect 48678 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48800 13628
rect 48800 13588 48802 13628
rect 48510 13546 48634 13588
rect 48678 13546 48802 13588
rect 63630 13628 63754 13670
rect 63798 13628 63922 13670
rect 63630 13588 63632 13628
rect 63632 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63754 13628
rect 63798 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63920 13628
rect 63920 13588 63922 13628
rect 63630 13546 63754 13588
rect 63798 13546 63922 13588
rect 78750 13628 78874 13670
rect 78918 13628 79042 13670
rect 78750 13588 78752 13628
rect 78752 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78874 13628
rect 78918 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79040 13628
rect 79040 13588 79042 13628
rect 78750 13546 78874 13588
rect 78918 13546 79042 13588
rect 93870 13628 93994 13670
rect 94038 13628 94162 13670
rect 93870 13588 93872 13628
rect 93872 13588 93914 13628
rect 93914 13588 93954 13628
rect 93954 13588 93994 13628
rect 94038 13588 94078 13628
rect 94078 13588 94118 13628
rect 94118 13588 94160 13628
rect 94160 13588 94162 13628
rect 93870 13546 93994 13588
rect 94038 13546 94162 13588
rect 4390 12872 4514 12914
rect 4558 12872 4682 12914
rect 4390 12832 4392 12872
rect 4392 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4514 12872
rect 4558 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4680 12872
rect 4680 12832 4682 12872
rect 4390 12790 4514 12832
rect 4558 12790 4682 12832
rect 19510 12872 19634 12914
rect 19678 12872 19802 12914
rect 19510 12832 19512 12872
rect 19512 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19634 12872
rect 19678 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19800 12872
rect 19800 12832 19802 12872
rect 19510 12790 19634 12832
rect 19678 12790 19802 12832
rect 34630 12872 34754 12914
rect 34798 12872 34922 12914
rect 34630 12832 34632 12872
rect 34632 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34754 12872
rect 34798 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34920 12872
rect 34920 12832 34922 12872
rect 34630 12790 34754 12832
rect 34798 12790 34922 12832
rect 49750 12872 49874 12914
rect 49918 12872 50042 12914
rect 49750 12832 49752 12872
rect 49752 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49874 12872
rect 49918 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50040 12872
rect 50040 12832 50042 12872
rect 49750 12790 49874 12832
rect 49918 12790 50042 12832
rect 64870 12872 64994 12914
rect 65038 12872 65162 12914
rect 64870 12832 64872 12872
rect 64872 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64994 12872
rect 65038 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65160 12872
rect 65160 12832 65162 12872
rect 64870 12790 64994 12832
rect 65038 12790 65162 12832
rect 79990 12872 80114 12914
rect 80158 12872 80282 12914
rect 79990 12832 79992 12872
rect 79992 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80114 12872
rect 80158 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80280 12872
rect 80280 12832 80282 12872
rect 79990 12790 80114 12832
rect 80158 12790 80282 12832
rect 95110 12872 95234 12914
rect 95278 12872 95402 12914
rect 95110 12832 95112 12872
rect 95112 12832 95154 12872
rect 95154 12832 95194 12872
rect 95194 12832 95234 12872
rect 95278 12832 95318 12872
rect 95318 12832 95358 12872
rect 95358 12832 95400 12872
rect 95400 12832 95402 12872
rect 95110 12790 95234 12832
rect 95278 12790 95402 12832
rect 3150 12116 3274 12158
rect 3318 12116 3442 12158
rect 3150 12076 3152 12116
rect 3152 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3274 12116
rect 3318 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3440 12116
rect 3440 12076 3442 12116
rect 3150 12034 3274 12076
rect 3318 12034 3442 12076
rect 18270 12116 18394 12158
rect 18438 12116 18562 12158
rect 18270 12076 18272 12116
rect 18272 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18394 12116
rect 18438 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18560 12116
rect 18560 12076 18562 12116
rect 18270 12034 18394 12076
rect 18438 12034 18562 12076
rect 33390 12116 33514 12158
rect 33558 12116 33682 12158
rect 33390 12076 33392 12116
rect 33392 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33514 12116
rect 33558 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33680 12116
rect 33680 12076 33682 12116
rect 33390 12034 33514 12076
rect 33558 12034 33682 12076
rect 48510 12116 48634 12158
rect 48678 12116 48802 12158
rect 48510 12076 48512 12116
rect 48512 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48634 12116
rect 48678 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48800 12116
rect 48800 12076 48802 12116
rect 48510 12034 48634 12076
rect 48678 12034 48802 12076
rect 63630 12116 63754 12158
rect 63798 12116 63922 12158
rect 63630 12076 63632 12116
rect 63632 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63754 12116
rect 63798 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63920 12116
rect 63920 12076 63922 12116
rect 63630 12034 63754 12076
rect 63798 12034 63922 12076
rect 78750 12116 78874 12158
rect 78918 12116 79042 12158
rect 78750 12076 78752 12116
rect 78752 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78874 12116
rect 78918 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79040 12116
rect 79040 12076 79042 12116
rect 78750 12034 78874 12076
rect 78918 12034 79042 12076
rect 93870 12116 93994 12158
rect 94038 12116 94162 12158
rect 93870 12076 93872 12116
rect 93872 12076 93914 12116
rect 93914 12076 93954 12116
rect 93954 12076 93994 12116
rect 94038 12076 94078 12116
rect 94078 12076 94118 12116
rect 94118 12076 94160 12116
rect 94160 12076 94162 12116
rect 93870 12034 93994 12076
rect 94038 12034 94162 12076
rect 4390 11360 4514 11402
rect 4558 11360 4682 11402
rect 4390 11320 4392 11360
rect 4392 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4514 11360
rect 4558 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4680 11360
rect 4680 11320 4682 11360
rect 4390 11278 4514 11320
rect 4558 11278 4682 11320
rect 19510 11360 19634 11402
rect 19678 11360 19802 11402
rect 19510 11320 19512 11360
rect 19512 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19634 11360
rect 19678 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19800 11360
rect 19800 11320 19802 11360
rect 19510 11278 19634 11320
rect 19678 11278 19802 11320
rect 34630 11360 34754 11402
rect 34798 11360 34922 11402
rect 34630 11320 34632 11360
rect 34632 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34754 11360
rect 34798 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34920 11360
rect 34920 11320 34922 11360
rect 34630 11278 34754 11320
rect 34798 11278 34922 11320
rect 49750 11360 49874 11402
rect 49918 11360 50042 11402
rect 49750 11320 49752 11360
rect 49752 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49874 11360
rect 49918 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50040 11360
rect 50040 11320 50042 11360
rect 49750 11278 49874 11320
rect 49918 11278 50042 11320
rect 64870 11360 64994 11402
rect 65038 11360 65162 11402
rect 64870 11320 64872 11360
rect 64872 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64994 11360
rect 65038 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65160 11360
rect 65160 11320 65162 11360
rect 64870 11278 64994 11320
rect 65038 11278 65162 11320
rect 79990 11360 80114 11402
rect 80158 11360 80282 11402
rect 79990 11320 79992 11360
rect 79992 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80114 11360
rect 80158 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80280 11360
rect 80280 11320 80282 11360
rect 79990 11278 80114 11320
rect 80158 11278 80282 11320
rect 95110 11360 95234 11402
rect 95278 11360 95402 11402
rect 95110 11320 95112 11360
rect 95112 11320 95154 11360
rect 95154 11320 95194 11360
rect 95194 11320 95234 11360
rect 95278 11320 95318 11360
rect 95318 11320 95358 11360
rect 95358 11320 95400 11360
rect 95400 11320 95402 11360
rect 95110 11278 95234 11320
rect 95278 11278 95402 11320
rect 3150 10604 3274 10646
rect 3318 10604 3442 10646
rect 3150 10564 3152 10604
rect 3152 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3274 10604
rect 3318 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3440 10604
rect 3440 10564 3442 10604
rect 3150 10522 3274 10564
rect 3318 10522 3442 10564
rect 18270 10604 18394 10646
rect 18438 10604 18562 10646
rect 18270 10564 18272 10604
rect 18272 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18394 10604
rect 18438 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18560 10604
rect 18560 10564 18562 10604
rect 18270 10522 18394 10564
rect 18438 10522 18562 10564
rect 33390 10604 33514 10646
rect 33558 10604 33682 10646
rect 33390 10564 33392 10604
rect 33392 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33514 10604
rect 33558 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33680 10604
rect 33680 10564 33682 10604
rect 33390 10522 33514 10564
rect 33558 10522 33682 10564
rect 48510 10604 48634 10646
rect 48678 10604 48802 10646
rect 48510 10564 48512 10604
rect 48512 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48634 10604
rect 48678 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48800 10604
rect 48800 10564 48802 10604
rect 48510 10522 48634 10564
rect 48678 10522 48802 10564
rect 63630 10604 63754 10646
rect 63798 10604 63922 10646
rect 63630 10564 63632 10604
rect 63632 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63754 10604
rect 63798 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63920 10604
rect 63920 10564 63922 10604
rect 63630 10522 63754 10564
rect 63798 10522 63922 10564
rect 78750 10604 78874 10646
rect 78918 10604 79042 10646
rect 78750 10564 78752 10604
rect 78752 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78874 10604
rect 78918 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79040 10604
rect 79040 10564 79042 10604
rect 78750 10522 78874 10564
rect 78918 10522 79042 10564
rect 93870 10604 93994 10646
rect 94038 10604 94162 10646
rect 93870 10564 93872 10604
rect 93872 10564 93914 10604
rect 93914 10564 93954 10604
rect 93954 10564 93994 10604
rect 94038 10564 94078 10604
rect 94078 10564 94118 10604
rect 94118 10564 94160 10604
rect 94160 10564 94162 10604
rect 93870 10522 93994 10564
rect 94038 10522 94162 10564
rect 4390 9848 4514 9890
rect 4558 9848 4682 9890
rect 4390 9808 4392 9848
rect 4392 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4514 9848
rect 4558 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4680 9848
rect 4680 9808 4682 9848
rect 4390 9766 4514 9808
rect 4558 9766 4682 9808
rect 19510 9848 19634 9890
rect 19678 9848 19802 9890
rect 19510 9808 19512 9848
rect 19512 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19634 9848
rect 19678 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19800 9848
rect 19800 9808 19802 9848
rect 19510 9766 19634 9808
rect 19678 9766 19802 9808
rect 34630 9848 34754 9890
rect 34798 9848 34922 9890
rect 34630 9808 34632 9848
rect 34632 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34754 9848
rect 34798 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34920 9848
rect 34920 9808 34922 9848
rect 34630 9766 34754 9808
rect 34798 9766 34922 9808
rect 49750 9848 49874 9890
rect 49918 9848 50042 9890
rect 49750 9808 49752 9848
rect 49752 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49874 9848
rect 49918 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50040 9848
rect 50040 9808 50042 9848
rect 49750 9766 49874 9808
rect 49918 9766 50042 9808
rect 64870 9848 64994 9890
rect 65038 9848 65162 9890
rect 64870 9808 64872 9848
rect 64872 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64994 9848
rect 65038 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65160 9848
rect 65160 9808 65162 9848
rect 64870 9766 64994 9808
rect 65038 9766 65162 9808
rect 79990 9848 80114 9890
rect 80158 9848 80282 9890
rect 79990 9808 79992 9848
rect 79992 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80114 9848
rect 80158 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80280 9848
rect 80280 9808 80282 9848
rect 79990 9766 80114 9808
rect 80158 9766 80282 9808
rect 95110 9848 95234 9890
rect 95278 9848 95402 9890
rect 95110 9808 95112 9848
rect 95112 9808 95154 9848
rect 95154 9808 95194 9848
rect 95194 9808 95234 9848
rect 95278 9808 95318 9848
rect 95318 9808 95358 9848
rect 95358 9808 95400 9848
rect 95400 9808 95402 9848
rect 95110 9766 95234 9808
rect 95278 9766 95402 9808
rect 3150 9092 3274 9134
rect 3318 9092 3442 9134
rect 3150 9052 3152 9092
rect 3152 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3274 9092
rect 3318 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3440 9092
rect 3440 9052 3442 9092
rect 3150 9010 3274 9052
rect 3318 9010 3442 9052
rect 18270 9092 18394 9134
rect 18438 9092 18562 9134
rect 18270 9052 18272 9092
rect 18272 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18394 9092
rect 18438 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18560 9092
rect 18560 9052 18562 9092
rect 18270 9010 18394 9052
rect 18438 9010 18562 9052
rect 33390 9092 33514 9134
rect 33558 9092 33682 9134
rect 33390 9052 33392 9092
rect 33392 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33514 9092
rect 33558 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33680 9092
rect 33680 9052 33682 9092
rect 33390 9010 33514 9052
rect 33558 9010 33682 9052
rect 48510 9092 48634 9134
rect 48678 9092 48802 9134
rect 48510 9052 48512 9092
rect 48512 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48634 9092
rect 48678 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48800 9092
rect 48800 9052 48802 9092
rect 48510 9010 48634 9052
rect 48678 9010 48802 9052
rect 63630 9092 63754 9134
rect 63798 9092 63922 9134
rect 63630 9052 63632 9092
rect 63632 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63754 9092
rect 63798 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63920 9092
rect 63920 9052 63922 9092
rect 63630 9010 63754 9052
rect 63798 9010 63922 9052
rect 78750 9092 78874 9134
rect 78918 9092 79042 9134
rect 78750 9052 78752 9092
rect 78752 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78874 9092
rect 78918 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79040 9092
rect 79040 9052 79042 9092
rect 78750 9010 78874 9052
rect 78918 9010 79042 9052
rect 93870 9092 93994 9134
rect 94038 9092 94162 9134
rect 93870 9052 93872 9092
rect 93872 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93994 9092
rect 94038 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94160 9092
rect 94160 9052 94162 9092
rect 93870 9010 93994 9052
rect 94038 9010 94162 9052
rect 4390 8336 4514 8378
rect 4558 8336 4682 8378
rect 4390 8296 4392 8336
rect 4392 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4514 8336
rect 4558 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4680 8336
rect 4680 8296 4682 8336
rect 4390 8254 4514 8296
rect 4558 8254 4682 8296
rect 19510 8336 19634 8378
rect 19678 8336 19802 8378
rect 19510 8296 19512 8336
rect 19512 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19634 8336
rect 19678 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19800 8336
rect 19800 8296 19802 8336
rect 19510 8254 19634 8296
rect 19678 8254 19802 8296
rect 34630 8336 34754 8378
rect 34798 8336 34922 8378
rect 34630 8296 34632 8336
rect 34632 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34754 8336
rect 34798 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34920 8336
rect 34920 8296 34922 8336
rect 34630 8254 34754 8296
rect 34798 8254 34922 8296
rect 49750 8336 49874 8378
rect 49918 8336 50042 8378
rect 49750 8296 49752 8336
rect 49752 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49874 8336
rect 49918 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50040 8336
rect 50040 8296 50042 8336
rect 49750 8254 49874 8296
rect 49918 8254 50042 8296
rect 64870 8336 64994 8378
rect 65038 8336 65162 8378
rect 64870 8296 64872 8336
rect 64872 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64994 8336
rect 65038 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65160 8336
rect 65160 8296 65162 8336
rect 64870 8254 64994 8296
rect 65038 8254 65162 8296
rect 79990 8336 80114 8378
rect 80158 8336 80282 8378
rect 79990 8296 79992 8336
rect 79992 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80114 8336
rect 80158 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80280 8336
rect 80280 8296 80282 8336
rect 79990 8254 80114 8296
rect 80158 8254 80282 8296
rect 95110 8336 95234 8378
rect 95278 8336 95402 8378
rect 95110 8296 95112 8336
rect 95112 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95234 8336
rect 95278 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95400 8336
rect 95400 8296 95402 8336
rect 95110 8254 95234 8296
rect 95278 8254 95402 8296
rect 3150 7580 3274 7622
rect 3318 7580 3442 7622
rect 3150 7540 3152 7580
rect 3152 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3274 7580
rect 3318 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3440 7580
rect 3440 7540 3442 7580
rect 3150 7498 3274 7540
rect 3318 7498 3442 7540
rect 18270 7580 18394 7622
rect 18438 7580 18562 7622
rect 18270 7540 18272 7580
rect 18272 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18394 7580
rect 18438 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18560 7580
rect 18560 7540 18562 7580
rect 18270 7498 18394 7540
rect 18438 7498 18562 7540
rect 33390 7580 33514 7622
rect 33558 7580 33682 7622
rect 33390 7540 33392 7580
rect 33392 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33514 7580
rect 33558 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33680 7580
rect 33680 7540 33682 7580
rect 33390 7498 33514 7540
rect 33558 7498 33682 7540
rect 48510 7580 48634 7622
rect 48678 7580 48802 7622
rect 48510 7540 48512 7580
rect 48512 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48634 7580
rect 48678 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48800 7580
rect 48800 7540 48802 7580
rect 48510 7498 48634 7540
rect 48678 7498 48802 7540
rect 63630 7580 63754 7622
rect 63798 7580 63922 7622
rect 63630 7540 63632 7580
rect 63632 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63754 7580
rect 63798 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63920 7580
rect 63920 7540 63922 7580
rect 63630 7498 63754 7540
rect 63798 7498 63922 7540
rect 78750 7580 78874 7622
rect 78918 7580 79042 7622
rect 78750 7540 78752 7580
rect 78752 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78874 7580
rect 78918 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79040 7580
rect 79040 7540 79042 7580
rect 78750 7498 78874 7540
rect 78918 7498 79042 7540
rect 93870 7580 93994 7622
rect 94038 7580 94162 7622
rect 93870 7540 93872 7580
rect 93872 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93994 7580
rect 94038 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94160 7580
rect 94160 7540 94162 7580
rect 93870 7498 93994 7540
rect 94038 7498 94162 7540
rect 4390 6824 4514 6866
rect 4558 6824 4682 6866
rect 4390 6784 4392 6824
rect 4392 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4514 6824
rect 4558 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4680 6824
rect 4680 6784 4682 6824
rect 4390 6742 4514 6784
rect 4558 6742 4682 6784
rect 19510 6824 19634 6866
rect 19678 6824 19802 6866
rect 19510 6784 19512 6824
rect 19512 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19634 6824
rect 19678 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19800 6824
rect 19800 6784 19802 6824
rect 19510 6742 19634 6784
rect 19678 6742 19802 6784
rect 34630 6824 34754 6866
rect 34798 6824 34922 6866
rect 34630 6784 34632 6824
rect 34632 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34754 6824
rect 34798 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34920 6824
rect 34920 6784 34922 6824
rect 34630 6742 34754 6784
rect 34798 6742 34922 6784
rect 49750 6824 49874 6866
rect 49918 6824 50042 6866
rect 49750 6784 49752 6824
rect 49752 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49874 6824
rect 49918 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50040 6824
rect 50040 6784 50042 6824
rect 49750 6742 49874 6784
rect 49918 6742 50042 6784
rect 64870 6824 64994 6866
rect 65038 6824 65162 6866
rect 64870 6784 64872 6824
rect 64872 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64994 6824
rect 65038 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65160 6824
rect 65160 6784 65162 6824
rect 64870 6742 64994 6784
rect 65038 6742 65162 6784
rect 79990 6824 80114 6866
rect 80158 6824 80282 6866
rect 79990 6784 79992 6824
rect 79992 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80114 6824
rect 80158 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80280 6824
rect 80280 6784 80282 6824
rect 79990 6742 80114 6784
rect 80158 6742 80282 6784
rect 95110 6824 95234 6866
rect 95278 6824 95402 6866
rect 95110 6784 95112 6824
rect 95112 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95234 6824
rect 95278 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95400 6824
rect 95400 6784 95402 6824
rect 95110 6742 95234 6784
rect 95278 6742 95402 6784
rect 3150 6068 3274 6110
rect 3318 6068 3442 6110
rect 3150 6028 3152 6068
rect 3152 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3274 6068
rect 3318 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3440 6068
rect 3440 6028 3442 6068
rect 3150 5986 3274 6028
rect 3318 5986 3442 6028
rect 18270 6068 18394 6110
rect 18438 6068 18562 6110
rect 18270 6028 18272 6068
rect 18272 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18394 6068
rect 18438 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18560 6068
rect 18560 6028 18562 6068
rect 18270 5986 18394 6028
rect 18438 5986 18562 6028
rect 33390 6068 33514 6110
rect 33558 6068 33682 6110
rect 33390 6028 33392 6068
rect 33392 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33514 6068
rect 33558 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33680 6068
rect 33680 6028 33682 6068
rect 33390 5986 33514 6028
rect 33558 5986 33682 6028
rect 48510 6068 48634 6110
rect 48678 6068 48802 6110
rect 48510 6028 48512 6068
rect 48512 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48634 6068
rect 48678 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48800 6068
rect 48800 6028 48802 6068
rect 48510 5986 48634 6028
rect 48678 5986 48802 6028
rect 63630 6068 63754 6110
rect 63798 6068 63922 6110
rect 63630 6028 63632 6068
rect 63632 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63754 6068
rect 63798 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63920 6068
rect 63920 6028 63922 6068
rect 63630 5986 63754 6028
rect 63798 5986 63922 6028
rect 78750 6068 78874 6110
rect 78918 6068 79042 6110
rect 78750 6028 78752 6068
rect 78752 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78874 6068
rect 78918 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79040 6068
rect 79040 6028 79042 6068
rect 78750 5986 78874 6028
rect 78918 5986 79042 6028
rect 93870 6068 93994 6110
rect 94038 6068 94162 6110
rect 93870 6028 93872 6068
rect 93872 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93994 6068
rect 94038 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94160 6068
rect 94160 6028 94162 6068
rect 93870 5986 93994 6028
rect 94038 5986 94162 6028
rect 4390 5312 4514 5354
rect 4558 5312 4682 5354
rect 4390 5272 4392 5312
rect 4392 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4514 5312
rect 4558 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4680 5312
rect 4680 5272 4682 5312
rect 4390 5230 4514 5272
rect 4558 5230 4682 5272
rect 19510 5312 19634 5354
rect 19678 5312 19802 5354
rect 19510 5272 19512 5312
rect 19512 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19634 5312
rect 19678 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19800 5312
rect 19800 5272 19802 5312
rect 19510 5230 19634 5272
rect 19678 5230 19802 5272
rect 34630 5312 34754 5354
rect 34798 5312 34922 5354
rect 34630 5272 34632 5312
rect 34632 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34754 5312
rect 34798 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34920 5312
rect 34920 5272 34922 5312
rect 34630 5230 34754 5272
rect 34798 5230 34922 5272
rect 49750 5312 49874 5354
rect 49918 5312 50042 5354
rect 49750 5272 49752 5312
rect 49752 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49874 5312
rect 49918 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50040 5312
rect 50040 5272 50042 5312
rect 49750 5230 49874 5272
rect 49918 5230 50042 5272
rect 64870 5312 64994 5354
rect 65038 5312 65162 5354
rect 64870 5272 64872 5312
rect 64872 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64994 5312
rect 65038 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65160 5312
rect 65160 5272 65162 5312
rect 64870 5230 64994 5272
rect 65038 5230 65162 5272
rect 79990 5312 80114 5354
rect 80158 5312 80282 5354
rect 79990 5272 79992 5312
rect 79992 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80114 5312
rect 80158 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80280 5312
rect 80280 5272 80282 5312
rect 79990 5230 80114 5272
rect 80158 5230 80282 5272
rect 95110 5312 95234 5354
rect 95278 5312 95402 5354
rect 95110 5272 95112 5312
rect 95112 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95234 5312
rect 95278 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95400 5312
rect 95400 5272 95402 5312
rect 95110 5230 95234 5272
rect 95278 5230 95402 5272
rect 3150 4556 3274 4598
rect 3318 4556 3442 4598
rect 3150 4516 3152 4556
rect 3152 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3274 4556
rect 3318 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3440 4556
rect 3440 4516 3442 4556
rect 3150 4474 3274 4516
rect 3318 4474 3442 4516
rect 18270 4556 18394 4598
rect 18438 4556 18562 4598
rect 18270 4516 18272 4556
rect 18272 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18394 4556
rect 18438 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18560 4556
rect 18560 4516 18562 4556
rect 18270 4474 18394 4516
rect 18438 4474 18562 4516
rect 33390 4556 33514 4598
rect 33558 4556 33682 4598
rect 33390 4516 33392 4556
rect 33392 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33514 4556
rect 33558 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33680 4556
rect 33680 4516 33682 4556
rect 33390 4474 33514 4516
rect 33558 4474 33682 4516
rect 48510 4556 48634 4598
rect 48678 4556 48802 4598
rect 48510 4516 48512 4556
rect 48512 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48634 4556
rect 48678 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48800 4556
rect 48800 4516 48802 4556
rect 48510 4474 48634 4516
rect 48678 4474 48802 4516
rect 63630 4556 63754 4598
rect 63798 4556 63922 4598
rect 63630 4516 63632 4556
rect 63632 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63754 4556
rect 63798 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63920 4556
rect 63920 4516 63922 4556
rect 63630 4474 63754 4516
rect 63798 4474 63922 4516
rect 78750 4556 78874 4598
rect 78918 4556 79042 4598
rect 78750 4516 78752 4556
rect 78752 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78874 4556
rect 78918 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79040 4556
rect 79040 4516 79042 4556
rect 78750 4474 78874 4516
rect 78918 4474 79042 4516
rect 93870 4556 93994 4598
rect 94038 4556 94162 4598
rect 93870 4516 93872 4556
rect 93872 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93994 4556
rect 94038 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94160 4556
rect 94160 4516 94162 4556
rect 93870 4474 93994 4516
rect 94038 4474 94162 4516
rect 4390 3800 4514 3842
rect 4558 3800 4682 3842
rect 4390 3760 4392 3800
rect 4392 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4514 3800
rect 4558 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4680 3800
rect 4680 3760 4682 3800
rect 4390 3718 4514 3760
rect 4558 3718 4682 3760
rect 19510 3800 19634 3842
rect 19678 3800 19802 3842
rect 19510 3760 19512 3800
rect 19512 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19634 3800
rect 19678 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19800 3800
rect 19800 3760 19802 3800
rect 19510 3718 19634 3760
rect 19678 3718 19802 3760
rect 34630 3800 34754 3842
rect 34798 3800 34922 3842
rect 34630 3760 34632 3800
rect 34632 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34754 3800
rect 34798 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34920 3800
rect 34920 3760 34922 3800
rect 34630 3718 34754 3760
rect 34798 3718 34922 3760
rect 49750 3800 49874 3842
rect 49918 3800 50042 3842
rect 49750 3760 49752 3800
rect 49752 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49874 3800
rect 49918 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50040 3800
rect 50040 3760 50042 3800
rect 49750 3718 49874 3760
rect 49918 3718 50042 3760
rect 64870 3800 64994 3842
rect 65038 3800 65162 3842
rect 64870 3760 64872 3800
rect 64872 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64994 3800
rect 65038 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65160 3800
rect 65160 3760 65162 3800
rect 64870 3718 64994 3760
rect 65038 3718 65162 3760
rect 79990 3800 80114 3842
rect 80158 3800 80282 3842
rect 79990 3760 79992 3800
rect 79992 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80114 3800
rect 80158 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80280 3800
rect 80280 3760 80282 3800
rect 79990 3718 80114 3760
rect 80158 3718 80282 3760
rect 95110 3800 95234 3842
rect 95278 3800 95402 3842
rect 95110 3760 95112 3800
rect 95112 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95234 3800
rect 95278 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95400 3800
rect 95400 3760 95402 3800
rect 95110 3718 95234 3760
rect 95278 3718 95402 3760
rect 3150 3044 3274 3086
rect 3318 3044 3442 3086
rect 3150 3004 3152 3044
rect 3152 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3274 3044
rect 3318 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3440 3044
rect 3440 3004 3442 3044
rect 3150 2962 3274 3004
rect 3318 2962 3442 3004
rect 18270 3044 18394 3086
rect 18438 3044 18562 3086
rect 18270 3004 18272 3044
rect 18272 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18394 3044
rect 18438 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18560 3044
rect 18560 3004 18562 3044
rect 18270 2962 18394 3004
rect 18438 2962 18562 3004
rect 33390 3044 33514 3086
rect 33558 3044 33682 3086
rect 33390 3004 33392 3044
rect 33392 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33514 3044
rect 33558 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33680 3044
rect 33680 3004 33682 3044
rect 33390 2962 33514 3004
rect 33558 2962 33682 3004
rect 48510 3044 48634 3086
rect 48678 3044 48802 3086
rect 48510 3004 48512 3044
rect 48512 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48634 3044
rect 48678 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48800 3044
rect 48800 3004 48802 3044
rect 48510 2962 48634 3004
rect 48678 2962 48802 3004
rect 63630 3044 63754 3086
rect 63798 3044 63922 3086
rect 63630 3004 63632 3044
rect 63632 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63754 3044
rect 63798 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63920 3044
rect 63920 3004 63922 3044
rect 63630 2962 63754 3004
rect 63798 2962 63922 3004
rect 78750 3044 78874 3086
rect 78918 3044 79042 3086
rect 78750 3004 78752 3044
rect 78752 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78874 3044
rect 78918 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79040 3044
rect 79040 3004 79042 3044
rect 78750 2962 78874 3004
rect 78918 2962 79042 3004
rect 93870 3044 93994 3086
rect 94038 3044 94162 3086
rect 93870 3004 93872 3044
rect 93872 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93994 3044
rect 94038 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94160 3044
rect 94160 3004 94162 3044
rect 93870 2962 93994 3004
rect 94038 2962 94162 3004
rect 4390 2288 4514 2330
rect 4558 2288 4682 2330
rect 4390 2248 4392 2288
rect 4392 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4514 2288
rect 4558 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4680 2288
rect 4680 2248 4682 2288
rect 4390 2206 4514 2248
rect 4558 2206 4682 2248
rect 19510 2288 19634 2330
rect 19678 2288 19802 2330
rect 19510 2248 19512 2288
rect 19512 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19634 2288
rect 19678 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19800 2288
rect 19800 2248 19802 2288
rect 19510 2206 19634 2248
rect 19678 2206 19802 2248
rect 34630 2288 34754 2330
rect 34798 2288 34922 2330
rect 34630 2248 34632 2288
rect 34632 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34754 2288
rect 34798 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34920 2288
rect 34920 2248 34922 2288
rect 34630 2206 34754 2248
rect 34798 2206 34922 2248
rect 49750 2288 49874 2330
rect 49918 2288 50042 2330
rect 49750 2248 49752 2288
rect 49752 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49874 2288
rect 49918 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50040 2288
rect 50040 2248 50042 2288
rect 49750 2206 49874 2248
rect 49918 2206 50042 2248
rect 64870 2288 64994 2330
rect 65038 2288 65162 2330
rect 64870 2248 64872 2288
rect 64872 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64994 2288
rect 65038 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65160 2288
rect 65160 2248 65162 2288
rect 64870 2206 64994 2248
rect 65038 2206 65162 2248
rect 79990 2288 80114 2330
rect 80158 2288 80282 2330
rect 79990 2248 79992 2288
rect 79992 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80114 2288
rect 80158 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80280 2288
rect 80280 2248 80282 2288
rect 79990 2206 80114 2248
rect 80158 2206 80282 2248
rect 95110 2288 95234 2330
rect 95278 2288 95402 2330
rect 95110 2248 95112 2288
rect 95112 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95234 2288
rect 95278 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95400 2288
rect 95400 2248 95402 2288
rect 95110 2206 95234 2248
rect 95278 2206 95402 2248
rect 3150 1532 3274 1574
rect 3318 1532 3442 1574
rect 3150 1492 3152 1532
rect 3152 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3274 1532
rect 3318 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3440 1532
rect 3440 1492 3442 1532
rect 3150 1450 3274 1492
rect 3318 1450 3442 1492
rect 18270 1532 18394 1574
rect 18438 1532 18562 1574
rect 18270 1492 18272 1532
rect 18272 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18394 1532
rect 18438 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18560 1532
rect 18560 1492 18562 1532
rect 18270 1450 18394 1492
rect 18438 1450 18562 1492
rect 33390 1532 33514 1574
rect 33558 1532 33682 1574
rect 33390 1492 33392 1532
rect 33392 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33514 1532
rect 33558 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33680 1532
rect 33680 1492 33682 1532
rect 33390 1450 33514 1492
rect 33558 1450 33682 1492
rect 48510 1532 48634 1574
rect 48678 1532 48802 1574
rect 48510 1492 48512 1532
rect 48512 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48634 1532
rect 48678 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48800 1532
rect 48800 1492 48802 1532
rect 48510 1450 48634 1492
rect 48678 1450 48802 1492
rect 63630 1532 63754 1574
rect 63798 1532 63922 1574
rect 63630 1492 63632 1532
rect 63632 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63754 1532
rect 63798 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63920 1532
rect 63920 1492 63922 1532
rect 63630 1450 63754 1492
rect 63798 1450 63922 1492
rect 78750 1532 78874 1574
rect 78918 1532 79042 1574
rect 78750 1492 78752 1532
rect 78752 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78874 1532
rect 78918 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79040 1532
rect 79040 1492 79042 1532
rect 78750 1450 78874 1492
rect 78918 1450 79042 1492
rect 93870 1532 93994 1574
rect 94038 1532 94162 1574
rect 93870 1492 93872 1532
rect 93872 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93994 1532
rect 94038 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94160 1532
rect 94160 1492 94162 1532
rect 93870 1450 93994 1492
rect 94038 1450 94162 1492
rect 4390 776 4514 818
rect 4558 776 4682 818
rect 4390 736 4392 776
rect 4392 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4514 776
rect 4558 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4680 776
rect 4680 736 4682 776
rect 4390 694 4514 736
rect 4558 694 4682 736
rect 19510 776 19634 818
rect 19678 776 19802 818
rect 19510 736 19512 776
rect 19512 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19634 776
rect 19678 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19800 776
rect 19800 736 19802 776
rect 19510 694 19634 736
rect 19678 694 19802 736
rect 34630 776 34754 818
rect 34798 776 34922 818
rect 34630 736 34632 776
rect 34632 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34754 776
rect 34798 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34920 776
rect 34920 736 34922 776
rect 34630 694 34754 736
rect 34798 694 34922 736
rect 49750 776 49874 818
rect 49918 776 50042 818
rect 49750 736 49752 776
rect 49752 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49874 776
rect 49918 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50040 776
rect 50040 736 50042 776
rect 49750 694 49874 736
rect 49918 694 50042 736
rect 64870 776 64994 818
rect 65038 776 65162 818
rect 64870 736 64872 776
rect 64872 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64994 776
rect 65038 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65160 776
rect 65160 736 65162 776
rect 64870 694 64994 736
rect 65038 694 65162 736
rect 79990 776 80114 818
rect 80158 776 80282 818
rect 79990 736 79992 776
rect 79992 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80114 776
rect 80158 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80280 776
rect 80280 736 80282 776
rect 79990 694 80114 736
rect 80158 694 80282 736
rect 95110 776 95234 818
rect 95278 776 95402 818
rect 95110 736 95112 776
rect 95112 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95234 776
rect 95278 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95400 776
rect 95400 736 95402 776
rect 95110 694 95234 736
rect 95278 694 95402 736
<< metal6 >>
rect 4316 38618 4756 38682
rect 3076 37862 3516 38600
rect 3076 37738 3150 37862
rect 3274 37738 3318 37862
rect 3442 37738 3516 37862
rect 3076 36350 3516 37738
rect 3076 36226 3150 36350
rect 3274 36226 3318 36350
rect 3442 36226 3516 36350
rect 3076 34838 3516 36226
rect 3076 34714 3150 34838
rect 3274 34714 3318 34838
rect 3442 34714 3516 34838
rect 3076 33326 3516 34714
rect 3076 33202 3150 33326
rect 3274 33202 3318 33326
rect 3442 33202 3516 33326
rect 3076 31814 3516 33202
rect 3076 31690 3150 31814
rect 3274 31690 3318 31814
rect 3442 31690 3516 31814
rect 3076 30302 3516 31690
rect 3076 30178 3150 30302
rect 3274 30178 3318 30302
rect 3442 30178 3516 30302
rect 3076 28790 3516 30178
rect 3076 28666 3150 28790
rect 3274 28666 3318 28790
rect 3442 28666 3516 28790
rect 3076 27278 3516 28666
rect 3076 27154 3150 27278
rect 3274 27154 3318 27278
rect 3442 27154 3516 27278
rect 3076 25766 3516 27154
rect 3076 25642 3150 25766
rect 3274 25642 3318 25766
rect 3442 25642 3516 25766
rect 3076 24254 3516 25642
rect 3076 24130 3150 24254
rect 3274 24130 3318 24254
rect 3442 24130 3516 24254
rect 3076 22742 3516 24130
rect 3076 22618 3150 22742
rect 3274 22618 3318 22742
rect 3442 22618 3516 22742
rect 3076 21230 3516 22618
rect 3076 21106 3150 21230
rect 3274 21106 3318 21230
rect 3442 21106 3516 21230
rect 3076 19718 3516 21106
rect 3076 19594 3150 19718
rect 3274 19594 3318 19718
rect 3442 19594 3516 19718
rect 3076 18206 3516 19594
rect 3076 18082 3150 18206
rect 3274 18082 3318 18206
rect 3442 18082 3516 18206
rect 3076 16694 3516 18082
rect 3076 16570 3150 16694
rect 3274 16570 3318 16694
rect 3442 16570 3516 16694
rect 3076 15182 3516 16570
rect 3076 15058 3150 15182
rect 3274 15058 3318 15182
rect 3442 15058 3516 15182
rect 3076 13670 3516 15058
rect 3076 13546 3150 13670
rect 3274 13546 3318 13670
rect 3442 13546 3516 13670
rect 3076 12158 3516 13546
rect 3076 12034 3150 12158
rect 3274 12034 3318 12158
rect 3442 12034 3516 12158
rect 3076 10646 3516 12034
rect 3076 10522 3150 10646
rect 3274 10522 3318 10646
rect 3442 10522 3516 10646
rect 3076 9134 3516 10522
rect 3076 9010 3150 9134
rect 3274 9010 3318 9134
rect 3442 9010 3516 9134
rect 3076 7622 3516 9010
rect 3076 7498 3150 7622
rect 3274 7498 3318 7622
rect 3442 7498 3516 7622
rect 3076 6110 3516 7498
rect 3076 5986 3150 6110
rect 3274 5986 3318 6110
rect 3442 5986 3516 6110
rect 3076 4598 3516 5986
rect 3076 4474 3150 4598
rect 3274 4474 3318 4598
rect 3442 4474 3516 4598
rect 3076 3086 3516 4474
rect 3076 2962 3150 3086
rect 3274 2962 3318 3086
rect 3442 2962 3516 3086
rect 3076 1574 3516 2962
rect 3076 1450 3150 1574
rect 3274 1450 3318 1574
rect 3442 1450 3516 1574
rect 3076 712 3516 1450
rect 4316 38494 4390 38618
rect 4514 38494 4558 38618
rect 4682 38494 4756 38618
rect 19436 38618 19876 38682
rect 4316 37106 4756 38494
rect 4316 36982 4390 37106
rect 4514 36982 4558 37106
rect 4682 36982 4756 37106
rect 4316 35594 4756 36982
rect 4316 35470 4390 35594
rect 4514 35470 4558 35594
rect 4682 35470 4756 35594
rect 4316 34082 4756 35470
rect 4316 33958 4390 34082
rect 4514 33958 4558 34082
rect 4682 33958 4756 34082
rect 4316 32570 4756 33958
rect 4316 32446 4390 32570
rect 4514 32446 4558 32570
rect 4682 32446 4756 32570
rect 4316 31058 4756 32446
rect 4316 30934 4390 31058
rect 4514 30934 4558 31058
rect 4682 30934 4756 31058
rect 4316 29546 4756 30934
rect 4316 29422 4390 29546
rect 4514 29422 4558 29546
rect 4682 29422 4756 29546
rect 4316 28034 4756 29422
rect 4316 27910 4390 28034
rect 4514 27910 4558 28034
rect 4682 27910 4756 28034
rect 4316 26522 4756 27910
rect 4316 26398 4390 26522
rect 4514 26398 4558 26522
rect 4682 26398 4756 26522
rect 4316 25010 4756 26398
rect 4316 24886 4390 25010
rect 4514 24886 4558 25010
rect 4682 24886 4756 25010
rect 4316 23498 4756 24886
rect 4316 23374 4390 23498
rect 4514 23374 4558 23498
rect 4682 23374 4756 23498
rect 4316 21986 4756 23374
rect 4316 21862 4390 21986
rect 4514 21862 4558 21986
rect 4682 21862 4756 21986
rect 4316 20474 4756 21862
rect 4316 20350 4390 20474
rect 4514 20350 4558 20474
rect 4682 20350 4756 20474
rect 4316 18962 4756 20350
rect 4316 18838 4390 18962
rect 4514 18838 4558 18962
rect 4682 18838 4756 18962
rect 4316 17450 4756 18838
rect 4316 17326 4390 17450
rect 4514 17326 4558 17450
rect 4682 17326 4756 17450
rect 4316 15938 4756 17326
rect 4316 15814 4390 15938
rect 4514 15814 4558 15938
rect 4682 15814 4756 15938
rect 4316 14426 4756 15814
rect 4316 14302 4390 14426
rect 4514 14302 4558 14426
rect 4682 14302 4756 14426
rect 4316 12914 4756 14302
rect 4316 12790 4390 12914
rect 4514 12790 4558 12914
rect 4682 12790 4756 12914
rect 4316 11402 4756 12790
rect 4316 11278 4390 11402
rect 4514 11278 4558 11402
rect 4682 11278 4756 11402
rect 4316 9890 4756 11278
rect 4316 9766 4390 9890
rect 4514 9766 4558 9890
rect 4682 9766 4756 9890
rect 4316 8378 4756 9766
rect 4316 8254 4390 8378
rect 4514 8254 4558 8378
rect 4682 8254 4756 8378
rect 4316 6866 4756 8254
rect 4316 6742 4390 6866
rect 4514 6742 4558 6866
rect 4682 6742 4756 6866
rect 4316 5354 4756 6742
rect 4316 5230 4390 5354
rect 4514 5230 4558 5354
rect 4682 5230 4756 5354
rect 4316 3842 4756 5230
rect 4316 3718 4390 3842
rect 4514 3718 4558 3842
rect 4682 3718 4756 3842
rect 4316 2330 4756 3718
rect 4316 2206 4390 2330
rect 4514 2206 4558 2330
rect 4682 2206 4756 2330
rect 4316 818 4756 2206
rect 4316 694 4390 818
rect 4514 694 4558 818
rect 4682 694 4756 818
rect 18196 37862 18636 38600
rect 18196 37738 18270 37862
rect 18394 37738 18438 37862
rect 18562 37738 18636 37862
rect 18196 36350 18636 37738
rect 18196 36226 18270 36350
rect 18394 36226 18438 36350
rect 18562 36226 18636 36350
rect 18196 34838 18636 36226
rect 18196 34714 18270 34838
rect 18394 34714 18438 34838
rect 18562 34714 18636 34838
rect 18196 33326 18636 34714
rect 18196 33202 18270 33326
rect 18394 33202 18438 33326
rect 18562 33202 18636 33326
rect 18196 31814 18636 33202
rect 18196 31690 18270 31814
rect 18394 31690 18438 31814
rect 18562 31690 18636 31814
rect 18196 30302 18636 31690
rect 18196 30178 18270 30302
rect 18394 30178 18438 30302
rect 18562 30178 18636 30302
rect 18196 28790 18636 30178
rect 18196 28666 18270 28790
rect 18394 28666 18438 28790
rect 18562 28666 18636 28790
rect 18196 27278 18636 28666
rect 18196 27154 18270 27278
rect 18394 27154 18438 27278
rect 18562 27154 18636 27278
rect 18196 25766 18636 27154
rect 18196 25642 18270 25766
rect 18394 25642 18438 25766
rect 18562 25642 18636 25766
rect 18196 24254 18636 25642
rect 18196 24130 18270 24254
rect 18394 24130 18438 24254
rect 18562 24130 18636 24254
rect 18196 22742 18636 24130
rect 18196 22618 18270 22742
rect 18394 22618 18438 22742
rect 18562 22618 18636 22742
rect 18196 21230 18636 22618
rect 18196 21106 18270 21230
rect 18394 21106 18438 21230
rect 18562 21106 18636 21230
rect 18196 19718 18636 21106
rect 18196 19594 18270 19718
rect 18394 19594 18438 19718
rect 18562 19594 18636 19718
rect 18196 18206 18636 19594
rect 18196 18082 18270 18206
rect 18394 18082 18438 18206
rect 18562 18082 18636 18206
rect 18196 16694 18636 18082
rect 18196 16570 18270 16694
rect 18394 16570 18438 16694
rect 18562 16570 18636 16694
rect 18196 15182 18636 16570
rect 18196 15058 18270 15182
rect 18394 15058 18438 15182
rect 18562 15058 18636 15182
rect 18196 13670 18636 15058
rect 18196 13546 18270 13670
rect 18394 13546 18438 13670
rect 18562 13546 18636 13670
rect 18196 12158 18636 13546
rect 18196 12034 18270 12158
rect 18394 12034 18438 12158
rect 18562 12034 18636 12158
rect 18196 10646 18636 12034
rect 18196 10522 18270 10646
rect 18394 10522 18438 10646
rect 18562 10522 18636 10646
rect 18196 9134 18636 10522
rect 18196 9010 18270 9134
rect 18394 9010 18438 9134
rect 18562 9010 18636 9134
rect 18196 7622 18636 9010
rect 18196 7498 18270 7622
rect 18394 7498 18438 7622
rect 18562 7498 18636 7622
rect 18196 6110 18636 7498
rect 18196 5986 18270 6110
rect 18394 5986 18438 6110
rect 18562 5986 18636 6110
rect 18196 4598 18636 5986
rect 18196 4474 18270 4598
rect 18394 4474 18438 4598
rect 18562 4474 18636 4598
rect 18196 3086 18636 4474
rect 18196 2962 18270 3086
rect 18394 2962 18438 3086
rect 18562 2962 18636 3086
rect 18196 1574 18636 2962
rect 18196 1450 18270 1574
rect 18394 1450 18438 1574
rect 18562 1450 18636 1574
rect 18196 712 18636 1450
rect 19436 38494 19510 38618
rect 19634 38494 19678 38618
rect 19802 38494 19876 38618
rect 34556 38618 34996 38682
rect 19436 37106 19876 38494
rect 19436 36982 19510 37106
rect 19634 36982 19678 37106
rect 19802 36982 19876 37106
rect 19436 35594 19876 36982
rect 19436 35470 19510 35594
rect 19634 35470 19678 35594
rect 19802 35470 19876 35594
rect 19436 34082 19876 35470
rect 19436 33958 19510 34082
rect 19634 33958 19678 34082
rect 19802 33958 19876 34082
rect 19436 32570 19876 33958
rect 19436 32446 19510 32570
rect 19634 32446 19678 32570
rect 19802 32446 19876 32570
rect 19436 31058 19876 32446
rect 19436 30934 19510 31058
rect 19634 30934 19678 31058
rect 19802 30934 19876 31058
rect 19436 29546 19876 30934
rect 19436 29422 19510 29546
rect 19634 29422 19678 29546
rect 19802 29422 19876 29546
rect 19436 28034 19876 29422
rect 19436 27910 19510 28034
rect 19634 27910 19678 28034
rect 19802 27910 19876 28034
rect 19436 26522 19876 27910
rect 19436 26398 19510 26522
rect 19634 26398 19678 26522
rect 19802 26398 19876 26522
rect 19436 25010 19876 26398
rect 19436 24886 19510 25010
rect 19634 24886 19678 25010
rect 19802 24886 19876 25010
rect 19436 23498 19876 24886
rect 19436 23374 19510 23498
rect 19634 23374 19678 23498
rect 19802 23374 19876 23498
rect 19436 21986 19876 23374
rect 19436 21862 19510 21986
rect 19634 21862 19678 21986
rect 19802 21862 19876 21986
rect 19436 20474 19876 21862
rect 19436 20350 19510 20474
rect 19634 20350 19678 20474
rect 19802 20350 19876 20474
rect 19436 18962 19876 20350
rect 19436 18838 19510 18962
rect 19634 18838 19678 18962
rect 19802 18838 19876 18962
rect 19436 17450 19876 18838
rect 19436 17326 19510 17450
rect 19634 17326 19678 17450
rect 19802 17326 19876 17450
rect 19436 15938 19876 17326
rect 19436 15814 19510 15938
rect 19634 15814 19678 15938
rect 19802 15814 19876 15938
rect 19436 14426 19876 15814
rect 19436 14302 19510 14426
rect 19634 14302 19678 14426
rect 19802 14302 19876 14426
rect 19436 12914 19876 14302
rect 19436 12790 19510 12914
rect 19634 12790 19678 12914
rect 19802 12790 19876 12914
rect 19436 11402 19876 12790
rect 19436 11278 19510 11402
rect 19634 11278 19678 11402
rect 19802 11278 19876 11402
rect 19436 9890 19876 11278
rect 19436 9766 19510 9890
rect 19634 9766 19678 9890
rect 19802 9766 19876 9890
rect 19436 8378 19876 9766
rect 19436 8254 19510 8378
rect 19634 8254 19678 8378
rect 19802 8254 19876 8378
rect 19436 6866 19876 8254
rect 19436 6742 19510 6866
rect 19634 6742 19678 6866
rect 19802 6742 19876 6866
rect 19436 5354 19876 6742
rect 19436 5230 19510 5354
rect 19634 5230 19678 5354
rect 19802 5230 19876 5354
rect 19436 3842 19876 5230
rect 19436 3718 19510 3842
rect 19634 3718 19678 3842
rect 19802 3718 19876 3842
rect 19436 2330 19876 3718
rect 19436 2206 19510 2330
rect 19634 2206 19678 2330
rect 19802 2206 19876 2330
rect 19436 818 19876 2206
rect 4316 630 4756 694
rect 19436 694 19510 818
rect 19634 694 19678 818
rect 19802 694 19876 818
rect 33316 37862 33756 38600
rect 33316 37738 33390 37862
rect 33514 37738 33558 37862
rect 33682 37738 33756 37862
rect 33316 36350 33756 37738
rect 33316 36226 33390 36350
rect 33514 36226 33558 36350
rect 33682 36226 33756 36350
rect 33316 34838 33756 36226
rect 33316 34714 33390 34838
rect 33514 34714 33558 34838
rect 33682 34714 33756 34838
rect 33316 33326 33756 34714
rect 33316 33202 33390 33326
rect 33514 33202 33558 33326
rect 33682 33202 33756 33326
rect 33316 31814 33756 33202
rect 33316 31690 33390 31814
rect 33514 31690 33558 31814
rect 33682 31690 33756 31814
rect 33316 30302 33756 31690
rect 33316 30178 33390 30302
rect 33514 30178 33558 30302
rect 33682 30178 33756 30302
rect 33316 28790 33756 30178
rect 33316 28666 33390 28790
rect 33514 28666 33558 28790
rect 33682 28666 33756 28790
rect 33316 27278 33756 28666
rect 33316 27154 33390 27278
rect 33514 27154 33558 27278
rect 33682 27154 33756 27278
rect 33316 25766 33756 27154
rect 33316 25642 33390 25766
rect 33514 25642 33558 25766
rect 33682 25642 33756 25766
rect 33316 24254 33756 25642
rect 33316 24130 33390 24254
rect 33514 24130 33558 24254
rect 33682 24130 33756 24254
rect 33316 22742 33756 24130
rect 33316 22618 33390 22742
rect 33514 22618 33558 22742
rect 33682 22618 33756 22742
rect 33316 21230 33756 22618
rect 33316 21106 33390 21230
rect 33514 21106 33558 21230
rect 33682 21106 33756 21230
rect 33316 19718 33756 21106
rect 33316 19594 33390 19718
rect 33514 19594 33558 19718
rect 33682 19594 33756 19718
rect 33316 18206 33756 19594
rect 33316 18082 33390 18206
rect 33514 18082 33558 18206
rect 33682 18082 33756 18206
rect 33316 16694 33756 18082
rect 33316 16570 33390 16694
rect 33514 16570 33558 16694
rect 33682 16570 33756 16694
rect 33316 15182 33756 16570
rect 33316 15058 33390 15182
rect 33514 15058 33558 15182
rect 33682 15058 33756 15182
rect 33316 13670 33756 15058
rect 33316 13546 33390 13670
rect 33514 13546 33558 13670
rect 33682 13546 33756 13670
rect 33316 12158 33756 13546
rect 33316 12034 33390 12158
rect 33514 12034 33558 12158
rect 33682 12034 33756 12158
rect 33316 10646 33756 12034
rect 33316 10522 33390 10646
rect 33514 10522 33558 10646
rect 33682 10522 33756 10646
rect 33316 9134 33756 10522
rect 33316 9010 33390 9134
rect 33514 9010 33558 9134
rect 33682 9010 33756 9134
rect 33316 7622 33756 9010
rect 33316 7498 33390 7622
rect 33514 7498 33558 7622
rect 33682 7498 33756 7622
rect 33316 6110 33756 7498
rect 33316 5986 33390 6110
rect 33514 5986 33558 6110
rect 33682 5986 33756 6110
rect 33316 4598 33756 5986
rect 33316 4474 33390 4598
rect 33514 4474 33558 4598
rect 33682 4474 33756 4598
rect 33316 3086 33756 4474
rect 33316 2962 33390 3086
rect 33514 2962 33558 3086
rect 33682 2962 33756 3086
rect 33316 1574 33756 2962
rect 33316 1450 33390 1574
rect 33514 1450 33558 1574
rect 33682 1450 33756 1574
rect 33316 712 33756 1450
rect 34556 38494 34630 38618
rect 34754 38494 34798 38618
rect 34922 38494 34996 38618
rect 49676 38618 50116 38682
rect 34556 37106 34996 38494
rect 34556 36982 34630 37106
rect 34754 36982 34798 37106
rect 34922 36982 34996 37106
rect 34556 35594 34996 36982
rect 34556 35470 34630 35594
rect 34754 35470 34798 35594
rect 34922 35470 34996 35594
rect 34556 34082 34996 35470
rect 34556 33958 34630 34082
rect 34754 33958 34798 34082
rect 34922 33958 34996 34082
rect 34556 32570 34996 33958
rect 34556 32446 34630 32570
rect 34754 32446 34798 32570
rect 34922 32446 34996 32570
rect 34556 31058 34996 32446
rect 34556 30934 34630 31058
rect 34754 30934 34798 31058
rect 34922 30934 34996 31058
rect 34556 29546 34996 30934
rect 34556 29422 34630 29546
rect 34754 29422 34798 29546
rect 34922 29422 34996 29546
rect 34556 28034 34996 29422
rect 34556 27910 34630 28034
rect 34754 27910 34798 28034
rect 34922 27910 34996 28034
rect 34556 26522 34996 27910
rect 34556 26398 34630 26522
rect 34754 26398 34798 26522
rect 34922 26398 34996 26522
rect 34556 25010 34996 26398
rect 34556 24886 34630 25010
rect 34754 24886 34798 25010
rect 34922 24886 34996 25010
rect 34556 23498 34996 24886
rect 34556 23374 34630 23498
rect 34754 23374 34798 23498
rect 34922 23374 34996 23498
rect 34556 21986 34996 23374
rect 34556 21862 34630 21986
rect 34754 21862 34798 21986
rect 34922 21862 34996 21986
rect 34556 20474 34996 21862
rect 34556 20350 34630 20474
rect 34754 20350 34798 20474
rect 34922 20350 34996 20474
rect 34556 18962 34996 20350
rect 34556 18838 34630 18962
rect 34754 18838 34798 18962
rect 34922 18838 34996 18962
rect 34556 17450 34996 18838
rect 34556 17326 34630 17450
rect 34754 17326 34798 17450
rect 34922 17326 34996 17450
rect 34556 15938 34996 17326
rect 34556 15814 34630 15938
rect 34754 15814 34798 15938
rect 34922 15814 34996 15938
rect 34556 14426 34996 15814
rect 34556 14302 34630 14426
rect 34754 14302 34798 14426
rect 34922 14302 34996 14426
rect 34556 12914 34996 14302
rect 34556 12790 34630 12914
rect 34754 12790 34798 12914
rect 34922 12790 34996 12914
rect 34556 11402 34996 12790
rect 34556 11278 34630 11402
rect 34754 11278 34798 11402
rect 34922 11278 34996 11402
rect 34556 9890 34996 11278
rect 34556 9766 34630 9890
rect 34754 9766 34798 9890
rect 34922 9766 34996 9890
rect 34556 8378 34996 9766
rect 34556 8254 34630 8378
rect 34754 8254 34798 8378
rect 34922 8254 34996 8378
rect 34556 6866 34996 8254
rect 34556 6742 34630 6866
rect 34754 6742 34798 6866
rect 34922 6742 34996 6866
rect 34556 5354 34996 6742
rect 34556 5230 34630 5354
rect 34754 5230 34798 5354
rect 34922 5230 34996 5354
rect 34556 3842 34996 5230
rect 34556 3718 34630 3842
rect 34754 3718 34798 3842
rect 34922 3718 34996 3842
rect 34556 2330 34996 3718
rect 34556 2206 34630 2330
rect 34754 2206 34798 2330
rect 34922 2206 34996 2330
rect 34556 818 34996 2206
rect 19436 630 19876 694
rect 34556 694 34630 818
rect 34754 694 34798 818
rect 34922 694 34996 818
rect 48436 37862 48876 38600
rect 48436 37738 48510 37862
rect 48634 37738 48678 37862
rect 48802 37738 48876 37862
rect 48436 36350 48876 37738
rect 48436 36226 48510 36350
rect 48634 36226 48678 36350
rect 48802 36226 48876 36350
rect 48436 34838 48876 36226
rect 48436 34714 48510 34838
rect 48634 34714 48678 34838
rect 48802 34714 48876 34838
rect 48436 33326 48876 34714
rect 48436 33202 48510 33326
rect 48634 33202 48678 33326
rect 48802 33202 48876 33326
rect 48436 31814 48876 33202
rect 48436 31690 48510 31814
rect 48634 31690 48678 31814
rect 48802 31690 48876 31814
rect 48436 30302 48876 31690
rect 48436 30178 48510 30302
rect 48634 30178 48678 30302
rect 48802 30178 48876 30302
rect 48436 28790 48876 30178
rect 48436 28666 48510 28790
rect 48634 28666 48678 28790
rect 48802 28666 48876 28790
rect 48436 27278 48876 28666
rect 48436 27154 48510 27278
rect 48634 27154 48678 27278
rect 48802 27154 48876 27278
rect 48436 25766 48876 27154
rect 48436 25642 48510 25766
rect 48634 25642 48678 25766
rect 48802 25642 48876 25766
rect 48436 24254 48876 25642
rect 48436 24130 48510 24254
rect 48634 24130 48678 24254
rect 48802 24130 48876 24254
rect 48436 22742 48876 24130
rect 48436 22618 48510 22742
rect 48634 22618 48678 22742
rect 48802 22618 48876 22742
rect 48436 21230 48876 22618
rect 48436 21106 48510 21230
rect 48634 21106 48678 21230
rect 48802 21106 48876 21230
rect 48436 19718 48876 21106
rect 48436 19594 48510 19718
rect 48634 19594 48678 19718
rect 48802 19594 48876 19718
rect 48436 18206 48876 19594
rect 48436 18082 48510 18206
rect 48634 18082 48678 18206
rect 48802 18082 48876 18206
rect 48436 16694 48876 18082
rect 48436 16570 48510 16694
rect 48634 16570 48678 16694
rect 48802 16570 48876 16694
rect 48436 15182 48876 16570
rect 48436 15058 48510 15182
rect 48634 15058 48678 15182
rect 48802 15058 48876 15182
rect 48436 13670 48876 15058
rect 48436 13546 48510 13670
rect 48634 13546 48678 13670
rect 48802 13546 48876 13670
rect 48436 12158 48876 13546
rect 48436 12034 48510 12158
rect 48634 12034 48678 12158
rect 48802 12034 48876 12158
rect 48436 10646 48876 12034
rect 48436 10522 48510 10646
rect 48634 10522 48678 10646
rect 48802 10522 48876 10646
rect 48436 9134 48876 10522
rect 48436 9010 48510 9134
rect 48634 9010 48678 9134
rect 48802 9010 48876 9134
rect 48436 7622 48876 9010
rect 48436 7498 48510 7622
rect 48634 7498 48678 7622
rect 48802 7498 48876 7622
rect 48436 6110 48876 7498
rect 48436 5986 48510 6110
rect 48634 5986 48678 6110
rect 48802 5986 48876 6110
rect 48436 4598 48876 5986
rect 48436 4474 48510 4598
rect 48634 4474 48678 4598
rect 48802 4474 48876 4598
rect 48436 3086 48876 4474
rect 48436 2962 48510 3086
rect 48634 2962 48678 3086
rect 48802 2962 48876 3086
rect 48436 1574 48876 2962
rect 48436 1450 48510 1574
rect 48634 1450 48678 1574
rect 48802 1450 48876 1574
rect 48436 712 48876 1450
rect 49676 38494 49750 38618
rect 49874 38494 49918 38618
rect 50042 38494 50116 38618
rect 64796 38618 65236 38682
rect 49676 37106 50116 38494
rect 49676 36982 49750 37106
rect 49874 36982 49918 37106
rect 50042 36982 50116 37106
rect 49676 35594 50116 36982
rect 49676 35470 49750 35594
rect 49874 35470 49918 35594
rect 50042 35470 50116 35594
rect 49676 34082 50116 35470
rect 49676 33958 49750 34082
rect 49874 33958 49918 34082
rect 50042 33958 50116 34082
rect 49676 32570 50116 33958
rect 49676 32446 49750 32570
rect 49874 32446 49918 32570
rect 50042 32446 50116 32570
rect 49676 31058 50116 32446
rect 49676 30934 49750 31058
rect 49874 30934 49918 31058
rect 50042 30934 50116 31058
rect 49676 29546 50116 30934
rect 49676 29422 49750 29546
rect 49874 29422 49918 29546
rect 50042 29422 50116 29546
rect 49676 28034 50116 29422
rect 49676 27910 49750 28034
rect 49874 27910 49918 28034
rect 50042 27910 50116 28034
rect 49676 26522 50116 27910
rect 49676 26398 49750 26522
rect 49874 26398 49918 26522
rect 50042 26398 50116 26522
rect 49676 25010 50116 26398
rect 49676 24886 49750 25010
rect 49874 24886 49918 25010
rect 50042 24886 50116 25010
rect 49676 23498 50116 24886
rect 49676 23374 49750 23498
rect 49874 23374 49918 23498
rect 50042 23374 50116 23498
rect 49676 21986 50116 23374
rect 49676 21862 49750 21986
rect 49874 21862 49918 21986
rect 50042 21862 50116 21986
rect 49676 20474 50116 21862
rect 49676 20350 49750 20474
rect 49874 20350 49918 20474
rect 50042 20350 50116 20474
rect 49676 18962 50116 20350
rect 49676 18838 49750 18962
rect 49874 18838 49918 18962
rect 50042 18838 50116 18962
rect 49676 17450 50116 18838
rect 49676 17326 49750 17450
rect 49874 17326 49918 17450
rect 50042 17326 50116 17450
rect 49676 15938 50116 17326
rect 49676 15814 49750 15938
rect 49874 15814 49918 15938
rect 50042 15814 50116 15938
rect 49676 14426 50116 15814
rect 49676 14302 49750 14426
rect 49874 14302 49918 14426
rect 50042 14302 50116 14426
rect 49676 12914 50116 14302
rect 49676 12790 49750 12914
rect 49874 12790 49918 12914
rect 50042 12790 50116 12914
rect 49676 11402 50116 12790
rect 49676 11278 49750 11402
rect 49874 11278 49918 11402
rect 50042 11278 50116 11402
rect 49676 9890 50116 11278
rect 49676 9766 49750 9890
rect 49874 9766 49918 9890
rect 50042 9766 50116 9890
rect 49676 8378 50116 9766
rect 49676 8254 49750 8378
rect 49874 8254 49918 8378
rect 50042 8254 50116 8378
rect 49676 6866 50116 8254
rect 49676 6742 49750 6866
rect 49874 6742 49918 6866
rect 50042 6742 50116 6866
rect 49676 5354 50116 6742
rect 49676 5230 49750 5354
rect 49874 5230 49918 5354
rect 50042 5230 50116 5354
rect 49676 3842 50116 5230
rect 49676 3718 49750 3842
rect 49874 3718 49918 3842
rect 50042 3718 50116 3842
rect 49676 2330 50116 3718
rect 49676 2206 49750 2330
rect 49874 2206 49918 2330
rect 50042 2206 50116 2330
rect 49676 818 50116 2206
rect 34556 630 34996 694
rect 49676 694 49750 818
rect 49874 694 49918 818
rect 50042 694 50116 818
rect 63556 37862 63996 38600
rect 63556 37738 63630 37862
rect 63754 37738 63798 37862
rect 63922 37738 63996 37862
rect 63556 36350 63996 37738
rect 63556 36226 63630 36350
rect 63754 36226 63798 36350
rect 63922 36226 63996 36350
rect 63556 34838 63996 36226
rect 63556 34714 63630 34838
rect 63754 34714 63798 34838
rect 63922 34714 63996 34838
rect 63556 33326 63996 34714
rect 63556 33202 63630 33326
rect 63754 33202 63798 33326
rect 63922 33202 63996 33326
rect 63556 31814 63996 33202
rect 63556 31690 63630 31814
rect 63754 31690 63798 31814
rect 63922 31690 63996 31814
rect 63556 30302 63996 31690
rect 63556 30178 63630 30302
rect 63754 30178 63798 30302
rect 63922 30178 63996 30302
rect 63556 28790 63996 30178
rect 63556 28666 63630 28790
rect 63754 28666 63798 28790
rect 63922 28666 63996 28790
rect 63556 27278 63996 28666
rect 63556 27154 63630 27278
rect 63754 27154 63798 27278
rect 63922 27154 63996 27278
rect 63556 25766 63996 27154
rect 63556 25642 63630 25766
rect 63754 25642 63798 25766
rect 63922 25642 63996 25766
rect 63556 24254 63996 25642
rect 63556 24130 63630 24254
rect 63754 24130 63798 24254
rect 63922 24130 63996 24254
rect 63556 22742 63996 24130
rect 63556 22618 63630 22742
rect 63754 22618 63798 22742
rect 63922 22618 63996 22742
rect 63556 21230 63996 22618
rect 63556 21106 63630 21230
rect 63754 21106 63798 21230
rect 63922 21106 63996 21230
rect 63556 19718 63996 21106
rect 63556 19594 63630 19718
rect 63754 19594 63798 19718
rect 63922 19594 63996 19718
rect 63556 18206 63996 19594
rect 63556 18082 63630 18206
rect 63754 18082 63798 18206
rect 63922 18082 63996 18206
rect 63556 16694 63996 18082
rect 63556 16570 63630 16694
rect 63754 16570 63798 16694
rect 63922 16570 63996 16694
rect 63556 15182 63996 16570
rect 63556 15058 63630 15182
rect 63754 15058 63798 15182
rect 63922 15058 63996 15182
rect 63556 13670 63996 15058
rect 63556 13546 63630 13670
rect 63754 13546 63798 13670
rect 63922 13546 63996 13670
rect 63556 12158 63996 13546
rect 63556 12034 63630 12158
rect 63754 12034 63798 12158
rect 63922 12034 63996 12158
rect 63556 10646 63996 12034
rect 63556 10522 63630 10646
rect 63754 10522 63798 10646
rect 63922 10522 63996 10646
rect 63556 9134 63996 10522
rect 63556 9010 63630 9134
rect 63754 9010 63798 9134
rect 63922 9010 63996 9134
rect 63556 7622 63996 9010
rect 63556 7498 63630 7622
rect 63754 7498 63798 7622
rect 63922 7498 63996 7622
rect 63556 6110 63996 7498
rect 63556 5986 63630 6110
rect 63754 5986 63798 6110
rect 63922 5986 63996 6110
rect 63556 4598 63996 5986
rect 63556 4474 63630 4598
rect 63754 4474 63798 4598
rect 63922 4474 63996 4598
rect 63556 3086 63996 4474
rect 63556 2962 63630 3086
rect 63754 2962 63798 3086
rect 63922 2962 63996 3086
rect 63556 1574 63996 2962
rect 63556 1450 63630 1574
rect 63754 1450 63798 1574
rect 63922 1450 63996 1574
rect 63556 712 63996 1450
rect 64796 38494 64870 38618
rect 64994 38494 65038 38618
rect 65162 38494 65236 38618
rect 79916 38618 80356 38682
rect 64796 37106 65236 38494
rect 64796 36982 64870 37106
rect 64994 36982 65038 37106
rect 65162 36982 65236 37106
rect 64796 35594 65236 36982
rect 64796 35470 64870 35594
rect 64994 35470 65038 35594
rect 65162 35470 65236 35594
rect 64796 34082 65236 35470
rect 64796 33958 64870 34082
rect 64994 33958 65038 34082
rect 65162 33958 65236 34082
rect 64796 32570 65236 33958
rect 64796 32446 64870 32570
rect 64994 32446 65038 32570
rect 65162 32446 65236 32570
rect 64796 31058 65236 32446
rect 64796 30934 64870 31058
rect 64994 30934 65038 31058
rect 65162 30934 65236 31058
rect 64796 29546 65236 30934
rect 64796 29422 64870 29546
rect 64994 29422 65038 29546
rect 65162 29422 65236 29546
rect 64796 28034 65236 29422
rect 64796 27910 64870 28034
rect 64994 27910 65038 28034
rect 65162 27910 65236 28034
rect 64796 26522 65236 27910
rect 64796 26398 64870 26522
rect 64994 26398 65038 26522
rect 65162 26398 65236 26522
rect 64796 25010 65236 26398
rect 64796 24886 64870 25010
rect 64994 24886 65038 25010
rect 65162 24886 65236 25010
rect 64796 23498 65236 24886
rect 64796 23374 64870 23498
rect 64994 23374 65038 23498
rect 65162 23374 65236 23498
rect 64796 21986 65236 23374
rect 64796 21862 64870 21986
rect 64994 21862 65038 21986
rect 65162 21862 65236 21986
rect 64796 20474 65236 21862
rect 64796 20350 64870 20474
rect 64994 20350 65038 20474
rect 65162 20350 65236 20474
rect 64796 18962 65236 20350
rect 64796 18838 64870 18962
rect 64994 18838 65038 18962
rect 65162 18838 65236 18962
rect 64796 17450 65236 18838
rect 64796 17326 64870 17450
rect 64994 17326 65038 17450
rect 65162 17326 65236 17450
rect 64796 15938 65236 17326
rect 64796 15814 64870 15938
rect 64994 15814 65038 15938
rect 65162 15814 65236 15938
rect 64796 14426 65236 15814
rect 64796 14302 64870 14426
rect 64994 14302 65038 14426
rect 65162 14302 65236 14426
rect 64796 12914 65236 14302
rect 64796 12790 64870 12914
rect 64994 12790 65038 12914
rect 65162 12790 65236 12914
rect 64796 11402 65236 12790
rect 64796 11278 64870 11402
rect 64994 11278 65038 11402
rect 65162 11278 65236 11402
rect 64796 9890 65236 11278
rect 64796 9766 64870 9890
rect 64994 9766 65038 9890
rect 65162 9766 65236 9890
rect 64796 8378 65236 9766
rect 64796 8254 64870 8378
rect 64994 8254 65038 8378
rect 65162 8254 65236 8378
rect 64796 6866 65236 8254
rect 64796 6742 64870 6866
rect 64994 6742 65038 6866
rect 65162 6742 65236 6866
rect 64796 5354 65236 6742
rect 64796 5230 64870 5354
rect 64994 5230 65038 5354
rect 65162 5230 65236 5354
rect 64796 3842 65236 5230
rect 64796 3718 64870 3842
rect 64994 3718 65038 3842
rect 65162 3718 65236 3842
rect 64796 2330 65236 3718
rect 64796 2206 64870 2330
rect 64994 2206 65038 2330
rect 65162 2206 65236 2330
rect 64796 818 65236 2206
rect 49676 630 50116 694
rect 64796 694 64870 818
rect 64994 694 65038 818
rect 65162 694 65236 818
rect 78676 37862 79116 38600
rect 78676 37738 78750 37862
rect 78874 37738 78918 37862
rect 79042 37738 79116 37862
rect 78676 36350 79116 37738
rect 78676 36226 78750 36350
rect 78874 36226 78918 36350
rect 79042 36226 79116 36350
rect 78676 34838 79116 36226
rect 78676 34714 78750 34838
rect 78874 34714 78918 34838
rect 79042 34714 79116 34838
rect 78676 33326 79116 34714
rect 78676 33202 78750 33326
rect 78874 33202 78918 33326
rect 79042 33202 79116 33326
rect 78676 31814 79116 33202
rect 78676 31690 78750 31814
rect 78874 31690 78918 31814
rect 79042 31690 79116 31814
rect 78676 30302 79116 31690
rect 78676 30178 78750 30302
rect 78874 30178 78918 30302
rect 79042 30178 79116 30302
rect 78676 28790 79116 30178
rect 78676 28666 78750 28790
rect 78874 28666 78918 28790
rect 79042 28666 79116 28790
rect 78676 27278 79116 28666
rect 78676 27154 78750 27278
rect 78874 27154 78918 27278
rect 79042 27154 79116 27278
rect 78676 25766 79116 27154
rect 78676 25642 78750 25766
rect 78874 25642 78918 25766
rect 79042 25642 79116 25766
rect 78676 24254 79116 25642
rect 78676 24130 78750 24254
rect 78874 24130 78918 24254
rect 79042 24130 79116 24254
rect 78676 22742 79116 24130
rect 78676 22618 78750 22742
rect 78874 22618 78918 22742
rect 79042 22618 79116 22742
rect 78676 21230 79116 22618
rect 78676 21106 78750 21230
rect 78874 21106 78918 21230
rect 79042 21106 79116 21230
rect 78676 19718 79116 21106
rect 78676 19594 78750 19718
rect 78874 19594 78918 19718
rect 79042 19594 79116 19718
rect 78676 18206 79116 19594
rect 78676 18082 78750 18206
rect 78874 18082 78918 18206
rect 79042 18082 79116 18206
rect 78676 16694 79116 18082
rect 78676 16570 78750 16694
rect 78874 16570 78918 16694
rect 79042 16570 79116 16694
rect 78676 15182 79116 16570
rect 78676 15058 78750 15182
rect 78874 15058 78918 15182
rect 79042 15058 79116 15182
rect 78676 13670 79116 15058
rect 78676 13546 78750 13670
rect 78874 13546 78918 13670
rect 79042 13546 79116 13670
rect 78676 12158 79116 13546
rect 78676 12034 78750 12158
rect 78874 12034 78918 12158
rect 79042 12034 79116 12158
rect 78676 10646 79116 12034
rect 78676 10522 78750 10646
rect 78874 10522 78918 10646
rect 79042 10522 79116 10646
rect 78676 9134 79116 10522
rect 78676 9010 78750 9134
rect 78874 9010 78918 9134
rect 79042 9010 79116 9134
rect 78676 7622 79116 9010
rect 78676 7498 78750 7622
rect 78874 7498 78918 7622
rect 79042 7498 79116 7622
rect 78676 6110 79116 7498
rect 78676 5986 78750 6110
rect 78874 5986 78918 6110
rect 79042 5986 79116 6110
rect 78676 4598 79116 5986
rect 78676 4474 78750 4598
rect 78874 4474 78918 4598
rect 79042 4474 79116 4598
rect 78676 3086 79116 4474
rect 78676 2962 78750 3086
rect 78874 2962 78918 3086
rect 79042 2962 79116 3086
rect 78676 1574 79116 2962
rect 78676 1450 78750 1574
rect 78874 1450 78918 1574
rect 79042 1450 79116 1574
rect 78676 712 79116 1450
rect 79916 38494 79990 38618
rect 80114 38494 80158 38618
rect 80282 38494 80356 38618
rect 95036 38618 95476 38682
rect 79916 37106 80356 38494
rect 79916 36982 79990 37106
rect 80114 36982 80158 37106
rect 80282 36982 80356 37106
rect 79916 35594 80356 36982
rect 79916 35470 79990 35594
rect 80114 35470 80158 35594
rect 80282 35470 80356 35594
rect 79916 34082 80356 35470
rect 79916 33958 79990 34082
rect 80114 33958 80158 34082
rect 80282 33958 80356 34082
rect 79916 32570 80356 33958
rect 79916 32446 79990 32570
rect 80114 32446 80158 32570
rect 80282 32446 80356 32570
rect 79916 31058 80356 32446
rect 79916 30934 79990 31058
rect 80114 30934 80158 31058
rect 80282 30934 80356 31058
rect 79916 29546 80356 30934
rect 79916 29422 79990 29546
rect 80114 29422 80158 29546
rect 80282 29422 80356 29546
rect 79916 28034 80356 29422
rect 79916 27910 79990 28034
rect 80114 27910 80158 28034
rect 80282 27910 80356 28034
rect 79916 26522 80356 27910
rect 79916 26398 79990 26522
rect 80114 26398 80158 26522
rect 80282 26398 80356 26522
rect 79916 25010 80356 26398
rect 79916 24886 79990 25010
rect 80114 24886 80158 25010
rect 80282 24886 80356 25010
rect 79916 23498 80356 24886
rect 79916 23374 79990 23498
rect 80114 23374 80158 23498
rect 80282 23374 80356 23498
rect 79916 21986 80356 23374
rect 79916 21862 79990 21986
rect 80114 21862 80158 21986
rect 80282 21862 80356 21986
rect 79916 20474 80356 21862
rect 79916 20350 79990 20474
rect 80114 20350 80158 20474
rect 80282 20350 80356 20474
rect 79916 18962 80356 20350
rect 79916 18838 79990 18962
rect 80114 18838 80158 18962
rect 80282 18838 80356 18962
rect 79916 17450 80356 18838
rect 79916 17326 79990 17450
rect 80114 17326 80158 17450
rect 80282 17326 80356 17450
rect 79916 15938 80356 17326
rect 79916 15814 79990 15938
rect 80114 15814 80158 15938
rect 80282 15814 80356 15938
rect 79916 14426 80356 15814
rect 79916 14302 79990 14426
rect 80114 14302 80158 14426
rect 80282 14302 80356 14426
rect 79916 12914 80356 14302
rect 79916 12790 79990 12914
rect 80114 12790 80158 12914
rect 80282 12790 80356 12914
rect 79916 11402 80356 12790
rect 79916 11278 79990 11402
rect 80114 11278 80158 11402
rect 80282 11278 80356 11402
rect 79916 9890 80356 11278
rect 79916 9766 79990 9890
rect 80114 9766 80158 9890
rect 80282 9766 80356 9890
rect 79916 8378 80356 9766
rect 79916 8254 79990 8378
rect 80114 8254 80158 8378
rect 80282 8254 80356 8378
rect 79916 6866 80356 8254
rect 79916 6742 79990 6866
rect 80114 6742 80158 6866
rect 80282 6742 80356 6866
rect 79916 5354 80356 6742
rect 79916 5230 79990 5354
rect 80114 5230 80158 5354
rect 80282 5230 80356 5354
rect 79916 3842 80356 5230
rect 79916 3718 79990 3842
rect 80114 3718 80158 3842
rect 80282 3718 80356 3842
rect 79916 2330 80356 3718
rect 79916 2206 79990 2330
rect 80114 2206 80158 2330
rect 80282 2206 80356 2330
rect 79916 818 80356 2206
rect 64796 630 65236 694
rect 79916 694 79990 818
rect 80114 694 80158 818
rect 80282 694 80356 818
rect 93796 37862 94236 38600
rect 93796 37738 93870 37862
rect 93994 37738 94038 37862
rect 94162 37738 94236 37862
rect 93796 36350 94236 37738
rect 93796 36226 93870 36350
rect 93994 36226 94038 36350
rect 94162 36226 94236 36350
rect 93796 34838 94236 36226
rect 93796 34714 93870 34838
rect 93994 34714 94038 34838
rect 94162 34714 94236 34838
rect 93796 33326 94236 34714
rect 93796 33202 93870 33326
rect 93994 33202 94038 33326
rect 94162 33202 94236 33326
rect 93796 31814 94236 33202
rect 93796 31690 93870 31814
rect 93994 31690 94038 31814
rect 94162 31690 94236 31814
rect 93796 30302 94236 31690
rect 93796 30178 93870 30302
rect 93994 30178 94038 30302
rect 94162 30178 94236 30302
rect 93796 28790 94236 30178
rect 93796 28666 93870 28790
rect 93994 28666 94038 28790
rect 94162 28666 94236 28790
rect 93796 27278 94236 28666
rect 93796 27154 93870 27278
rect 93994 27154 94038 27278
rect 94162 27154 94236 27278
rect 93796 25766 94236 27154
rect 93796 25642 93870 25766
rect 93994 25642 94038 25766
rect 94162 25642 94236 25766
rect 93796 24254 94236 25642
rect 93796 24130 93870 24254
rect 93994 24130 94038 24254
rect 94162 24130 94236 24254
rect 93796 22742 94236 24130
rect 93796 22618 93870 22742
rect 93994 22618 94038 22742
rect 94162 22618 94236 22742
rect 93796 21230 94236 22618
rect 93796 21106 93870 21230
rect 93994 21106 94038 21230
rect 94162 21106 94236 21230
rect 93796 19718 94236 21106
rect 93796 19594 93870 19718
rect 93994 19594 94038 19718
rect 94162 19594 94236 19718
rect 93796 18206 94236 19594
rect 93796 18082 93870 18206
rect 93994 18082 94038 18206
rect 94162 18082 94236 18206
rect 93796 16694 94236 18082
rect 93796 16570 93870 16694
rect 93994 16570 94038 16694
rect 94162 16570 94236 16694
rect 93796 15182 94236 16570
rect 93796 15058 93870 15182
rect 93994 15058 94038 15182
rect 94162 15058 94236 15182
rect 93796 13670 94236 15058
rect 93796 13546 93870 13670
rect 93994 13546 94038 13670
rect 94162 13546 94236 13670
rect 93796 12158 94236 13546
rect 93796 12034 93870 12158
rect 93994 12034 94038 12158
rect 94162 12034 94236 12158
rect 93796 10646 94236 12034
rect 93796 10522 93870 10646
rect 93994 10522 94038 10646
rect 94162 10522 94236 10646
rect 93796 9134 94236 10522
rect 93796 9010 93870 9134
rect 93994 9010 94038 9134
rect 94162 9010 94236 9134
rect 93796 7622 94236 9010
rect 93796 7498 93870 7622
rect 93994 7498 94038 7622
rect 94162 7498 94236 7622
rect 93796 6110 94236 7498
rect 93796 5986 93870 6110
rect 93994 5986 94038 6110
rect 94162 5986 94236 6110
rect 93796 4598 94236 5986
rect 93796 4474 93870 4598
rect 93994 4474 94038 4598
rect 94162 4474 94236 4598
rect 93796 3086 94236 4474
rect 93796 2962 93870 3086
rect 93994 2962 94038 3086
rect 94162 2962 94236 3086
rect 93796 1574 94236 2962
rect 93796 1450 93870 1574
rect 93994 1450 94038 1574
rect 94162 1450 94236 1574
rect 93796 712 94236 1450
rect 95036 38494 95110 38618
rect 95234 38494 95278 38618
rect 95402 38494 95476 38618
rect 95036 37106 95476 38494
rect 95036 36982 95110 37106
rect 95234 36982 95278 37106
rect 95402 36982 95476 37106
rect 95036 35594 95476 36982
rect 95036 35470 95110 35594
rect 95234 35470 95278 35594
rect 95402 35470 95476 35594
rect 95036 34082 95476 35470
rect 95036 33958 95110 34082
rect 95234 33958 95278 34082
rect 95402 33958 95476 34082
rect 95036 32570 95476 33958
rect 95036 32446 95110 32570
rect 95234 32446 95278 32570
rect 95402 32446 95476 32570
rect 95036 31058 95476 32446
rect 95036 30934 95110 31058
rect 95234 30934 95278 31058
rect 95402 30934 95476 31058
rect 95036 29546 95476 30934
rect 95036 29422 95110 29546
rect 95234 29422 95278 29546
rect 95402 29422 95476 29546
rect 95036 28034 95476 29422
rect 95036 27910 95110 28034
rect 95234 27910 95278 28034
rect 95402 27910 95476 28034
rect 95036 26522 95476 27910
rect 95036 26398 95110 26522
rect 95234 26398 95278 26522
rect 95402 26398 95476 26522
rect 95036 25010 95476 26398
rect 95036 24886 95110 25010
rect 95234 24886 95278 25010
rect 95402 24886 95476 25010
rect 95036 23498 95476 24886
rect 95036 23374 95110 23498
rect 95234 23374 95278 23498
rect 95402 23374 95476 23498
rect 95036 21986 95476 23374
rect 95036 21862 95110 21986
rect 95234 21862 95278 21986
rect 95402 21862 95476 21986
rect 95036 20474 95476 21862
rect 95036 20350 95110 20474
rect 95234 20350 95278 20474
rect 95402 20350 95476 20474
rect 95036 18962 95476 20350
rect 95036 18838 95110 18962
rect 95234 18838 95278 18962
rect 95402 18838 95476 18962
rect 95036 17450 95476 18838
rect 95036 17326 95110 17450
rect 95234 17326 95278 17450
rect 95402 17326 95476 17450
rect 95036 15938 95476 17326
rect 95036 15814 95110 15938
rect 95234 15814 95278 15938
rect 95402 15814 95476 15938
rect 95036 14426 95476 15814
rect 95036 14302 95110 14426
rect 95234 14302 95278 14426
rect 95402 14302 95476 14426
rect 95036 12914 95476 14302
rect 95036 12790 95110 12914
rect 95234 12790 95278 12914
rect 95402 12790 95476 12914
rect 95036 11402 95476 12790
rect 95036 11278 95110 11402
rect 95234 11278 95278 11402
rect 95402 11278 95476 11402
rect 95036 9890 95476 11278
rect 95036 9766 95110 9890
rect 95234 9766 95278 9890
rect 95402 9766 95476 9890
rect 95036 8378 95476 9766
rect 95036 8254 95110 8378
rect 95234 8254 95278 8378
rect 95402 8254 95476 8378
rect 95036 6866 95476 8254
rect 95036 6742 95110 6866
rect 95234 6742 95278 6866
rect 95402 6742 95476 6866
rect 95036 5354 95476 6742
rect 95036 5230 95110 5354
rect 95234 5230 95278 5354
rect 95402 5230 95476 5354
rect 95036 3842 95476 5230
rect 95036 3718 95110 3842
rect 95234 3718 95278 3842
rect 95402 3718 95476 3842
rect 95036 2330 95476 3718
rect 95036 2206 95110 2330
rect 95234 2206 95278 2330
rect 95402 2206 95476 2330
rect 95036 818 95476 2206
rect 79916 630 80356 694
rect 95036 694 95110 818
rect 95234 694 95278 818
rect 95402 694 95476 818
rect 95036 630 95476 694
use sg13g2_inv_1  _31_
timestamp 1676386529
transform 1 0 8352 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _32_
timestamp 1676386529
transform 1 0 4032 0 -1 9828
box -48 -56 336 834
use sg13g2_and3_1  _33_
timestamp 1676975269
transform 1 0 2688 0 1 11340
box -48 -56 720 834
use sg13g2_and3_1  _34_
timestamp 1676975269
transform 1 0 6816 0 1 8316
box -48 -56 720 834
use sg13g2_and2_1  _35_
timestamp 1676905363
transform 1 0 9120 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _36_
timestamp 1685182643
transform -1 0 10560 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _37_
timestamp 1683980220
transform -1 0 11520 0 -1 14364
box -48 -56 528 834
use sg13g2_a21oi_1  _38_
timestamp 1683980220
transform -1 0 10080 0 1 11340
box -48 -56 528 834
use sg13g2_and4_1  _39_
timestamp 1676989577
transform -1 0 9216 0 1 11340
box -48 -56 816 834
use sg13g2_nor3_1  _40_
timestamp 1676643042
transform 1 0 9600 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _41_
timestamp 1685182643
transform -1 0 9312 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _42_
timestamp 1683980220
transform 1 0 8352 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _43_
timestamp 1685182643
transform 1 0 2496 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _44_
timestamp 1683980220
transform 1 0 3168 0 1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _45_
timestamp 1683980220
transform -1 0 2688 0 1 11340
box -48 -56 528 834
use sg13g2_nor3_1  _46_
timestamp 1676643042
transform -1 0 4704 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _47_
timestamp 1685182643
transform -1 0 9600 0 -1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _48_
timestamp 1683980220
transform 1 0 9216 0 1 3780
box -48 -56 528 834
use sg13g2_a21oi_1  _49_
timestamp 1683980220
transform -1 0 4224 0 -1 5292
box -48 -56 528 834
use sg13g2_nand3_1  _50_
timestamp 1683995554
transform 1 0 5184 0 1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _51_
timestamp 1676560849
transform -1 0 5088 0 -1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _52_
timestamp 1676630787
transform 1 0 4224 0 -1 5292
box -48 -56 432 834
use sg13g2_a221oi_1  _53_
timestamp 1685204697
transform 1 0 8640 0 -1 8316
box -48 -56 816 834
use sg13g2_tiehi  _54__26
timestamp 1680007851
transform -1 0 13920 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _54_
timestamp 1746542328
transform 1 0 13056 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _55_
timestamp 1746542328
transform 1 0 14016 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _55__25
timestamp 1680007851
transform -1 0 14880 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _56_
timestamp 1746542328
transform 1 0 7584 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _56__23
timestamp 1680007851
transform 1 0 7680 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  _57__21
timestamp 1680007851
transform 1 0 5088 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _57_
timestamp 1746542328
transform 1 0 4896 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _58_
timestamp 1746542328
transform -1 0 5280 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _58__19
timestamp 1680007851
transform 1 0 3744 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _59_
timestamp 1746542328
transform 1 0 9120 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _59__24
timestamp 1680007851
transform -1 0 9984 0 1 2268
box -48 -56 432 834
use sg13g2_tiehi  _60__20
timestamp 1680007851
transform -1 0 4416 0 -1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _60_
timestamp 1746542328
transform 1 0 3552 0 1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _61__22
timestamp 1680007851
transform -1 0 12576 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _61_
timestamp 1746542328
transform 1 0 11616 0 1 6804
box -48 -56 2640 834
use sg13g2_buf_1  _78_
timestamp 1676385511
transform -1 0 2976 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _79_
timestamp 1676385511
transform -1 0 2976 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _80_
timestamp 1676385511
transform -1 0 2976 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _81_
timestamp 1676385511
transform -1 0 2976 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _82_
timestamp 1676385511
transform -1 0 2976 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _83_
timestamp 1676385511
transform -1 0 2592 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _84_
timestamp 1676385511
transform -1 0 2976 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _85_
timestamp 1676385511
transform -1 0 2976 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_16  clkbuf_0_clk
timestamp 1676557096
transform -1 0 12096 0 -1 12852
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_0__f_clk
timestamp 1676557096
transform -1 0 12672 0 -1 9828
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_1__f_clk
timestamp 1676557096
transform 1 0 8832 0 -1 15876
box -48 -56 2448 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679585382
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679585382
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679585382
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679585382
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679585382
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679585382
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679585382
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679585382
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679585382
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679585382
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679585382
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679585382
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679585382
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679585382
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679585382
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679585382
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679585382
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679585382
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679585382
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679585382
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679585382
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679585382
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679585382
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679585382
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679585382
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679585382
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679585382
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679585382
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679585382
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679585382
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679585382
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679585382
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679585382
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679585382
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679585382
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679585382
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679585382
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679585382
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679585382
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679585382
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679585382
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679585382
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679585382
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679585382
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679585382
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679585382
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679585382
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679585382
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679585382
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679585382
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679585382
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679585382
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679585382
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679585382
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679585382
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679585382
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679585382
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679585382
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679585382
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679585382
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679585382
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679585382
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679585382
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679585382
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679585382
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679585382
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679585382
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679585382
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679585382
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679585382
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679585382
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679585382
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679585382
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679585382
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679585382
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679585382
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679585382
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679585382
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679585382
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679585382
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679585382
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679585382
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679585382
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679585382
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679585382
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679585382
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679585382
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679585382
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679585382
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679585382
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679585382
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679585382
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679585382
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679585382
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679585382
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679585382
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679585382
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679585382
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679585382
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679585382
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679585382
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679585382
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679585382
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679585382
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679585382
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679585382
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679585382
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679585382
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679585382
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679585382
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679585382
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679585382
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679585382
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679585382
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679585382
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679585382
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679585382
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679585382
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679585382
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679585382
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679585382
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679585382
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679585382
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679585382
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679585382
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679585382
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679585382
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679585382
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679585382
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679585382
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679585382
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679585382
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_924
timestamp 1679585382
transform 1 0 89280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_931
timestamp 1679585382
transform 1 0 89952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_938
timestamp 1679585382
transform 1 0 90624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_945
timestamp 1679585382
transform 1 0 91296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_952
timestamp 1679585382
transform 1 0 91968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_959
timestamp 1679585382
transform 1 0 92640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_966
timestamp 1679585382
transform 1 0 93312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_973
timestamp 1679585382
transform 1 0 93984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_980
timestamp 1679585382
transform 1 0 94656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_987
timestamp 1679585382
transform 1 0 95328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_994
timestamp 1679585382
transform 1 0 96000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1001
timestamp 1679585382
transform 1 0 96672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1008
timestamp 1679585382
transform 1 0 97344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1015
timestamp 1679585382
transform 1 0 98016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1022
timestamp 1679585382
transform 1 0 98688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679585382
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679585382
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679585382
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679585382
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679585382
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679585382
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679585382
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679585382
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679585382
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679585382
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679585382
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679585382
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679585382
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679585382
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679585382
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679585382
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679585382
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679585382
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679585382
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679585382
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679585382
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679585382
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679585382
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679585382
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679585382
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679585382
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679585382
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679585382
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679585382
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679585382
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679585382
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679585382
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679585382
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679585382
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679585382
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679585382
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679585382
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679585382
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679585382
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679585382
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679585382
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679585382
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679585382
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679585382
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679585382
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679585382
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679585382
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679585382
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679585382
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679585382
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679585382
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679585382
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679585382
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679585382
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679585382
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679585382
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679585382
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679585382
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679585382
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679585382
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679585382
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679585382
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679585382
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679585382
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679585382
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679585382
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679585382
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679585382
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679585382
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679585382
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679585382
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679585382
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679585382
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679585382
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679585382
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679585382
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679585382
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679585382
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679585382
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679585382
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679585382
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679585382
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679585382
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679585382
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679585382
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679585382
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679585382
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679585382
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679585382
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679585382
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679585382
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679585382
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679585382
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679585382
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679585382
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679585382
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679585382
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679585382
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679585382
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679585382
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679585382
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679585382
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679585382
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679585382
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679585382
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679585382
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679585382
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679585382
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679585382
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679585382
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679585382
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679585382
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679585382
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679585382
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679585382
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679585382
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679585382
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679585382
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679585382
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679585382
transform 1 0 80544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_840
timestamp 1679585382
transform 1 0 81216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_847
timestamp 1679585382
transform 1 0 81888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_854
timestamp 1679585382
transform 1 0 82560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_861
timestamp 1679585382
transform 1 0 83232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_868
timestamp 1679585382
transform 1 0 83904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_875
timestamp 1679585382
transform 1 0 84576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_882
timestamp 1679585382
transform 1 0 85248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_889
timestamp 1679585382
transform 1 0 85920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_896
timestamp 1679585382
transform 1 0 86592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_903
timestamp 1679585382
transform 1 0 87264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_910
timestamp 1679585382
transform 1 0 87936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_917
timestamp 1679585382
transform 1 0 88608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_924
timestamp 1679585382
transform 1 0 89280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_931
timestamp 1679585382
transform 1 0 89952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_938
timestamp 1679585382
transform 1 0 90624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_945
timestamp 1679585382
transform 1 0 91296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_952
timestamp 1679585382
transform 1 0 91968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_959
timestamp 1679585382
transform 1 0 92640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_966
timestamp 1679585382
transform 1 0 93312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_973
timestamp 1679585382
transform 1 0 93984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_980
timestamp 1679585382
transform 1 0 94656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_987
timestamp 1679585382
transform 1 0 95328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_994
timestamp 1679585382
transform 1 0 96000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1001
timestamp 1679585382
transform 1 0 96672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1008
timestamp 1679585382
transform 1 0 97344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1015
timestamp 1679585382
transform 1 0 98016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1022
timestamp 1679585382
transform 1 0 98688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679585382
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679585382
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_18
timestamp 1677583704
transform 1 0 2304 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_20
timestamp 1677583258
transform 1 0 2496 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_25
timestamp 1679581501
transform 1 0 2976 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_29
timestamp 1677583704
transform 1 0 3360 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_58
timestamp 1679585382
transform 1 0 6144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_65
timestamp 1679585382
transform 1 0 6816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_72
timestamp 1679585382
transform 1 0 7488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_79
timestamp 1679585382
transform 1 0 8160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_86
timestamp 1679585382
transform 1 0 8832 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_93
timestamp 1677583258
transform 1 0 9504 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679585382
transform 1 0 9984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679585382
transform 1 0 10656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679585382
transform 1 0 11328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679585382
transform 1 0 12000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679585382
transform 1 0 12672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679585382
transform 1 0 13344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679585382
transform 1 0 14016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679585382
transform 1 0 14688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679585382
transform 1 0 15360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679585382
transform 1 0 16032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679585382
transform 1 0 16704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679585382
transform 1 0 17376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679585382
transform 1 0 18048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679585382
transform 1 0 18720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1679585382
transform 1 0 19392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1679585382
transform 1 0 20064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1679585382
transform 1 0 20736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1679585382
transform 1 0 21408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679585382
transform 1 0 22080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1679585382
transform 1 0 22752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1679585382
transform 1 0 23424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1679585382
transform 1 0 24096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_252
timestamp 1679585382
transform 1 0 24768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_259
timestamp 1679585382
transform 1 0 25440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_266
timestamp 1679585382
transform 1 0 26112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_273
timestamp 1679585382
transform 1 0 26784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_280
timestamp 1679585382
transform 1 0 27456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_287
timestamp 1679585382
transform 1 0 28128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_294
timestamp 1679585382
transform 1 0 28800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_301
timestamp 1679585382
transform 1 0 29472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_308
timestamp 1679585382
transform 1 0 30144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_315
timestamp 1679585382
transform 1 0 30816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_322
timestamp 1679585382
transform 1 0 31488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_329
timestamp 1679585382
transform 1 0 32160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_336
timestamp 1679585382
transform 1 0 32832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_343
timestamp 1679585382
transform 1 0 33504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_350
timestamp 1679585382
transform 1 0 34176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_357
timestamp 1679585382
transform 1 0 34848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_364
timestamp 1679585382
transform 1 0 35520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_371
timestamp 1679585382
transform 1 0 36192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_378
timestamp 1679585382
transform 1 0 36864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_385
timestamp 1679585382
transform 1 0 37536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_392
timestamp 1679585382
transform 1 0 38208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_399
timestamp 1679585382
transform 1 0 38880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_406
timestamp 1679585382
transform 1 0 39552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_413
timestamp 1679585382
transform 1 0 40224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_420
timestamp 1679585382
transform 1 0 40896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_427
timestamp 1679585382
transform 1 0 41568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_434
timestamp 1679585382
transform 1 0 42240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_441
timestamp 1679585382
transform 1 0 42912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_448
timestamp 1679585382
transform 1 0 43584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_455
timestamp 1679585382
transform 1 0 44256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_462
timestamp 1679585382
transform 1 0 44928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_469
timestamp 1679585382
transform 1 0 45600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_476
timestamp 1679585382
transform 1 0 46272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_483
timestamp 1679585382
transform 1 0 46944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_490
timestamp 1679585382
transform 1 0 47616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_497
timestamp 1679585382
transform 1 0 48288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_504
timestamp 1679585382
transform 1 0 48960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_511
timestamp 1679585382
transform 1 0 49632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_518
timestamp 1679585382
transform 1 0 50304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_525
timestamp 1679585382
transform 1 0 50976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_532
timestamp 1679585382
transform 1 0 51648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_539
timestamp 1679585382
transform 1 0 52320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_546
timestamp 1679585382
transform 1 0 52992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_553
timestamp 1679585382
transform 1 0 53664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_560
timestamp 1679585382
transform 1 0 54336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_567
timestamp 1679585382
transform 1 0 55008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_574
timestamp 1679585382
transform 1 0 55680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_581
timestamp 1679585382
transform 1 0 56352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_588
timestamp 1679585382
transform 1 0 57024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_595
timestamp 1679585382
transform 1 0 57696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_602
timestamp 1679585382
transform 1 0 58368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_609
timestamp 1679585382
transform 1 0 59040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_616
timestamp 1679585382
transform 1 0 59712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_623
timestamp 1679585382
transform 1 0 60384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_630
timestamp 1679585382
transform 1 0 61056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_637
timestamp 1679585382
transform 1 0 61728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_644
timestamp 1679585382
transform 1 0 62400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_651
timestamp 1679585382
transform 1 0 63072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_658
timestamp 1679585382
transform 1 0 63744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_665
timestamp 1679585382
transform 1 0 64416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_672
timestamp 1679585382
transform 1 0 65088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_679
timestamp 1679585382
transform 1 0 65760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_686
timestamp 1679585382
transform 1 0 66432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_693
timestamp 1679585382
transform 1 0 67104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_700
timestamp 1679585382
transform 1 0 67776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_707
timestamp 1679585382
transform 1 0 68448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_714
timestamp 1679585382
transform 1 0 69120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_721
timestamp 1679585382
transform 1 0 69792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_728
timestamp 1679585382
transform 1 0 70464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_735
timestamp 1679585382
transform 1 0 71136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_742
timestamp 1679585382
transform 1 0 71808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_749
timestamp 1679585382
transform 1 0 72480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_756
timestamp 1679585382
transform 1 0 73152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_763
timestamp 1679585382
transform 1 0 73824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_770
timestamp 1679585382
transform 1 0 74496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_777
timestamp 1679585382
transform 1 0 75168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_784
timestamp 1679585382
transform 1 0 75840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_791
timestamp 1679585382
transform 1 0 76512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_798
timestamp 1679585382
transform 1 0 77184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_805
timestamp 1679585382
transform 1 0 77856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_812
timestamp 1679585382
transform 1 0 78528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_819
timestamp 1679585382
transform 1 0 79200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_826
timestamp 1679585382
transform 1 0 79872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_833
timestamp 1679585382
transform 1 0 80544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_840
timestamp 1679585382
transform 1 0 81216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_847
timestamp 1679585382
transform 1 0 81888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_854
timestamp 1679585382
transform 1 0 82560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_861
timestamp 1679585382
transform 1 0 83232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_868
timestamp 1679585382
transform 1 0 83904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_875
timestamp 1679585382
transform 1 0 84576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_882
timestamp 1679585382
transform 1 0 85248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_889
timestamp 1679585382
transform 1 0 85920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_896
timestamp 1679585382
transform 1 0 86592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_903
timestamp 1679585382
transform 1 0 87264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_910
timestamp 1679585382
transform 1 0 87936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_917
timestamp 1679585382
transform 1 0 88608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_924
timestamp 1679585382
transform 1 0 89280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_931
timestamp 1679585382
transform 1 0 89952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_938
timestamp 1679585382
transform 1 0 90624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_945
timestamp 1679585382
transform 1 0 91296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_952
timestamp 1679585382
transform 1 0 91968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_959
timestamp 1679585382
transform 1 0 92640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_966
timestamp 1679585382
transform 1 0 93312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_973
timestamp 1679585382
transform 1 0 93984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_980
timestamp 1679585382
transform 1 0 94656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_987
timestamp 1679585382
transform 1 0 95328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_994
timestamp 1679585382
transform 1 0 96000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1001
timestamp 1679585382
transform 1 0 96672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1008
timestamp 1679585382
transform 1 0 97344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1015
timestamp 1679585382
transform 1 0 98016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1022
timestamp 1679585382
transform 1 0 98688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679585382
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679585382
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679585382
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679585382
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_32
timestamp 1679581501
transform 1 0 3648 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_40
timestamp 1679585382
transform 1 0 4416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_47
timestamp 1679585382
transform 1 0 5088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_54
timestamp 1679585382
transform 1 0 5760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_61
timestamp 1679585382
transform 1 0 6432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_68
timestamp 1679585382
transform 1 0 7104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_75
timestamp 1679585382
transform 1 0 7776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_82
timestamp 1679585382
transform 1 0 8448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679585382
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679585382
transform 1 0 12384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679585382
transform 1 0 13056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679585382
transform 1 0 13728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679585382
transform 1 0 14400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679585382
transform 1 0 15072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679585382
transform 1 0 15744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679585382
transform 1 0 16416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679585382
transform 1 0 17088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679585382
transform 1 0 17760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679585382
transform 1 0 18432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679585382
transform 1 0 19104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_200
timestamp 1679585382
transform 1 0 19776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_207
timestamp 1679585382
transform 1 0 20448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_214
timestamp 1679585382
transform 1 0 21120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_221
timestamp 1679585382
transform 1 0 21792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_228
timestamp 1679585382
transform 1 0 22464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_235
timestamp 1679585382
transform 1 0 23136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_242
timestamp 1679585382
transform 1 0 23808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_249
timestamp 1679585382
transform 1 0 24480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_256
timestamp 1679585382
transform 1 0 25152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_263
timestamp 1679585382
transform 1 0 25824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_270
timestamp 1679585382
transform 1 0 26496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_277
timestamp 1679585382
transform 1 0 27168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_284
timestamp 1679585382
transform 1 0 27840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_291
timestamp 1679585382
transform 1 0 28512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679585382
transform 1 0 29184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679585382
transform 1 0 29856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_312
timestamp 1679585382
transform 1 0 30528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_319
timestamp 1679585382
transform 1 0 31200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_326
timestamp 1679585382
transform 1 0 31872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_333
timestamp 1679585382
transform 1 0 32544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_340
timestamp 1679585382
transform 1 0 33216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_347
timestamp 1679585382
transform 1 0 33888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_354
timestamp 1679585382
transform 1 0 34560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_361
timestamp 1679585382
transform 1 0 35232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_368
timestamp 1679585382
transform 1 0 35904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_375
timestamp 1679585382
transform 1 0 36576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_382
timestamp 1679585382
transform 1 0 37248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_389
timestamp 1679585382
transform 1 0 37920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_396
timestamp 1679585382
transform 1 0 38592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_403
timestamp 1679585382
transform 1 0 39264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_410
timestamp 1679585382
transform 1 0 39936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_417
timestamp 1679585382
transform 1 0 40608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_424
timestamp 1679585382
transform 1 0 41280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_431
timestamp 1679585382
transform 1 0 41952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_438
timestamp 1679585382
transform 1 0 42624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_445
timestamp 1679585382
transform 1 0 43296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_452
timestamp 1679585382
transform 1 0 43968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_459
timestamp 1679585382
transform 1 0 44640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_466
timestamp 1679585382
transform 1 0 45312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_473
timestamp 1679585382
transform 1 0 45984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_480
timestamp 1679585382
transform 1 0 46656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_487
timestamp 1679585382
transform 1 0 47328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_494
timestamp 1679585382
transform 1 0 48000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_501
timestamp 1679585382
transform 1 0 48672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_508
timestamp 1679585382
transform 1 0 49344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_515
timestamp 1679585382
transform 1 0 50016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_522
timestamp 1679585382
transform 1 0 50688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_529
timestamp 1679585382
transform 1 0 51360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_536
timestamp 1679585382
transform 1 0 52032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_543
timestamp 1679585382
transform 1 0 52704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_550
timestamp 1679585382
transform 1 0 53376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_557
timestamp 1679585382
transform 1 0 54048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_564
timestamp 1679585382
transform 1 0 54720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_571
timestamp 1679585382
transform 1 0 55392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_578
timestamp 1679585382
transform 1 0 56064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_585
timestamp 1679585382
transform 1 0 56736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_592
timestamp 1679585382
transform 1 0 57408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_599
timestamp 1679585382
transform 1 0 58080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_606
timestamp 1679585382
transform 1 0 58752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_613
timestamp 1679585382
transform 1 0 59424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_620
timestamp 1679585382
transform 1 0 60096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_627
timestamp 1679585382
transform 1 0 60768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_634
timestamp 1679585382
transform 1 0 61440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_641
timestamp 1679585382
transform 1 0 62112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_648
timestamp 1679585382
transform 1 0 62784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_655
timestamp 1679585382
transform 1 0 63456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_662
timestamp 1679585382
transform 1 0 64128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_669
timestamp 1679585382
transform 1 0 64800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_676
timestamp 1679585382
transform 1 0 65472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_683
timestamp 1679585382
transform 1 0 66144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_690
timestamp 1679585382
transform 1 0 66816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_697
timestamp 1679585382
transform 1 0 67488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_704
timestamp 1679585382
transform 1 0 68160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_711
timestamp 1679585382
transform 1 0 68832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_718
timestamp 1679585382
transform 1 0 69504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_725
timestamp 1679585382
transform 1 0 70176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_732
timestamp 1679585382
transform 1 0 70848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_739
timestamp 1679585382
transform 1 0 71520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_746
timestamp 1679585382
transform 1 0 72192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_753
timestamp 1679585382
transform 1 0 72864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_760
timestamp 1679585382
transform 1 0 73536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_767
timestamp 1679585382
transform 1 0 74208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_774
timestamp 1679585382
transform 1 0 74880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_781
timestamp 1679585382
transform 1 0 75552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_788
timestamp 1679585382
transform 1 0 76224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_795
timestamp 1679585382
transform 1 0 76896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_802
timestamp 1679585382
transform 1 0 77568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679585382
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679585382
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_823
timestamp 1679585382
transform 1 0 79584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_830
timestamp 1679585382
transform 1 0 80256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_837
timestamp 1679585382
transform 1 0 80928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_844
timestamp 1679585382
transform 1 0 81600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_851
timestamp 1679585382
transform 1 0 82272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_858
timestamp 1679585382
transform 1 0 82944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_865
timestamp 1679585382
transform 1 0 83616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_872
timestamp 1679585382
transform 1 0 84288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_879
timestamp 1679585382
transform 1 0 84960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_886
timestamp 1679585382
transform 1 0 85632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_893
timestamp 1679585382
transform 1 0 86304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_900
timestamp 1679585382
transform 1 0 86976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_907
timestamp 1679585382
transform 1 0 87648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_914
timestamp 1679585382
transform 1 0 88320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_921
timestamp 1679585382
transform 1 0 88992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_928
timestamp 1679585382
transform 1 0 89664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_935
timestamp 1679585382
transform 1 0 90336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_942
timestamp 1679585382
transform 1 0 91008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_949
timestamp 1679585382
transform 1 0 91680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_956
timestamp 1679585382
transform 1 0 92352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_963
timestamp 1679585382
transform 1 0 93024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_970
timestamp 1679585382
transform 1 0 93696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_977
timestamp 1679585382
transform 1 0 94368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_984
timestamp 1679585382
transform 1 0 95040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_991
timestamp 1679585382
transform 1 0 95712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_998
timestamp 1679585382
transform 1 0 96384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1005
timestamp 1679585382
transform 1 0 97056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1012
timestamp 1679585382
transform 1 0 97728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1019
timestamp 1679585382
transform 1 0 98400 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_1026
timestamp 1677583704
transform 1 0 99072 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_1028
timestamp 1677583258
transform 1 0 99264 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679585382
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679585382
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_18
timestamp 1677583704
transform 1 0 2304 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_20
timestamp 1677583258
transform 1 0 2496 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679585382
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_32
timestamp 1679581501
transform 1 0 3648 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_45
timestamp 1677583704
transform 1 0 4896 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679585382
transform 1 0 5952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679585382
transform 1 0 6624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679585382
transform 1 0 7296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679585382
transform 1 0 7968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_84
timestamp 1679581501
transform 1 0 8640 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_88
timestamp 1677583704
transform 1 0 9024 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679585382
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_102
timestamp 1677583704
transform 1 0 10368 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_113
timestamp 1679585382
transform 1 0 11424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_120
timestamp 1679585382
transform 1 0 12096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_127
timestamp 1679585382
transform 1 0 12768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_134
timestamp 1679585382
transform 1 0 13440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_141
timestamp 1679585382
transform 1 0 14112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_148
timestamp 1679585382
transform 1 0 14784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_155
timestamp 1679585382
transform 1 0 15456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_162
timestamp 1679585382
transform 1 0 16128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_169
timestamp 1679585382
transform 1 0 16800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_176
timestamp 1679585382
transform 1 0 17472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_183
timestamp 1679585382
transform 1 0 18144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_190
timestamp 1679585382
transform 1 0 18816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_197
timestamp 1679585382
transform 1 0 19488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_204
timestamp 1679585382
transform 1 0 20160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_211
timestamp 1679585382
transform 1 0 20832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_218
timestamp 1679585382
transform 1 0 21504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_225
timestamp 1679585382
transform 1 0 22176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_232
timestamp 1679585382
transform 1 0 22848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_239
timestamp 1679585382
transform 1 0 23520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_246
timestamp 1679585382
transform 1 0 24192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_253
timestamp 1679585382
transform 1 0 24864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_260
timestamp 1679585382
transform 1 0 25536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_267
timestamp 1679585382
transform 1 0 26208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_274
timestamp 1679585382
transform 1 0 26880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_281
timestamp 1679585382
transform 1 0 27552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_288
timestamp 1679585382
transform 1 0 28224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_295
timestamp 1679585382
transform 1 0 28896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_302
timestamp 1679585382
transform 1 0 29568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_309
timestamp 1679585382
transform 1 0 30240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_316
timestamp 1679585382
transform 1 0 30912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_323
timestamp 1679585382
transform 1 0 31584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_330
timestamp 1679585382
transform 1 0 32256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_337
timestamp 1679585382
transform 1 0 32928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_344
timestamp 1679585382
transform 1 0 33600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_351
timestamp 1679585382
transform 1 0 34272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_358
timestamp 1679585382
transform 1 0 34944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_365
timestamp 1679585382
transform 1 0 35616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_372
timestamp 1679585382
transform 1 0 36288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_379
timestamp 1679585382
transform 1 0 36960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_386
timestamp 1679585382
transform 1 0 37632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_393
timestamp 1679585382
transform 1 0 38304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_400
timestamp 1679585382
transform 1 0 38976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_407
timestamp 1679585382
transform 1 0 39648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_414
timestamp 1679585382
transform 1 0 40320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_421
timestamp 1679585382
transform 1 0 40992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_428
timestamp 1679585382
transform 1 0 41664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_435
timestamp 1679585382
transform 1 0 42336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_442
timestamp 1679585382
transform 1 0 43008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_449
timestamp 1679585382
transform 1 0 43680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_456
timestamp 1679585382
transform 1 0 44352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_463
timestamp 1679585382
transform 1 0 45024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_470
timestamp 1679585382
transform 1 0 45696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_477
timestamp 1679585382
transform 1 0 46368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_484
timestamp 1679585382
transform 1 0 47040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_491
timestamp 1679585382
transform 1 0 47712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_498
timestamp 1679585382
transform 1 0 48384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_505
timestamp 1679585382
transform 1 0 49056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_512
timestamp 1679585382
transform 1 0 49728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_519
timestamp 1679585382
transform 1 0 50400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_526
timestamp 1679585382
transform 1 0 51072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_533
timestamp 1679585382
transform 1 0 51744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_540
timestamp 1679585382
transform 1 0 52416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_547
timestamp 1679585382
transform 1 0 53088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_554
timestamp 1679585382
transform 1 0 53760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_561
timestamp 1679585382
transform 1 0 54432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_568
timestamp 1679585382
transform 1 0 55104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_575
timestamp 1679585382
transform 1 0 55776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_582
timestamp 1679585382
transform 1 0 56448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_589
timestamp 1679585382
transform 1 0 57120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_596
timestamp 1679585382
transform 1 0 57792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_603
timestamp 1679585382
transform 1 0 58464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_610
timestamp 1679585382
transform 1 0 59136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_617
timestamp 1679585382
transform 1 0 59808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_624
timestamp 1679585382
transform 1 0 60480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_631
timestamp 1679585382
transform 1 0 61152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_638
timestamp 1679585382
transform 1 0 61824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_645
timestamp 1679585382
transform 1 0 62496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_652
timestamp 1679585382
transform 1 0 63168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_659
timestamp 1679585382
transform 1 0 63840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_666
timestamp 1679585382
transform 1 0 64512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_673
timestamp 1679585382
transform 1 0 65184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_680
timestamp 1679585382
transform 1 0 65856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_687
timestamp 1679585382
transform 1 0 66528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_694
timestamp 1679585382
transform 1 0 67200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_701
timestamp 1679585382
transform 1 0 67872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_708
timestamp 1679585382
transform 1 0 68544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_715
timestamp 1679585382
transform 1 0 69216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_722
timestamp 1679585382
transform 1 0 69888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_729
timestamp 1679585382
transform 1 0 70560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_736
timestamp 1679585382
transform 1 0 71232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_743
timestamp 1679585382
transform 1 0 71904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_750
timestamp 1679585382
transform 1 0 72576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_757
timestamp 1679585382
transform 1 0 73248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_764
timestamp 1679585382
transform 1 0 73920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_771
timestamp 1679585382
transform 1 0 74592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_778
timestamp 1679585382
transform 1 0 75264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_785
timestamp 1679585382
transform 1 0 75936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_792
timestamp 1679585382
transform 1 0 76608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_799
timestamp 1679585382
transform 1 0 77280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_806
timestamp 1679585382
transform 1 0 77952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_813
timestamp 1679585382
transform 1 0 78624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_820
timestamp 1679585382
transform 1 0 79296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_827
timestamp 1679585382
transform 1 0 79968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_834
timestamp 1679585382
transform 1 0 80640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_841
timestamp 1679585382
transform 1 0 81312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_848
timestamp 1679585382
transform 1 0 81984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_855
timestamp 1679585382
transform 1 0 82656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_862
timestamp 1679585382
transform 1 0 83328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_869
timestamp 1679585382
transform 1 0 84000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_876
timestamp 1679585382
transform 1 0 84672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_883
timestamp 1679585382
transform 1 0 85344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_890
timestamp 1679585382
transform 1 0 86016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_897
timestamp 1679585382
transform 1 0 86688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_904
timestamp 1679585382
transform 1 0 87360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_911
timestamp 1679585382
transform 1 0 88032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_918
timestamp 1679585382
transform 1 0 88704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_925
timestamp 1679585382
transform 1 0 89376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_932
timestamp 1679585382
transform 1 0 90048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_939
timestamp 1679585382
transform 1 0 90720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_946
timestamp 1679585382
transform 1 0 91392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_953
timestamp 1679585382
transform 1 0 92064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_960
timestamp 1679585382
transform 1 0 92736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_967
timestamp 1679585382
transform 1 0 93408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_974
timestamp 1679585382
transform 1 0 94080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_981
timestamp 1679585382
transform 1 0 94752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_988
timestamp 1679585382
transform 1 0 95424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_995
timestamp 1679585382
transform 1 0 96096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1002
timestamp 1679585382
transform 1 0 96768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1009
timestamp 1679585382
transform 1 0 97440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1016
timestamp 1679585382
transform 1 0 98112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_1023
timestamp 1679581501
transform 1 0 98784 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_1027
timestamp 1677583704
transform 1 0 99168 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679585382
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679585382
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_18
timestamp 1677583704
transform 1 0 2304 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_20
timestamp 1677583258
transform 1 0 2496 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679585382
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_32
timestamp 1677583258
transform 1 0 3648 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679585382
transform 1 0 4608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679585382
transform 1 0 5280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679585382
transform 1 0 5952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679585382
transform 1 0 6624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679585382
transform 1 0 7296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679585382
transform 1 0 7968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_84
timestamp 1679581501
transform 1 0 8640 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_88
timestamp 1677583258
transform 1 0 9024 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_94
timestamp 1679585382
transform 1 0 9600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_101
timestamp 1679585382
transform 1 0 10272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_108
timestamp 1679585382
transform 1 0 10944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_115
timestamp 1679585382
transform 1 0 11616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_122
timestamp 1679585382
transform 1 0 12288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_129
timestamp 1679585382
transform 1 0 12960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_136
timestamp 1679585382
transform 1 0 13632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_143
timestamp 1679585382
transform 1 0 14304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_150
timestamp 1679585382
transform 1 0 14976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_157
timestamp 1679585382
transform 1 0 15648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_164
timestamp 1679585382
transform 1 0 16320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_171
timestamp 1679585382
transform 1 0 16992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_178
timestamp 1679585382
transform 1 0 17664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_185
timestamp 1679585382
transform 1 0 18336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_192
timestamp 1679585382
transform 1 0 19008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_199
timestamp 1679585382
transform 1 0 19680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_206
timestamp 1679585382
transform 1 0 20352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_213
timestamp 1679585382
transform 1 0 21024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_220
timestamp 1679585382
transform 1 0 21696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_227
timestamp 1679585382
transform 1 0 22368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_234
timestamp 1679585382
transform 1 0 23040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_241
timestamp 1679585382
transform 1 0 23712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_248
timestamp 1679585382
transform 1 0 24384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_255
timestamp 1679585382
transform 1 0 25056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_262
timestamp 1679585382
transform 1 0 25728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_269
timestamp 1679585382
transform 1 0 26400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_276
timestamp 1679585382
transform 1 0 27072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_283
timestamp 1679585382
transform 1 0 27744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_290
timestamp 1679585382
transform 1 0 28416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_297
timestamp 1679585382
transform 1 0 29088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_304
timestamp 1679585382
transform 1 0 29760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_311
timestamp 1679585382
transform 1 0 30432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_318
timestamp 1679585382
transform 1 0 31104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_325
timestamp 1679585382
transform 1 0 31776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_332
timestamp 1679585382
transform 1 0 32448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_339
timestamp 1679585382
transform 1 0 33120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_346
timestamp 1679585382
transform 1 0 33792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_353
timestamp 1679585382
transform 1 0 34464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_360
timestamp 1679585382
transform 1 0 35136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_367
timestamp 1679585382
transform 1 0 35808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_374
timestamp 1679585382
transform 1 0 36480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_381
timestamp 1679585382
transform 1 0 37152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_388
timestamp 1679585382
transform 1 0 37824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_395
timestamp 1679585382
transform 1 0 38496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_402
timestamp 1679585382
transform 1 0 39168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_409
timestamp 1679585382
transform 1 0 39840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_416
timestamp 1679585382
transform 1 0 40512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_423
timestamp 1679585382
transform 1 0 41184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_430
timestamp 1679585382
transform 1 0 41856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_437
timestamp 1679585382
transform 1 0 42528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_444
timestamp 1679585382
transform 1 0 43200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_451
timestamp 1679585382
transform 1 0 43872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_458
timestamp 1679585382
transform 1 0 44544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_465
timestamp 1679585382
transform 1 0 45216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_472
timestamp 1679585382
transform 1 0 45888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_479
timestamp 1679585382
transform 1 0 46560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_486
timestamp 1679585382
transform 1 0 47232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_493
timestamp 1679585382
transform 1 0 47904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_500
timestamp 1679585382
transform 1 0 48576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_507
timestamp 1679585382
transform 1 0 49248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_514
timestamp 1679585382
transform 1 0 49920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_521
timestamp 1679585382
transform 1 0 50592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_528
timestamp 1679585382
transform 1 0 51264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_535
timestamp 1679585382
transform 1 0 51936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_542
timestamp 1679585382
transform 1 0 52608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_549
timestamp 1679585382
transform 1 0 53280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_556
timestamp 1679585382
transform 1 0 53952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_563
timestamp 1679585382
transform 1 0 54624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_570
timestamp 1679585382
transform 1 0 55296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_577
timestamp 1679585382
transform 1 0 55968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_584
timestamp 1679585382
transform 1 0 56640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_591
timestamp 1679585382
transform 1 0 57312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_598
timestamp 1679585382
transform 1 0 57984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_605
timestamp 1679585382
transform 1 0 58656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_612
timestamp 1679585382
transform 1 0 59328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_619
timestamp 1679585382
transform 1 0 60000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_626
timestamp 1679585382
transform 1 0 60672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_633
timestamp 1679585382
transform 1 0 61344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_640
timestamp 1679585382
transform 1 0 62016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_647
timestamp 1679585382
transform 1 0 62688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_654
timestamp 1679585382
transform 1 0 63360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_661
timestamp 1679585382
transform 1 0 64032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_668
timestamp 1679585382
transform 1 0 64704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_675
timestamp 1679585382
transform 1 0 65376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_682
timestamp 1679585382
transform 1 0 66048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_689
timestamp 1679585382
transform 1 0 66720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_696
timestamp 1679585382
transform 1 0 67392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_703
timestamp 1679585382
transform 1 0 68064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_710
timestamp 1679585382
transform 1 0 68736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_717
timestamp 1679585382
transform 1 0 69408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_724
timestamp 1679585382
transform 1 0 70080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_731
timestamp 1679585382
transform 1 0 70752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_738
timestamp 1679585382
transform 1 0 71424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_745
timestamp 1679585382
transform 1 0 72096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_752
timestamp 1679585382
transform 1 0 72768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_759
timestamp 1679585382
transform 1 0 73440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_766
timestamp 1679585382
transform 1 0 74112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_773
timestamp 1679585382
transform 1 0 74784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_780
timestamp 1679585382
transform 1 0 75456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_787
timestamp 1679585382
transform 1 0 76128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_794
timestamp 1679585382
transform 1 0 76800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_801
timestamp 1679585382
transform 1 0 77472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_808
timestamp 1679585382
transform 1 0 78144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_815
timestamp 1679585382
transform 1 0 78816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_822
timestamp 1679585382
transform 1 0 79488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_829
timestamp 1679585382
transform 1 0 80160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_836
timestamp 1679585382
transform 1 0 80832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_843
timestamp 1679585382
transform 1 0 81504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_850
timestamp 1679585382
transform 1 0 82176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_857
timestamp 1679585382
transform 1 0 82848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_864
timestamp 1679585382
transform 1 0 83520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_871
timestamp 1679585382
transform 1 0 84192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_878
timestamp 1679585382
transform 1 0 84864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_885
timestamp 1679585382
transform 1 0 85536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_892
timestamp 1679585382
transform 1 0 86208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_899
timestamp 1679585382
transform 1 0 86880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_906
timestamp 1679585382
transform 1 0 87552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_913
timestamp 1679585382
transform 1 0 88224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_920
timestamp 1679585382
transform 1 0 88896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_927
timestamp 1679585382
transform 1 0 89568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_934
timestamp 1679585382
transform 1 0 90240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_941
timestamp 1679585382
transform 1 0 90912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_948
timestamp 1679585382
transform 1 0 91584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_955
timestamp 1679585382
transform 1 0 92256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_962
timestamp 1679585382
transform 1 0 92928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_969
timestamp 1679585382
transform 1 0 93600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_976
timestamp 1679585382
transform 1 0 94272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_983
timestamp 1679585382
transform 1 0 94944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_990
timestamp 1679585382
transform 1 0 95616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_997
timestamp 1679585382
transform 1 0 96288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1004
timestamp 1679585382
transform 1 0 96960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1011
timestamp 1679585382
transform 1 0 97632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1018
timestamp 1679585382
transform 1 0 98304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_1025
timestamp 1679581501
transform 1 0 98976 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679585382
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679585382
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679585382
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679585382
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_32
timestamp 1679581501
transform 1 0 3648 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_36
timestamp 1677583704
transform 1 0 4032 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_47
timestamp 1679585382
transform 1 0 5088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_54
timestamp 1679585382
transform 1 0 5760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_61
timestamp 1679585382
transform 1 0 6432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_68
timestamp 1679585382
transform 1 0 7104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_75
timestamp 1679585382
transform 1 0 7776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_82
timestamp 1679585382
transform 1 0 8448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_89
timestamp 1679585382
transform 1 0 9120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_96
timestamp 1679585382
transform 1 0 9792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_103
timestamp 1679585382
transform 1 0 10464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_110
timestamp 1679585382
transform 1 0 11136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_117
timestamp 1679585382
transform 1 0 11808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_124
timestamp 1679585382
transform 1 0 12480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_131
timestamp 1679585382
transform 1 0 13152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_138
timestamp 1679585382
transform 1 0 13824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_145
timestamp 1679585382
transform 1 0 14496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_152
timestamp 1679585382
transform 1 0 15168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_159
timestamp 1679585382
transform 1 0 15840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_166
timestamp 1679585382
transform 1 0 16512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_173
timestamp 1679585382
transform 1 0 17184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_180
timestamp 1679585382
transform 1 0 17856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_187
timestamp 1679585382
transform 1 0 18528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_194
timestamp 1679585382
transform 1 0 19200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_201
timestamp 1679585382
transform 1 0 19872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_208
timestamp 1679585382
transform 1 0 20544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_215
timestamp 1679585382
transform 1 0 21216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_222
timestamp 1679585382
transform 1 0 21888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_229
timestamp 1679585382
transform 1 0 22560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_236
timestamp 1679585382
transform 1 0 23232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_243
timestamp 1679585382
transform 1 0 23904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_250
timestamp 1679585382
transform 1 0 24576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_257
timestamp 1679585382
transform 1 0 25248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_264
timestamp 1679585382
transform 1 0 25920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_271
timestamp 1679585382
transform 1 0 26592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_278
timestamp 1679585382
transform 1 0 27264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_285
timestamp 1679585382
transform 1 0 27936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_292
timestamp 1679585382
transform 1 0 28608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_299
timestamp 1679585382
transform 1 0 29280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_306
timestamp 1679585382
transform 1 0 29952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_313
timestamp 1679585382
transform 1 0 30624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_320
timestamp 1679585382
transform 1 0 31296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_327
timestamp 1679585382
transform 1 0 31968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_334
timestamp 1679585382
transform 1 0 32640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_341
timestamp 1679585382
transform 1 0 33312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_348
timestamp 1679585382
transform 1 0 33984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_355
timestamp 1679585382
transform 1 0 34656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_362
timestamp 1679585382
transform 1 0 35328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_369
timestamp 1679585382
transform 1 0 36000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_376
timestamp 1679585382
transform 1 0 36672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_383
timestamp 1679585382
transform 1 0 37344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_390
timestamp 1679585382
transform 1 0 38016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_397
timestamp 1679585382
transform 1 0 38688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_404
timestamp 1679585382
transform 1 0 39360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_411
timestamp 1679585382
transform 1 0 40032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_418
timestamp 1679585382
transform 1 0 40704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_425
timestamp 1679585382
transform 1 0 41376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_432
timestamp 1679585382
transform 1 0 42048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_439
timestamp 1679585382
transform 1 0 42720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_446
timestamp 1679585382
transform 1 0 43392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_453
timestamp 1679585382
transform 1 0 44064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_460
timestamp 1679585382
transform 1 0 44736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_467
timestamp 1679585382
transform 1 0 45408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_474
timestamp 1679585382
transform 1 0 46080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_481
timestamp 1679585382
transform 1 0 46752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_488
timestamp 1679585382
transform 1 0 47424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_495
timestamp 1679585382
transform 1 0 48096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_502
timestamp 1679585382
transform 1 0 48768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_509
timestamp 1679585382
transform 1 0 49440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_516
timestamp 1679585382
transform 1 0 50112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_523
timestamp 1679585382
transform 1 0 50784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_530
timestamp 1679585382
transform 1 0 51456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_537
timestamp 1679585382
transform 1 0 52128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_544
timestamp 1679585382
transform 1 0 52800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_551
timestamp 1679585382
transform 1 0 53472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_558
timestamp 1679585382
transform 1 0 54144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_565
timestamp 1679585382
transform 1 0 54816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_572
timestamp 1679585382
transform 1 0 55488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_579
timestamp 1679585382
transform 1 0 56160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_586
timestamp 1679585382
transform 1 0 56832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_593
timestamp 1679585382
transform 1 0 57504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_600
timestamp 1679585382
transform 1 0 58176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_607
timestamp 1679585382
transform 1 0 58848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_614
timestamp 1679585382
transform 1 0 59520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_621
timestamp 1679585382
transform 1 0 60192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_628
timestamp 1679585382
transform 1 0 60864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_635
timestamp 1679585382
transform 1 0 61536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_642
timestamp 1679585382
transform 1 0 62208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_649
timestamp 1679585382
transform 1 0 62880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_656
timestamp 1679585382
transform 1 0 63552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_663
timestamp 1679585382
transform 1 0 64224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_670
timestamp 1679585382
transform 1 0 64896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_677
timestamp 1679585382
transform 1 0 65568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_684
timestamp 1679585382
transform 1 0 66240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_691
timestamp 1679585382
transform 1 0 66912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_698
timestamp 1679585382
transform 1 0 67584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_705
timestamp 1679585382
transform 1 0 68256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_712
timestamp 1679585382
transform 1 0 68928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_719
timestamp 1679585382
transform 1 0 69600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_726
timestamp 1679585382
transform 1 0 70272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_733
timestamp 1679585382
transform 1 0 70944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_740
timestamp 1679585382
transform 1 0 71616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_747
timestamp 1679585382
transform 1 0 72288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_754
timestamp 1679585382
transform 1 0 72960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_761
timestamp 1679585382
transform 1 0 73632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_768
timestamp 1679585382
transform 1 0 74304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_775
timestamp 1679585382
transform 1 0 74976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_782
timestamp 1679585382
transform 1 0 75648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_789
timestamp 1679585382
transform 1 0 76320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_796
timestamp 1679585382
transform 1 0 76992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_803
timestamp 1679585382
transform 1 0 77664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_810
timestamp 1679585382
transform 1 0 78336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_817
timestamp 1679585382
transform 1 0 79008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_824
timestamp 1679585382
transform 1 0 79680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_831
timestamp 1679585382
transform 1 0 80352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_838
timestamp 1679585382
transform 1 0 81024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_845
timestamp 1679585382
transform 1 0 81696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_852
timestamp 1679585382
transform 1 0 82368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_859
timestamp 1679585382
transform 1 0 83040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_866
timestamp 1679585382
transform 1 0 83712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_873
timestamp 1679585382
transform 1 0 84384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_880
timestamp 1679585382
transform 1 0 85056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_887
timestamp 1679585382
transform 1 0 85728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_894
timestamp 1679585382
transform 1 0 86400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_901
timestamp 1679585382
transform 1 0 87072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_908
timestamp 1679585382
transform 1 0 87744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_915
timestamp 1679585382
transform 1 0 88416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_922
timestamp 1679585382
transform 1 0 89088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_929
timestamp 1679585382
transform 1 0 89760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_936
timestamp 1679585382
transform 1 0 90432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_943
timestamp 1679585382
transform 1 0 91104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_950
timestamp 1679585382
transform 1 0 91776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_957
timestamp 1679585382
transform 1 0 92448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_964
timestamp 1679585382
transform 1 0 93120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_971
timestamp 1679585382
transform 1 0 93792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_978
timestamp 1679585382
transform 1 0 94464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_985
timestamp 1679585382
transform 1 0 95136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_992
timestamp 1679585382
transform 1 0 95808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_999
timestamp 1679585382
transform 1 0 96480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1006
timestamp 1679585382
transform 1 0 97152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1013
timestamp 1679585382
transform 1 0 97824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1020
timestamp 1679585382
transform 1 0 98496 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_1027
timestamp 1677583704
transform 1 0 99168 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679585382
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679585382
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679585382
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_25
timestamp 1679585382
transform 1 0 2976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_32
timestamp 1679585382
transform 1 0 3648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_39
timestamp 1679581501
transform 1 0 4320 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_47
timestamp 1679585382
transform 1 0 5088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_54
timestamp 1679585382
transform 1 0 5760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_61
timestamp 1679585382
transform 1 0 6432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_68
timestamp 1679585382
transform 1 0 7104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_75
timestamp 1679585382
transform 1 0 7776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_82
timestamp 1679585382
transform 1 0 8448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_89
timestamp 1679585382
transform 1 0 9120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_96
timestamp 1679585382
transform 1 0 9792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_103
timestamp 1679585382
transform 1 0 10464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_110
timestamp 1679585382
transform 1 0 11136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_117
timestamp 1679585382
transform 1 0 11808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_124
timestamp 1679585382
transform 1 0 12480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_131
timestamp 1679585382
transform 1 0 13152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_138
timestamp 1679585382
transform 1 0 13824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_145
timestamp 1679585382
transform 1 0 14496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_152
timestamp 1679585382
transform 1 0 15168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_159
timestamp 1679585382
transform 1 0 15840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_166
timestamp 1679585382
transform 1 0 16512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_173
timestamp 1679585382
transform 1 0 17184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_180
timestamp 1679585382
transform 1 0 17856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_187
timestamp 1679585382
transform 1 0 18528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_194
timestamp 1679585382
transform 1 0 19200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_201
timestamp 1679585382
transform 1 0 19872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_208
timestamp 1679585382
transform 1 0 20544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_215
timestamp 1679585382
transform 1 0 21216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_222
timestamp 1679585382
transform 1 0 21888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_229
timestamp 1679585382
transform 1 0 22560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_236
timestamp 1679585382
transform 1 0 23232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_243
timestamp 1679585382
transform 1 0 23904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_250
timestamp 1679585382
transform 1 0 24576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_257
timestamp 1679585382
transform 1 0 25248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_264
timestamp 1679585382
transform 1 0 25920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_271
timestamp 1679585382
transform 1 0 26592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_278
timestamp 1679585382
transform 1 0 27264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_285
timestamp 1679585382
transform 1 0 27936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_292
timestamp 1679585382
transform 1 0 28608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_299
timestamp 1679585382
transform 1 0 29280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_306
timestamp 1679585382
transform 1 0 29952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_313
timestamp 1679585382
transform 1 0 30624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_320
timestamp 1679585382
transform 1 0 31296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_327
timestamp 1679585382
transform 1 0 31968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_334
timestamp 1679585382
transform 1 0 32640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_341
timestamp 1679585382
transform 1 0 33312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_348
timestamp 1679585382
transform 1 0 33984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_355
timestamp 1679585382
transform 1 0 34656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_362
timestamp 1679585382
transform 1 0 35328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_369
timestamp 1679585382
transform 1 0 36000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_376
timestamp 1679585382
transform 1 0 36672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_383
timestamp 1679585382
transform 1 0 37344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_390
timestamp 1679585382
transform 1 0 38016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_397
timestamp 1679585382
transform 1 0 38688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_404
timestamp 1679585382
transform 1 0 39360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_411
timestamp 1679585382
transform 1 0 40032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_418
timestamp 1679585382
transform 1 0 40704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_425
timestamp 1679585382
transform 1 0 41376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_432
timestamp 1679585382
transform 1 0 42048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_439
timestamp 1679585382
transform 1 0 42720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_446
timestamp 1679585382
transform 1 0 43392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_453
timestamp 1679585382
transform 1 0 44064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_460
timestamp 1679585382
transform 1 0 44736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_467
timestamp 1679585382
transform 1 0 45408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_474
timestamp 1679585382
transform 1 0 46080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_481
timestamp 1679585382
transform 1 0 46752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_488
timestamp 1679585382
transform 1 0 47424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_495
timestamp 1679585382
transform 1 0 48096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_502
timestamp 1679585382
transform 1 0 48768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_509
timestamp 1679585382
transform 1 0 49440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_516
timestamp 1679585382
transform 1 0 50112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_523
timestamp 1679585382
transform 1 0 50784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_530
timestamp 1679585382
transform 1 0 51456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_537
timestamp 1679585382
transform 1 0 52128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_544
timestamp 1679585382
transform 1 0 52800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_551
timestamp 1679585382
transform 1 0 53472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_558
timestamp 1679585382
transform 1 0 54144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_565
timestamp 1679585382
transform 1 0 54816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_572
timestamp 1679585382
transform 1 0 55488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_579
timestamp 1679585382
transform 1 0 56160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_586
timestamp 1679585382
transform 1 0 56832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_593
timestamp 1679585382
transform 1 0 57504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_600
timestamp 1679585382
transform 1 0 58176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_607
timestamp 1679585382
transform 1 0 58848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_614
timestamp 1679585382
transform 1 0 59520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_621
timestamp 1679585382
transform 1 0 60192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_628
timestamp 1679585382
transform 1 0 60864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_635
timestamp 1679585382
transform 1 0 61536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_642
timestamp 1679585382
transform 1 0 62208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_649
timestamp 1679585382
transform 1 0 62880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_656
timestamp 1679585382
transform 1 0 63552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_663
timestamp 1679585382
transform 1 0 64224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_670
timestamp 1679585382
transform 1 0 64896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_677
timestamp 1679585382
transform 1 0 65568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_684
timestamp 1679585382
transform 1 0 66240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_691
timestamp 1679585382
transform 1 0 66912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_698
timestamp 1679585382
transform 1 0 67584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_705
timestamp 1679585382
transform 1 0 68256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_712
timestamp 1679585382
transform 1 0 68928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_719
timestamp 1679585382
transform 1 0 69600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_726
timestamp 1679585382
transform 1 0 70272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_733
timestamp 1679585382
transform 1 0 70944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_740
timestamp 1679585382
transform 1 0 71616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_747
timestamp 1679585382
transform 1 0 72288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_754
timestamp 1679585382
transform 1 0 72960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_761
timestamp 1679585382
transform 1 0 73632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_768
timestamp 1679585382
transform 1 0 74304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_775
timestamp 1679585382
transform 1 0 74976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_782
timestamp 1679585382
transform 1 0 75648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_789
timestamp 1679585382
transform 1 0 76320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_796
timestamp 1679585382
transform 1 0 76992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_803
timestamp 1679585382
transform 1 0 77664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_810
timestamp 1679585382
transform 1 0 78336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_817
timestamp 1679585382
transform 1 0 79008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_824
timestamp 1679585382
transform 1 0 79680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_831
timestamp 1679585382
transform 1 0 80352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_838
timestamp 1679585382
transform 1 0 81024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_845
timestamp 1679585382
transform 1 0 81696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_852
timestamp 1679585382
transform 1 0 82368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_859
timestamp 1679585382
transform 1 0 83040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_866
timestamp 1679585382
transform 1 0 83712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_873
timestamp 1679585382
transform 1 0 84384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_880
timestamp 1679585382
transform 1 0 85056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_887
timestamp 1679585382
transform 1 0 85728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_894
timestamp 1679585382
transform 1 0 86400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_901
timestamp 1679585382
transform 1 0 87072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_908
timestamp 1679585382
transform 1 0 87744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_915
timestamp 1679585382
transform 1 0 88416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_922
timestamp 1679585382
transform 1 0 89088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_929
timestamp 1679585382
transform 1 0 89760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_936
timestamp 1679585382
transform 1 0 90432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_943
timestamp 1679585382
transform 1 0 91104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_950
timestamp 1679585382
transform 1 0 91776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_957
timestamp 1679585382
transform 1 0 92448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_964
timestamp 1679585382
transform 1 0 93120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_971
timestamp 1679585382
transform 1 0 93792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_978
timestamp 1679585382
transform 1 0 94464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_985
timestamp 1679585382
transform 1 0 95136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_992
timestamp 1679585382
transform 1 0 95808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_999
timestamp 1679585382
transform 1 0 96480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1006
timestamp 1679585382
transform 1 0 97152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1013
timestamp 1679585382
transform 1 0 97824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1020
timestamp 1679585382
transform 1 0 98496 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_1027
timestamp 1677583704
transform 1 0 99168 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679585382
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679585382
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679585382
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679585382
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679585382
transform 1 0 3648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679585382
transform 1 0 4320 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_46
timestamp 1677583704
transform 1 0 4992 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679585382
transform 1 0 5664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679585382
transform 1 0 6336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679585382
transform 1 0 7008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679585382
transform 1 0 7680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679585382
transform 1 0 8352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679585382
transform 1 0 9024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679585382
transform 1 0 9696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679585382
transform 1 0 10368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_109
timestamp 1679581501
transform 1 0 11040 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_113
timestamp 1677583704
transform 1 0 11424 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_142
timestamp 1679585382
transform 1 0 14208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_149
timestamp 1679585382
transform 1 0 14880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_156
timestamp 1679585382
transform 1 0 15552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_163
timestamp 1679585382
transform 1 0 16224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_170
timestamp 1679585382
transform 1 0 16896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_177
timestamp 1679585382
transform 1 0 17568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_184
timestamp 1679585382
transform 1 0 18240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_191
timestamp 1679585382
transform 1 0 18912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_198
timestamp 1679585382
transform 1 0 19584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_205
timestamp 1679585382
transform 1 0 20256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_212
timestamp 1679585382
transform 1 0 20928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_219
timestamp 1679585382
transform 1 0 21600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_226
timestamp 1679585382
transform 1 0 22272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_233
timestamp 1679585382
transform 1 0 22944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_240
timestamp 1679585382
transform 1 0 23616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_247
timestamp 1679585382
transform 1 0 24288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_254
timestamp 1679585382
transform 1 0 24960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_261
timestamp 1679585382
transform 1 0 25632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_268
timestamp 1679585382
transform 1 0 26304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_275
timestamp 1679585382
transform 1 0 26976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_282
timestamp 1679585382
transform 1 0 27648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_289
timestamp 1679585382
transform 1 0 28320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_296
timestamp 1679585382
transform 1 0 28992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_303
timestamp 1679585382
transform 1 0 29664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_310
timestamp 1679585382
transform 1 0 30336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_317
timestamp 1679585382
transform 1 0 31008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_324
timestamp 1679585382
transform 1 0 31680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_331
timestamp 1679585382
transform 1 0 32352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_338
timestamp 1679585382
transform 1 0 33024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_345
timestamp 1679585382
transform 1 0 33696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_352
timestamp 1679585382
transform 1 0 34368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_359
timestamp 1679585382
transform 1 0 35040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_366
timestamp 1679585382
transform 1 0 35712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_373
timestamp 1679585382
transform 1 0 36384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_380
timestamp 1679585382
transform 1 0 37056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_387
timestamp 1679585382
transform 1 0 37728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_394
timestamp 1679585382
transform 1 0 38400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_401
timestamp 1679585382
transform 1 0 39072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_408
timestamp 1679585382
transform 1 0 39744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_415
timestamp 1679585382
transform 1 0 40416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_422
timestamp 1679585382
transform 1 0 41088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_429
timestamp 1679585382
transform 1 0 41760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_436
timestamp 1679585382
transform 1 0 42432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_443
timestamp 1679585382
transform 1 0 43104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_450
timestamp 1679585382
transform 1 0 43776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_457
timestamp 1679585382
transform 1 0 44448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_464
timestamp 1679585382
transform 1 0 45120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_471
timestamp 1679585382
transform 1 0 45792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_478
timestamp 1679585382
transform 1 0 46464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_485
timestamp 1679585382
transform 1 0 47136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_492
timestamp 1679585382
transform 1 0 47808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_499
timestamp 1679585382
transform 1 0 48480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_506
timestamp 1679585382
transform 1 0 49152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_513
timestamp 1679585382
transform 1 0 49824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_520
timestamp 1679585382
transform 1 0 50496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_527
timestamp 1679585382
transform 1 0 51168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_534
timestamp 1679585382
transform 1 0 51840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_541
timestamp 1679585382
transform 1 0 52512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_548
timestamp 1679585382
transform 1 0 53184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_555
timestamp 1679585382
transform 1 0 53856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_562
timestamp 1679585382
transform 1 0 54528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_569
timestamp 1679585382
transform 1 0 55200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_576
timestamp 1679585382
transform 1 0 55872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_583
timestamp 1679585382
transform 1 0 56544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_590
timestamp 1679585382
transform 1 0 57216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_597
timestamp 1679585382
transform 1 0 57888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_604
timestamp 1679585382
transform 1 0 58560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_611
timestamp 1679585382
transform 1 0 59232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_618
timestamp 1679585382
transform 1 0 59904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_625
timestamp 1679585382
transform 1 0 60576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_632
timestamp 1679585382
transform 1 0 61248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_639
timestamp 1679585382
transform 1 0 61920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_646
timestamp 1679585382
transform 1 0 62592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_653
timestamp 1679585382
transform 1 0 63264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_660
timestamp 1679585382
transform 1 0 63936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_667
timestamp 1679585382
transform 1 0 64608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_674
timestamp 1679585382
transform 1 0 65280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_681
timestamp 1679585382
transform 1 0 65952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_688
timestamp 1679585382
transform 1 0 66624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_695
timestamp 1679585382
transform 1 0 67296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_702
timestamp 1679585382
transform 1 0 67968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_709
timestamp 1679585382
transform 1 0 68640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_716
timestamp 1679585382
transform 1 0 69312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_723
timestamp 1679585382
transform 1 0 69984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_730
timestamp 1679585382
transform 1 0 70656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_737
timestamp 1679585382
transform 1 0 71328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_744
timestamp 1679585382
transform 1 0 72000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_751
timestamp 1679585382
transform 1 0 72672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_758
timestamp 1679585382
transform 1 0 73344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_765
timestamp 1679585382
transform 1 0 74016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_772
timestamp 1679585382
transform 1 0 74688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_779
timestamp 1679585382
transform 1 0 75360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_786
timestamp 1679585382
transform 1 0 76032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_793
timestamp 1679585382
transform 1 0 76704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_800
timestamp 1679585382
transform 1 0 77376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_807
timestamp 1679585382
transform 1 0 78048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_814
timestamp 1679585382
transform 1 0 78720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_821
timestamp 1679585382
transform 1 0 79392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_828
timestamp 1679585382
transform 1 0 80064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_835
timestamp 1679585382
transform 1 0 80736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_842
timestamp 1679585382
transform 1 0 81408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_849
timestamp 1679585382
transform 1 0 82080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_856
timestamp 1679585382
transform 1 0 82752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_863
timestamp 1679585382
transform 1 0 83424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_870
timestamp 1679585382
transform 1 0 84096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_877
timestamp 1679585382
transform 1 0 84768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_884
timestamp 1679585382
transform 1 0 85440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_891
timestamp 1679585382
transform 1 0 86112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_898
timestamp 1679585382
transform 1 0 86784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_905
timestamp 1679585382
transform 1 0 87456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_912
timestamp 1679585382
transform 1 0 88128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_919
timestamp 1679585382
transform 1 0 88800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_926
timestamp 1679585382
transform 1 0 89472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_933
timestamp 1679585382
transform 1 0 90144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_940
timestamp 1679585382
transform 1 0 90816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_947
timestamp 1679585382
transform 1 0 91488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_954
timestamp 1679585382
transform 1 0 92160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_961
timestamp 1679585382
transform 1 0 92832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_968
timestamp 1679585382
transform 1 0 93504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_975
timestamp 1679585382
transform 1 0 94176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_982
timestamp 1679585382
transform 1 0 94848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_989
timestamp 1679585382
transform 1 0 95520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_996
timestamp 1679585382
transform 1 0 96192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1003
timestamp 1679585382
transform 1 0 96864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1010
timestamp 1679585382
transform 1 0 97536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1017
timestamp 1679585382
transform 1 0 98208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_1024
timestamp 1679581501
transform 1 0 98880 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_1028
timestamp 1677583258
transform 1 0 99264 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679585382
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679585382
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_18
timestamp 1677583704
transform 1 0 2304 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_20
timestamp 1677583258
transform 1 0 2496 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_25
timestamp 1679585382
transform 1 0 2976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_32
timestamp 1679585382
transform 1 0 3648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_39
timestamp 1679585382
transform 1 0 4320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_46
timestamp 1679585382
transform 1 0 4992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_53
timestamp 1679585382
transform 1 0 5664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_60
timestamp 1679585382
transform 1 0 6336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_67
timestamp 1679585382
transform 1 0 7008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_74
timestamp 1679585382
transform 1 0 7680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_92
timestamp 1679585382
transform 1 0 9408 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_99
timestamp 1677583704
transform 1 0 10080 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_101
timestamp 1677583258
transform 1 0 10272 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_111
timestamp 1677583258
transform 1 0 11232 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_125
timestamp 1679585382
transform 1 0 12576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_132
timestamp 1679585382
transform 1 0 13248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_139
timestamp 1679585382
transform 1 0 13920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_146
timestamp 1679585382
transform 1 0 14592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_153
timestamp 1679585382
transform 1 0 15264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_160
timestamp 1679585382
transform 1 0 15936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_167
timestamp 1679585382
transform 1 0 16608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_174
timestamp 1679585382
transform 1 0 17280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_181
timestamp 1679585382
transform 1 0 17952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_188
timestamp 1679585382
transform 1 0 18624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_195
timestamp 1679585382
transform 1 0 19296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_202
timestamp 1679585382
transform 1 0 19968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_209
timestamp 1679585382
transform 1 0 20640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_216
timestamp 1679585382
transform 1 0 21312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_223
timestamp 1679585382
transform 1 0 21984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_230
timestamp 1679585382
transform 1 0 22656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_237
timestamp 1679585382
transform 1 0 23328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_244
timestamp 1679585382
transform 1 0 24000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_251
timestamp 1679585382
transform 1 0 24672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_258
timestamp 1679585382
transform 1 0 25344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_265
timestamp 1679585382
transform 1 0 26016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_272
timestamp 1679585382
transform 1 0 26688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_279
timestamp 1679585382
transform 1 0 27360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_286
timestamp 1679585382
transform 1 0 28032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_293
timestamp 1679585382
transform 1 0 28704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_300
timestamp 1679585382
transform 1 0 29376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_307
timestamp 1679585382
transform 1 0 30048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_314
timestamp 1679585382
transform 1 0 30720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_321
timestamp 1679585382
transform 1 0 31392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_328
timestamp 1679585382
transform 1 0 32064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_335
timestamp 1679585382
transform 1 0 32736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_342
timestamp 1679585382
transform 1 0 33408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_349
timestamp 1679585382
transform 1 0 34080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_356
timestamp 1679585382
transform 1 0 34752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_363
timestamp 1679585382
transform 1 0 35424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_370
timestamp 1679585382
transform 1 0 36096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_377
timestamp 1679585382
transform 1 0 36768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_384
timestamp 1679585382
transform 1 0 37440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_391
timestamp 1679585382
transform 1 0 38112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_398
timestamp 1679585382
transform 1 0 38784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_405
timestamp 1679585382
transform 1 0 39456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_412
timestamp 1679585382
transform 1 0 40128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_419
timestamp 1679585382
transform 1 0 40800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_426
timestamp 1679585382
transform 1 0 41472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_433
timestamp 1679585382
transform 1 0 42144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_440
timestamp 1679585382
transform 1 0 42816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_447
timestamp 1679585382
transform 1 0 43488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_454
timestamp 1679585382
transform 1 0 44160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_461
timestamp 1679585382
transform 1 0 44832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_468
timestamp 1679585382
transform 1 0 45504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_475
timestamp 1679585382
transform 1 0 46176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_482
timestamp 1679585382
transform 1 0 46848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_489
timestamp 1679585382
transform 1 0 47520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_496
timestamp 1679585382
transform 1 0 48192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_503
timestamp 1679585382
transform 1 0 48864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_510
timestamp 1679585382
transform 1 0 49536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_517
timestamp 1679585382
transform 1 0 50208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_524
timestamp 1679585382
transform 1 0 50880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_531
timestamp 1679585382
transform 1 0 51552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_538
timestamp 1679585382
transform 1 0 52224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_545
timestamp 1679585382
transform 1 0 52896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_552
timestamp 1679585382
transform 1 0 53568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_559
timestamp 1679585382
transform 1 0 54240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_566
timestamp 1679585382
transform 1 0 54912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_573
timestamp 1679585382
transform 1 0 55584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_580
timestamp 1679585382
transform 1 0 56256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_587
timestamp 1679585382
transform 1 0 56928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_594
timestamp 1679585382
transform 1 0 57600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_601
timestamp 1679585382
transform 1 0 58272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_608
timestamp 1679585382
transform 1 0 58944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_615
timestamp 1679585382
transform 1 0 59616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_622
timestamp 1679585382
transform 1 0 60288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_629
timestamp 1679585382
transform 1 0 60960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_636
timestamp 1679585382
transform 1 0 61632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_643
timestamp 1679585382
transform 1 0 62304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_650
timestamp 1679585382
transform 1 0 62976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_657
timestamp 1679585382
transform 1 0 63648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_664
timestamp 1679585382
transform 1 0 64320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_671
timestamp 1679585382
transform 1 0 64992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_678
timestamp 1679585382
transform 1 0 65664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_685
timestamp 1679585382
transform 1 0 66336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_692
timestamp 1679585382
transform 1 0 67008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_699
timestamp 1679585382
transform 1 0 67680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_706
timestamp 1679585382
transform 1 0 68352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_713
timestamp 1679585382
transform 1 0 69024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_720
timestamp 1679585382
transform 1 0 69696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_727
timestamp 1679585382
transform 1 0 70368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_734
timestamp 1679585382
transform 1 0 71040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_741
timestamp 1679585382
transform 1 0 71712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_748
timestamp 1679585382
transform 1 0 72384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_755
timestamp 1679585382
transform 1 0 73056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_762
timestamp 1679585382
transform 1 0 73728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_769
timestamp 1679585382
transform 1 0 74400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_776
timestamp 1679585382
transform 1 0 75072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_783
timestamp 1679585382
transform 1 0 75744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_790
timestamp 1679585382
transform 1 0 76416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_797
timestamp 1679585382
transform 1 0 77088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_804
timestamp 1679585382
transform 1 0 77760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_811
timestamp 1679585382
transform 1 0 78432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_818
timestamp 1679585382
transform 1 0 79104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_825
timestamp 1679585382
transform 1 0 79776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_832
timestamp 1679585382
transform 1 0 80448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_839
timestamp 1679585382
transform 1 0 81120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_846
timestamp 1679585382
transform 1 0 81792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_853
timestamp 1679585382
transform 1 0 82464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_860
timestamp 1679585382
transform 1 0 83136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_867
timestamp 1679585382
transform 1 0 83808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_874
timestamp 1679585382
transform 1 0 84480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_881
timestamp 1679585382
transform 1 0 85152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_888
timestamp 1679585382
transform 1 0 85824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_895
timestamp 1679585382
transform 1 0 86496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_902
timestamp 1679585382
transform 1 0 87168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_909
timestamp 1679585382
transform 1 0 87840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_916
timestamp 1679585382
transform 1 0 88512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_923
timestamp 1679585382
transform 1 0 89184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_930
timestamp 1679585382
transform 1 0 89856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_937
timestamp 1679585382
transform 1 0 90528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_944
timestamp 1679585382
transform 1 0 91200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_951
timestamp 1679585382
transform 1 0 91872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_958
timestamp 1679585382
transform 1 0 92544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_965
timestamp 1679585382
transform 1 0 93216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_972
timestamp 1679585382
transform 1 0 93888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_979
timestamp 1679585382
transform 1 0 94560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_986
timestamp 1679585382
transform 1 0 95232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_993
timestamp 1679585382
transform 1 0 95904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1000
timestamp 1679585382
transform 1 0 96576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1007
timestamp 1679585382
transform 1 0 97248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1014
timestamp 1679585382
transform 1 0 97920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1021
timestamp 1679585382
transform 1 0 98592 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_1028
timestamp 1677583258
transform 1 0 99264 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679585382
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_11
timestamp 1679581501
transform 1 0 1632 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_15
timestamp 1677583704
transform 1 0 2016 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679585382
transform 1 0 2976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679585382
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679585382
transform 1 0 4320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_46
timestamp 1679585382
transform 1 0 4992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_53
timestamp 1679585382
transform 1 0 5664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_60
timestamp 1679581501
transform 1 0 6336 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_64
timestamp 1677583258
transform 1 0 6720 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_72
timestamp 1679585382
transform 1 0 7488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_79
timestamp 1679585382
transform 1 0 8160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_86
timestamp 1679585382
transform 1 0 8832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_93
timestamp 1679585382
transform 1 0 9504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_100
timestamp 1679585382
transform 1 0 10176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_107
timestamp 1679585382
transform 1 0 10848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_114
timestamp 1679585382
transform 1 0 11520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_121
timestamp 1679585382
transform 1 0 12192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_128
timestamp 1679585382
transform 1 0 12864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_135
timestamp 1679585382
transform 1 0 13536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_142
timestamp 1679585382
transform 1 0 14208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_149
timestamp 1679585382
transform 1 0 14880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_156
timestamp 1679585382
transform 1 0 15552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_163
timestamp 1679585382
transform 1 0 16224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_170
timestamp 1679585382
transform 1 0 16896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_177
timestamp 1679585382
transform 1 0 17568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_184
timestamp 1679585382
transform 1 0 18240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_191
timestamp 1679585382
transform 1 0 18912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_198
timestamp 1679585382
transform 1 0 19584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_205
timestamp 1679585382
transform 1 0 20256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_212
timestamp 1679585382
transform 1 0 20928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_219
timestamp 1679585382
transform 1 0 21600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_226
timestamp 1679585382
transform 1 0 22272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_233
timestamp 1679585382
transform 1 0 22944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_240
timestamp 1679585382
transform 1 0 23616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_247
timestamp 1679585382
transform 1 0 24288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_254
timestamp 1679585382
transform 1 0 24960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_261
timestamp 1679585382
transform 1 0 25632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_268
timestamp 1679585382
transform 1 0 26304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_275
timestamp 1679585382
transform 1 0 26976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_282
timestamp 1679585382
transform 1 0 27648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_289
timestamp 1679585382
transform 1 0 28320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_296
timestamp 1679585382
transform 1 0 28992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_303
timestamp 1679585382
transform 1 0 29664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_310
timestamp 1679585382
transform 1 0 30336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_317
timestamp 1679585382
transform 1 0 31008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_324
timestamp 1679585382
transform 1 0 31680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_331
timestamp 1679585382
transform 1 0 32352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_338
timestamp 1679585382
transform 1 0 33024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_345
timestamp 1679585382
transform 1 0 33696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_352
timestamp 1679585382
transform 1 0 34368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_359
timestamp 1679585382
transform 1 0 35040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_366
timestamp 1679585382
transform 1 0 35712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_373
timestamp 1679585382
transform 1 0 36384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_380
timestamp 1679585382
transform 1 0 37056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_387
timestamp 1679585382
transform 1 0 37728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_394
timestamp 1679585382
transform 1 0 38400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_401
timestamp 1679585382
transform 1 0 39072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_408
timestamp 1679585382
transform 1 0 39744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_415
timestamp 1679585382
transform 1 0 40416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_422
timestamp 1679585382
transform 1 0 41088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_429
timestamp 1679585382
transform 1 0 41760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_436
timestamp 1679585382
transform 1 0 42432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_443
timestamp 1679585382
transform 1 0 43104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_450
timestamp 1679585382
transform 1 0 43776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_457
timestamp 1679585382
transform 1 0 44448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_464
timestamp 1679585382
transform 1 0 45120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_471
timestamp 1679585382
transform 1 0 45792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_478
timestamp 1679585382
transform 1 0 46464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_485
timestamp 1679585382
transform 1 0 47136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_492
timestamp 1679585382
transform 1 0 47808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_499
timestamp 1679585382
transform 1 0 48480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_506
timestamp 1679585382
transform 1 0 49152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_513
timestamp 1679585382
transform 1 0 49824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_520
timestamp 1679585382
transform 1 0 50496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_527
timestamp 1679585382
transform 1 0 51168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_534
timestamp 1679585382
transform 1 0 51840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_541
timestamp 1679585382
transform 1 0 52512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_548
timestamp 1679585382
transform 1 0 53184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_555
timestamp 1679585382
transform 1 0 53856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_562
timestamp 1679585382
transform 1 0 54528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_569
timestamp 1679585382
transform 1 0 55200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_576
timestamp 1679585382
transform 1 0 55872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_583
timestamp 1679585382
transform 1 0 56544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_590
timestamp 1679585382
transform 1 0 57216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_597
timestamp 1679585382
transform 1 0 57888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_604
timestamp 1679585382
transform 1 0 58560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_611
timestamp 1679585382
transform 1 0 59232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_618
timestamp 1679585382
transform 1 0 59904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_625
timestamp 1679585382
transform 1 0 60576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_632
timestamp 1679585382
transform 1 0 61248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_639
timestamp 1679585382
transform 1 0 61920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_646
timestamp 1679585382
transform 1 0 62592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_653
timestamp 1679585382
transform 1 0 63264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_660
timestamp 1679585382
transform 1 0 63936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_667
timestamp 1679585382
transform 1 0 64608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_674
timestamp 1679585382
transform 1 0 65280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_681
timestamp 1679585382
transform 1 0 65952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_688
timestamp 1679585382
transform 1 0 66624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_695
timestamp 1679585382
transform 1 0 67296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_702
timestamp 1679585382
transform 1 0 67968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_709
timestamp 1679585382
transform 1 0 68640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_716
timestamp 1679585382
transform 1 0 69312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_723
timestamp 1679585382
transform 1 0 69984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_730
timestamp 1679585382
transform 1 0 70656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_737
timestamp 1679585382
transform 1 0 71328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_744
timestamp 1679585382
transform 1 0 72000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_751
timestamp 1679585382
transform 1 0 72672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_758
timestamp 1679585382
transform 1 0 73344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_765
timestamp 1679585382
transform 1 0 74016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_772
timestamp 1679585382
transform 1 0 74688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_779
timestamp 1679585382
transform 1 0 75360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_786
timestamp 1679585382
transform 1 0 76032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_793
timestamp 1679585382
transform 1 0 76704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_800
timestamp 1679585382
transform 1 0 77376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_807
timestamp 1679585382
transform 1 0 78048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_814
timestamp 1679585382
transform 1 0 78720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_821
timestamp 1679585382
transform 1 0 79392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_828
timestamp 1679585382
transform 1 0 80064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_835
timestamp 1679585382
transform 1 0 80736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_842
timestamp 1679585382
transform 1 0 81408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_849
timestamp 1679585382
transform 1 0 82080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_856
timestamp 1679585382
transform 1 0 82752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_863
timestamp 1679585382
transform 1 0 83424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_870
timestamp 1679585382
transform 1 0 84096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_877
timestamp 1679585382
transform 1 0 84768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_884
timestamp 1679585382
transform 1 0 85440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_891
timestamp 1679585382
transform 1 0 86112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_898
timestamp 1679585382
transform 1 0 86784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_905
timestamp 1679585382
transform 1 0 87456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_912
timestamp 1679585382
transform 1 0 88128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_919
timestamp 1679585382
transform 1 0 88800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_926
timestamp 1679585382
transform 1 0 89472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_933
timestamp 1679585382
transform 1 0 90144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_940
timestamp 1679585382
transform 1 0 90816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_947
timestamp 1679585382
transform 1 0 91488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_954
timestamp 1679585382
transform 1 0 92160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_961
timestamp 1679585382
transform 1 0 92832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_968
timestamp 1679585382
transform 1 0 93504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_975
timestamp 1679585382
transform 1 0 94176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_982
timestamp 1679585382
transform 1 0 94848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_989
timestamp 1679585382
transform 1 0 95520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_996
timestamp 1679585382
transform 1 0 96192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1003
timestamp 1679585382
transform 1 0 96864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1010
timestamp 1679585382
transform 1 0 97536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1017
timestamp 1679585382
transform 1 0 98208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_1024
timestamp 1679581501
transform 1 0 98880 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_1028
timestamp 1677583258
transform 1 0 99264 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679585382
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679585382
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_18
timestamp 1677583704
transform 1 0 2304 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_20
timestamp 1677583258
transform 1 0 2496 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679585382
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_32
timestamp 1679581501
transform 1 0 3648 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_39
timestamp 1679585382
transform 1 0 4320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_46
timestamp 1679585382
transform 1 0 4992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679585382
transform 1 0 5664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679585382
transform 1 0 6336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_67
timestamp 1679585382
transform 1 0 7008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_74
timestamp 1679585382
transform 1 0 7680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_81
timestamp 1679585382
transform 1 0 8352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_88
timestamp 1679585382
transform 1 0 9024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_95
timestamp 1679581501
transform 1 0 9696 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_99
timestamp 1677583704
transform 1 0 10080 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_126
timestamp 1679585382
transform 1 0 12672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_133
timestamp 1679585382
transform 1 0 13344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_140
timestamp 1679585382
transform 1 0 14016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_147
timestamp 1679585382
transform 1 0 14688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_154
timestamp 1679585382
transform 1 0 15360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_161
timestamp 1679585382
transform 1 0 16032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_168
timestamp 1679585382
transform 1 0 16704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_175
timestamp 1679585382
transform 1 0 17376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_182
timestamp 1679585382
transform 1 0 18048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679585382
transform 1 0 18720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_196
timestamp 1679585382
transform 1 0 19392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_203
timestamp 1679585382
transform 1 0 20064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_210
timestamp 1679585382
transform 1 0 20736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_217
timestamp 1679585382
transform 1 0 21408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_224
timestamp 1679585382
transform 1 0 22080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_231
timestamp 1679585382
transform 1 0 22752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_238
timestamp 1679585382
transform 1 0 23424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_245
timestamp 1679585382
transform 1 0 24096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_252
timestamp 1679585382
transform 1 0 24768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_259
timestamp 1679585382
transform 1 0 25440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_266
timestamp 1679585382
transform 1 0 26112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_273
timestamp 1679585382
transform 1 0 26784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_280
timestamp 1679585382
transform 1 0 27456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_287
timestamp 1679585382
transform 1 0 28128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_294
timestamp 1679585382
transform 1 0 28800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_301
timestamp 1679585382
transform 1 0 29472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_308
timestamp 1679585382
transform 1 0 30144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_315
timestamp 1679585382
transform 1 0 30816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_322
timestamp 1679585382
transform 1 0 31488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_329
timestamp 1679585382
transform 1 0 32160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_336
timestamp 1679585382
transform 1 0 32832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_343
timestamp 1679585382
transform 1 0 33504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_350
timestamp 1679585382
transform 1 0 34176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_357
timestamp 1679585382
transform 1 0 34848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_364
timestamp 1679585382
transform 1 0 35520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_371
timestamp 1679585382
transform 1 0 36192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_378
timestamp 1679585382
transform 1 0 36864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_385
timestamp 1679585382
transform 1 0 37536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_392
timestamp 1679585382
transform 1 0 38208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_399
timestamp 1679585382
transform 1 0 38880 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_406
timestamp 1679585382
transform 1 0 39552 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_413
timestamp 1679585382
transform 1 0 40224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_420
timestamp 1679585382
transform 1 0 40896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_427
timestamp 1679585382
transform 1 0 41568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_434
timestamp 1679585382
transform 1 0 42240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_441
timestamp 1679585382
transform 1 0 42912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_448
timestamp 1679585382
transform 1 0 43584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_455
timestamp 1679585382
transform 1 0 44256 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_462
timestamp 1679585382
transform 1 0 44928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_469
timestamp 1679585382
transform 1 0 45600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_476
timestamp 1679585382
transform 1 0 46272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_483
timestamp 1679585382
transform 1 0 46944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_490
timestamp 1679585382
transform 1 0 47616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_497
timestamp 1679585382
transform 1 0 48288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_504
timestamp 1679585382
transform 1 0 48960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_511
timestamp 1679585382
transform 1 0 49632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_518
timestamp 1679585382
transform 1 0 50304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_525
timestamp 1679585382
transform 1 0 50976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_532
timestamp 1679585382
transform 1 0 51648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_539
timestamp 1679585382
transform 1 0 52320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_546
timestamp 1679585382
transform 1 0 52992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_553
timestamp 1679585382
transform 1 0 53664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_560
timestamp 1679585382
transform 1 0 54336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_567
timestamp 1679585382
transform 1 0 55008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_574
timestamp 1679585382
transform 1 0 55680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_581
timestamp 1679585382
transform 1 0 56352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_588
timestamp 1679585382
transform 1 0 57024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_595
timestamp 1679585382
transform 1 0 57696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_602
timestamp 1679585382
transform 1 0 58368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_609
timestamp 1679585382
transform 1 0 59040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_616
timestamp 1679585382
transform 1 0 59712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_623
timestamp 1679585382
transform 1 0 60384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_630
timestamp 1679585382
transform 1 0 61056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_637
timestamp 1679585382
transform 1 0 61728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_644
timestamp 1679585382
transform 1 0 62400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_651
timestamp 1679585382
transform 1 0 63072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_658
timestamp 1679585382
transform 1 0 63744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_665
timestamp 1679585382
transform 1 0 64416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_672
timestamp 1679585382
transform 1 0 65088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_679
timestamp 1679585382
transform 1 0 65760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_686
timestamp 1679585382
transform 1 0 66432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_693
timestamp 1679585382
transform 1 0 67104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_700
timestamp 1679585382
transform 1 0 67776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_707
timestamp 1679585382
transform 1 0 68448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_714
timestamp 1679585382
transform 1 0 69120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_721
timestamp 1679585382
transform 1 0 69792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_728
timestamp 1679585382
transform 1 0 70464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_735
timestamp 1679585382
transform 1 0 71136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_742
timestamp 1679585382
transform 1 0 71808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_749
timestamp 1679585382
transform 1 0 72480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_756
timestamp 1679585382
transform 1 0 73152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_763
timestamp 1679585382
transform 1 0 73824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_770
timestamp 1679585382
transform 1 0 74496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_777
timestamp 1679585382
transform 1 0 75168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_784
timestamp 1679585382
transform 1 0 75840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_791
timestamp 1679585382
transform 1 0 76512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_798
timestamp 1679585382
transform 1 0 77184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_805
timestamp 1679585382
transform 1 0 77856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_812
timestamp 1679585382
transform 1 0 78528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_819
timestamp 1679585382
transform 1 0 79200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_826
timestamp 1679585382
transform 1 0 79872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_833
timestamp 1679585382
transform 1 0 80544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_840
timestamp 1679585382
transform 1 0 81216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_847
timestamp 1679585382
transform 1 0 81888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_854
timestamp 1679585382
transform 1 0 82560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_861
timestamp 1679585382
transform 1 0 83232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_868
timestamp 1679585382
transform 1 0 83904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_875
timestamp 1679585382
transform 1 0 84576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_882
timestamp 1679585382
transform 1 0 85248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_889
timestamp 1679585382
transform 1 0 85920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_896
timestamp 1679585382
transform 1 0 86592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_903
timestamp 1679585382
transform 1 0 87264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_910
timestamp 1679585382
transform 1 0 87936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_917
timestamp 1679585382
transform 1 0 88608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_924
timestamp 1679585382
transform 1 0 89280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_931
timestamp 1679585382
transform 1 0 89952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_938
timestamp 1679585382
transform 1 0 90624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_945
timestamp 1679585382
transform 1 0 91296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_952
timestamp 1679585382
transform 1 0 91968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_959
timestamp 1679585382
transform 1 0 92640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_966
timestamp 1679585382
transform 1 0 93312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_973
timestamp 1679585382
transform 1 0 93984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_980
timestamp 1679585382
transform 1 0 94656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_987
timestamp 1679585382
transform 1 0 95328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_994
timestamp 1679585382
transform 1 0 96000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1001
timestamp 1679585382
transform 1 0 96672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1008
timestamp 1679585382
transform 1 0 97344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1015
timestamp 1679585382
transform 1 0 98016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1022
timestamp 1679585382
transform 1 0 98688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679585382
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679585382
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679585382
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_25
timestamp 1679585382
transform 1 0 2976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_32
timestamp 1679585382
transform 1 0 3648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_39
timestamp 1679585382
transform 1 0 4320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_46
timestamp 1679585382
transform 1 0 4992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_53
timestamp 1679585382
transform 1 0 5664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_60
timestamp 1679585382
transform 1 0 6336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_67
timestamp 1679585382
transform 1 0 7008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_74
timestamp 1679585382
transform 1 0 7680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_81
timestamp 1679585382
transform 1 0 8352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_88
timestamp 1679585382
transform 1 0 9024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_95
timestamp 1679585382
transform 1 0 9696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_102
timestamp 1679585382
transform 1 0 10368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_109
timestamp 1679585382
transform 1 0 11040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_116
timestamp 1679585382
transform 1 0 11712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_123
timestamp 1679585382
transform 1 0 12384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_130
timestamp 1679585382
transform 1 0 13056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_137
timestamp 1679585382
transform 1 0 13728 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_144
timestamp 1677583258
transform 1 0 14400 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_149
timestamp 1679585382
transform 1 0 14880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_156
timestamp 1679585382
transform 1 0 15552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_163
timestamp 1679585382
transform 1 0 16224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_170
timestamp 1679585382
transform 1 0 16896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_177
timestamp 1679585382
transform 1 0 17568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_184
timestamp 1679585382
transform 1 0 18240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_191
timestamp 1679585382
transform 1 0 18912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_198
timestamp 1679585382
transform 1 0 19584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_205
timestamp 1679585382
transform 1 0 20256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_212
timestamp 1679585382
transform 1 0 20928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_219
timestamp 1679585382
transform 1 0 21600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_226
timestamp 1679585382
transform 1 0 22272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_233
timestamp 1679585382
transform 1 0 22944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_240
timestamp 1679585382
transform 1 0 23616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_247
timestamp 1679585382
transform 1 0 24288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_254
timestamp 1679585382
transform 1 0 24960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_261
timestamp 1679585382
transform 1 0 25632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_268
timestamp 1679585382
transform 1 0 26304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_275
timestamp 1679585382
transform 1 0 26976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_282
timestamp 1679585382
transform 1 0 27648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_289
timestamp 1679585382
transform 1 0 28320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_296
timestamp 1679585382
transform 1 0 28992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_303
timestamp 1679585382
transform 1 0 29664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_310
timestamp 1679585382
transform 1 0 30336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_317
timestamp 1679585382
transform 1 0 31008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_324
timestamp 1679585382
transform 1 0 31680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_331
timestamp 1679585382
transform 1 0 32352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_338
timestamp 1679585382
transform 1 0 33024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_345
timestamp 1679585382
transform 1 0 33696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_352
timestamp 1679585382
transform 1 0 34368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_359
timestamp 1679585382
transform 1 0 35040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_366
timestamp 1679585382
transform 1 0 35712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_373
timestamp 1679585382
transform 1 0 36384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_380
timestamp 1679585382
transform 1 0 37056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_387
timestamp 1679585382
transform 1 0 37728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_394
timestamp 1679585382
transform 1 0 38400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_401
timestamp 1679585382
transform 1 0 39072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_408
timestamp 1679585382
transform 1 0 39744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_415
timestamp 1679585382
transform 1 0 40416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_422
timestamp 1679585382
transform 1 0 41088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_429
timestamp 1679585382
transform 1 0 41760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_436
timestamp 1679585382
transform 1 0 42432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_443
timestamp 1679585382
transform 1 0 43104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_450
timestamp 1679585382
transform 1 0 43776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_457
timestamp 1679585382
transform 1 0 44448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_464
timestamp 1679585382
transform 1 0 45120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_471
timestamp 1679585382
transform 1 0 45792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_478
timestamp 1679585382
transform 1 0 46464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_485
timestamp 1679585382
transform 1 0 47136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_492
timestamp 1679585382
transform 1 0 47808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_499
timestamp 1679585382
transform 1 0 48480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_506
timestamp 1679585382
transform 1 0 49152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_513
timestamp 1679585382
transform 1 0 49824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_520
timestamp 1679585382
transform 1 0 50496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_527
timestamp 1679585382
transform 1 0 51168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_534
timestamp 1679585382
transform 1 0 51840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_541
timestamp 1679585382
transform 1 0 52512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_548
timestamp 1679585382
transform 1 0 53184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_555
timestamp 1679585382
transform 1 0 53856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_562
timestamp 1679585382
transform 1 0 54528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_569
timestamp 1679585382
transform 1 0 55200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_576
timestamp 1679585382
transform 1 0 55872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_583
timestamp 1679585382
transform 1 0 56544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_590
timestamp 1679585382
transform 1 0 57216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_597
timestamp 1679585382
transform 1 0 57888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_604
timestamp 1679585382
transform 1 0 58560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_611
timestamp 1679585382
transform 1 0 59232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_618
timestamp 1679585382
transform 1 0 59904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_625
timestamp 1679585382
transform 1 0 60576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_632
timestamp 1679585382
transform 1 0 61248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_639
timestamp 1679585382
transform 1 0 61920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_646
timestamp 1679585382
transform 1 0 62592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_653
timestamp 1679585382
transform 1 0 63264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_660
timestamp 1679585382
transform 1 0 63936 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_667
timestamp 1679585382
transform 1 0 64608 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_674
timestamp 1679585382
transform 1 0 65280 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_681
timestamp 1679585382
transform 1 0 65952 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_688
timestamp 1679585382
transform 1 0 66624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_695
timestamp 1679585382
transform 1 0 67296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_702
timestamp 1679585382
transform 1 0 67968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_709
timestamp 1679585382
transform 1 0 68640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_716
timestamp 1679585382
transform 1 0 69312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_723
timestamp 1679585382
transform 1 0 69984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_730
timestamp 1679585382
transform 1 0 70656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_737
timestamp 1679585382
transform 1 0 71328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_744
timestamp 1679585382
transform 1 0 72000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_751
timestamp 1679585382
transform 1 0 72672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_758
timestamp 1679585382
transform 1 0 73344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_765
timestamp 1679585382
transform 1 0 74016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_772
timestamp 1679585382
transform 1 0 74688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_779
timestamp 1679585382
transform 1 0 75360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_786
timestamp 1679585382
transform 1 0 76032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_793
timestamp 1679585382
transform 1 0 76704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_800
timestamp 1679585382
transform 1 0 77376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_807
timestamp 1679585382
transform 1 0 78048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_814
timestamp 1679585382
transform 1 0 78720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_821
timestamp 1679585382
transform 1 0 79392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_828
timestamp 1679585382
transform 1 0 80064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_835
timestamp 1679585382
transform 1 0 80736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_842
timestamp 1679585382
transform 1 0 81408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_849
timestamp 1679585382
transform 1 0 82080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_856
timestamp 1679585382
transform 1 0 82752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_863
timestamp 1679585382
transform 1 0 83424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_870
timestamp 1679585382
transform 1 0 84096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_877
timestamp 1679585382
transform 1 0 84768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_884
timestamp 1679585382
transform 1 0 85440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_891
timestamp 1679585382
transform 1 0 86112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_898
timestamp 1679585382
transform 1 0 86784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_905
timestamp 1679585382
transform 1 0 87456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_912
timestamp 1679585382
transform 1 0 88128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_919
timestamp 1679585382
transform 1 0 88800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_926
timestamp 1679585382
transform 1 0 89472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_933
timestamp 1679585382
transform 1 0 90144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_940
timestamp 1679585382
transform 1 0 90816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_947
timestamp 1679585382
transform 1 0 91488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_954
timestamp 1679585382
transform 1 0 92160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_961
timestamp 1679585382
transform 1 0 92832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_968
timestamp 1679585382
transform 1 0 93504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_975
timestamp 1679585382
transform 1 0 94176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_982
timestamp 1679585382
transform 1 0 94848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_989
timestamp 1679585382
transform 1 0 95520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_996
timestamp 1679585382
transform 1 0 96192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1003
timestamp 1679585382
transform 1 0 96864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1010
timestamp 1679585382
transform 1 0 97536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1017
timestamp 1679585382
transform 1 0 98208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_1024
timestamp 1679581501
transform 1 0 98880 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_1028
timestamp 1677583258
transform 1 0 99264 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679585382
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679585382
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_18
timestamp 1679585382
transform 1 0 2304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_25
timestamp 1679585382
transform 1 0 2976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_32
timestamp 1679585382
transform 1 0 3648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_39
timestamp 1679585382
transform 1 0 4320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679585382
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_53
timestamp 1679585382
transform 1 0 5664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_60
timestamp 1679585382
transform 1 0 6336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_67
timestamp 1679585382
transform 1 0 7008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_74
timestamp 1679585382
transform 1 0 7680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_81
timestamp 1679585382
transform 1 0 8352 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_88
timestamp 1677583258
transform 1 0 9024 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_99
timestamp 1679585382
transform 1 0 10080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_106
timestamp 1679585382
transform 1 0 10752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_113
timestamp 1679585382
transform 1 0 11424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_120
timestamp 1679585382
transform 1 0 12096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_127
timestamp 1679585382
transform 1 0 12768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_134
timestamp 1679581501
transform 1 0 13440 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_138
timestamp 1677583704
transform 1 0 13824 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_167
timestamp 1679585382
transform 1 0 16608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_174
timestamp 1679585382
transform 1 0 17280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_181
timestamp 1679585382
transform 1 0 17952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_188
timestamp 1679585382
transform 1 0 18624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_195
timestamp 1679585382
transform 1 0 19296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_202
timestamp 1679585382
transform 1 0 19968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_209
timestamp 1679585382
transform 1 0 20640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_216
timestamp 1679585382
transform 1 0 21312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_223
timestamp 1679585382
transform 1 0 21984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_230
timestamp 1679585382
transform 1 0 22656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_237
timestamp 1679585382
transform 1 0 23328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_244
timestamp 1679585382
transform 1 0 24000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_251
timestamp 1679585382
transform 1 0 24672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_258
timestamp 1679585382
transform 1 0 25344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_265
timestamp 1679585382
transform 1 0 26016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_272
timestamp 1679585382
transform 1 0 26688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_279
timestamp 1679585382
transform 1 0 27360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_286
timestamp 1679585382
transform 1 0 28032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_293
timestamp 1679585382
transform 1 0 28704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_300
timestamp 1679585382
transform 1 0 29376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_307
timestamp 1679585382
transform 1 0 30048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_314
timestamp 1679585382
transform 1 0 30720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_321
timestamp 1679585382
transform 1 0 31392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_328
timestamp 1679585382
transform 1 0 32064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_335
timestamp 1679585382
transform 1 0 32736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_342
timestamp 1679585382
transform 1 0 33408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_349
timestamp 1679585382
transform 1 0 34080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_356
timestamp 1679585382
transform 1 0 34752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_363
timestamp 1679585382
transform 1 0 35424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_370
timestamp 1679585382
transform 1 0 36096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_377
timestamp 1679585382
transform 1 0 36768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_384
timestamp 1679585382
transform 1 0 37440 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_391
timestamp 1679585382
transform 1 0 38112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_398
timestamp 1679585382
transform 1 0 38784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_405
timestamp 1679585382
transform 1 0 39456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_412
timestamp 1679585382
transform 1 0 40128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_419
timestamp 1679585382
transform 1 0 40800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_426
timestamp 1679585382
transform 1 0 41472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_433
timestamp 1679585382
transform 1 0 42144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_440
timestamp 1679585382
transform 1 0 42816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_447
timestamp 1679585382
transform 1 0 43488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_454
timestamp 1679585382
transform 1 0 44160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_461
timestamp 1679585382
transform 1 0 44832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_468
timestamp 1679585382
transform 1 0 45504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_475
timestamp 1679585382
transform 1 0 46176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_482
timestamp 1679585382
transform 1 0 46848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_489
timestamp 1679585382
transform 1 0 47520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_496
timestamp 1679585382
transform 1 0 48192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_503
timestamp 1679585382
transform 1 0 48864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_510
timestamp 1679585382
transform 1 0 49536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_517
timestamp 1679585382
transform 1 0 50208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_524
timestamp 1679585382
transform 1 0 50880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_531
timestamp 1679585382
transform 1 0 51552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_538
timestamp 1679585382
transform 1 0 52224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_545
timestamp 1679585382
transform 1 0 52896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_552
timestamp 1679585382
transform 1 0 53568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_559
timestamp 1679585382
transform 1 0 54240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_566
timestamp 1679585382
transform 1 0 54912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_573
timestamp 1679585382
transform 1 0 55584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_580
timestamp 1679585382
transform 1 0 56256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_587
timestamp 1679585382
transform 1 0 56928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_594
timestamp 1679585382
transform 1 0 57600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_601
timestamp 1679585382
transform 1 0 58272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_608
timestamp 1679585382
transform 1 0 58944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_615
timestamp 1679585382
transform 1 0 59616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_622
timestamp 1679585382
transform 1 0 60288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_629
timestamp 1679585382
transform 1 0 60960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_636
timestamp 1679585382
transform 1 0 61632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_643
timestamp 1679585382
transform 1 0 62304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_650
timestamp 1679585382
transform 1 0 62976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_657
timestamp 1679585382
transform 1 0 63648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_664
timestamp 1679585382
transform 1 0 64320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_671
timestamp 1679585382
transform 1 0 64992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_678
timestamp 1679585382
transform 1 0 65664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_685
timestamp 1679585382
transform 1 0 66336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_692
timestamp 1679585382
transform 1 0 67008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_699
timestamp 1679585382
transform 1 0 67680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_706
timestamp 1679585382
transform 1 0 68352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_713
timestamp 1679585382
transform 1 0 69024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_720
timestamp 1679585382
transform 1 0 69696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_727
timestamp 1679585382
transform 1 0 70368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_734
timestamp 1679585382
transform 1 0 71040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_741
timestamp 1679585382
transform 1 0 71712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_748
timestamp 1679585382
transform 1 0 72384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_755
timestamp 1679585382
transform 1 0 73056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_762
timestamp 1679585382
transform 1 0 73728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_769
timestamp 1679585382
transform 1 0 74400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_776
timestamp 1679585382
transform 1 0 75072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_783
timestamp 1679585382
transform 1 0 75744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_790
timestamp 1679585382
transform 1 0 76416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_797
timestamp 1679585382
transform 1 0 77088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_804
timestamp 1679585382
transform 1 0 77760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_811
timestamp 1679585382
transform 1 0 78432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_818
timestamp 1679585382
transform 1 0 79104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_825
timestamp 1679585382
transform 1 0 79776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_832
timestamp 1679585382
transform 1 0 80448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_839
timestamp 1679585382
transform 1 0 81120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_846
timestamp 1679585382
transform 1 0 81792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_853
timestamp 1679585382
transform 1 0 82464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_860
timestamp 1679585382
transform 1 0 83136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_867
timestamp 1679585382
transform 1 0 83808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_874
timestamp 1679585382
transform 1 0 84480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_881
timestamp 1679585382
transform 1 0 85152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_888
timestamp 1679585382
transform 1 0 85824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_895
timestamp 1679585382
transform 1 0 86496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_902
timestamp 1679585382
transform 1 0 87168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_909
timestamp 1679585382
transform 1 0 87840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_916
timestamp 1679585382
transform 1 0 88512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_923
timestamp 1679585382
transform 1 0 89184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_930
timestamp 1679585382
transform 1 0 89856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_937
timestamp 1679585382
transform 1 0 90528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_944
timestamp 1679585382
transform 1 0 91200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_951
timestamp 1679585382
transform 1 0 91872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_958
timestamp 1679585382
transform 1 0 92544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_965
timestamp 1679585382
transform 1 0 93216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_972
timestamp 1679585382
transform 1 0 93888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_979
timestamp 1679585382
transform 1 0 94560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_986
timestamp 1679585382
transform 1 0 95232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_993
timestamp 1679585382
transform 1 0 95904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1000
timestamp 1679585382
transform 1 0 96576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1007
timestamp 1679585382
transform 1 0 97248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1014
timestamp 1679585382
transform 1 0 97920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1021
timestamp 1679585382
transform 1 0 98592 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_1028
timestamp 1677583258
transform 1 0 99264 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679585382
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_11
timestamp 1679581501
transform 1 0 1632 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_15
timestamp 1677583704
transform 1 0 2016 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_43
timestamp 1679585382
transform 1 0 4704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_50
timestamp 1679585382
transform 1 0 5376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_57
timestamp 1679585382
transform 1 0 6048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_64
timestamp 1679585382
transform 1 0 6720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_71
timestamp 1679585382
transform 1 0 7392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_78
timestamp 1679581501
transform 1 0 8064 0 1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_14_90
timestamp 1679581501
transform 1 0 9216 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_108
timestamp 1679585382
transform 1 0 10944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_115
timestamp 1679581501
transform 1 0 11616 0 1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_14_128
timestamp 1679581501
transform 1 0 12864 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_132
timestamp 1677583258
transform 1 0 13248 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_142
timestamp 1679585382
transform 1 0 14208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_149
timestamp 1679585382
transform 1 0 14880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_156
timestamp 1679585382
transform 1 0 15552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_163
timestamp 1679585382
transform 1 0 16224 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_170
timestamp 1679585382
transform 1 0 16896 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_177
timestamp 1679585382
transform 1 0 17568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_184
timestamp 1679585382
transform 1 0 18240 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_191
timestamp 1679585382
transform 1 0 18912 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_198
timestamp 1679585382
transform 1 0 19584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_205
timestamp 1679585382
transform 1 0 20256 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_212
timestamp 1679585382
transform 1 0 20928 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_219
timestamp 1679585382
transform 1 0 21600 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_226
timestamp 1679585382
transform 1 0 22272 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_233
timestamp 1679585382
transform 1 0 22944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_240
timestamp 1679585382
transform 1 0 23616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_247
timestamp 1679585382
transform 1 0 24288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_254
timestamp 1679585382
transform 1 0 24960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_261
timestamp 1679585382
transform 1 0 25632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_268
timestamp 1679585382
transform 1 0 26304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_275
timestamp 1679585382
transform 1 0 26976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_282
timestamp 1679585382
transform 1 0 27648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_289
timestamp 1679585382
transform 1 0 28320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_296
timestamp 1679585382
transform 1 0 28992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_303
timestamp 1679585382
transform 1 0 29664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_310
timestamp 1679585382
transform 1 0 30336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_317
timestamp 1679585382
transform 1 0 31008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_324
timestamp 1679585382
transform 1 0 31680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_331
timestamp 1679585382
transform 1 0 32352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_338
timestamp 1679585382
transform 1 0 33024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_345
timestamp 1679585382
transform 1 0 33696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_352
timestamp 1679585382
transform 1 0 34368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_359
timestamp 1679585382
transform 1 0 35040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_366
timestamp 1679585382
transform 1 0 35712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_373
timestamp 1679585382
transform 1 0 36384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_380
timestamp 1679585382
transform 1 0 37056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_387
timestamp 1679585382
transform 1 0 37728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_394
timestamp 1679585382
transform 1 0 38400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_401
timestamp 1679585382
transform 1 0 39072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_408
timestamp 1679585382
transform 1 0 39744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_415
timestamp 1679585382
transform 1 0 40416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_422
timestamp 1679585382
transform 1 0 41088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_429
timestamp 1679585382
transform 1 0 41760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_436
timestamp 1679585382
transform 1 0 42432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_443
timestamp 1679585382
transform 1 0 43104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_450
timestamp 1679585382
transform 1 0 43776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_457
timestamp 1679585382
transform 1 0 44448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_464
timestamp 1679585382
transform 1 0 45120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_471
timestamp 1679585382
transform 1 0 45792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_478
timestamp 1679585382
transform 1 0 46464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_485
timestamp 1679585382
transform 1 0 47136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_492
timestamp 1679585382
transform 1 0 47808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_499
timestamp 1679585382
transform 1 0 48480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_506
timestamp 1679585382
transform 1 0 49152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_513
timestamp 1679585382
transform 1 0 49824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_520
timestamp 1679585382
transform 1 0 50496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_527
timestamp 1679585382
transform 1 0 51168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_534
timestamp 1679585382
transform 1 0 51840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_541
timestamp 1679585382
transform 1 0 52512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_548
timestamp 1679585382
transform 1 0 53184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_555
timestamp 1679585382
transform 1 0 53856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_562
timestamp 1679585382
transform 1 0 54528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_569
timestamp 1679585382
transform 1 0 55200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_576
timestamp 1679585382
transform 1 0 55872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_583
timestamp 1679585382
transform 1 0 56544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_590
timestamp 1679585382
transform 1 0 57216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_597
timestamp 1679585382
transform 1 0 57888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_604
timestamp 1679585382
transform 1 0 58560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_611
timestamp 1679585382
transform 1 0 59232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_618
timestamp 1679585382
transform 1 0 59904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_625
timestamp 1679585382
transform 1 0 60576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_632
timestamp 1679585382
transform 1 0 61248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_639
timestamp 1679585382
transform 1 0 61920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_646
timestamp 1679585382
transform 1 0 62592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_653
timestamp 1679585382
transform 1 0 63264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_660
timestamp 1679585382
transform 1 0 63936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_667
timestamp 1679585382
transform 1 0 64608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_674
timestamp 1679585382
transform 1 0 65280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_681
timestamp 1679585382
transform 1 0 65952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_688
timestamp 1679585382
transform 1 0 66624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_695
timestamp 1679585382
transform 1 0 67296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_702
timestamp 1679585382
transform 1 0 67968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_709
timestamp 1679585382
transform 1 0 68640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_716
timestamp 1679585382
transform 1 0 69312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_723
timestamp 1679585382
transform 1 0 69984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_730
timestamp 1679585382
transform 1 0 70656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_737
timestamp 1679585382
transform 1 0 71328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_744
timestamp 1679585382
transform 1 0 72000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_751
timestamp 1679585382
transform 1 0 72672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_758
timestamp 1679585382
transform 1 0 73344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_765
timestamp 1679585382
transform 1 0 74016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_772
timestamp 1679585382
transform 1 0 74688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_779
timestamp 1679585382
transform 1 0 75360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_786
timestamp 1679585382
transform 1 0 76032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_793
timestamp 1679585382
transform 1 0 76704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_800
timestamp 1679585382
transform 1 0 77376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_807
timestamp 1679585382
transform 1 0 78048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_814
timestamp 1679585382
transform 1 0 78720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_821
timestamp 1679585382
transform 1 0 79392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_828
timestamp 1679585382
transform 1 0 80064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_835
timestamp 1679585382
transform 1 0 80736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_842
timestamp 1679585382
transform 1 0 81408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_849
timestamp 1679585382
transform 1 0 82080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_856
timestamp 1679585382
transform 1 0 82752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_863
timestamp 1679585382
transform 1 0 83424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_870
timestamp 1679585382
transform 1 0 84096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_877
timestamp 1679585382
transform 1 0 84768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_884
timestamp 1679585382
transform 1 0 85440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_891
timestamp 1679585382
transform 1 0 86112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_898
timestamp 1679585382
transform 1 0 86784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_905
timestamp 1679585382
transform 1 0 87456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_912
timestamp 1679585382
transform 1 0 88128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_919
timestamp 1679585382
transform 1 0 88800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_926
timestamp 1679585382
transform 1 0 89472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_933
timestamp 1679585382
transform 1 0 90144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_940
timestamp 1679585382
transform 1 0 90816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_947
timestamp 1679585382
transform 1 0 91488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_954
timestamp 1679585382
transform 1 0 92160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_961
timestamp 1679585382
transform 1 0 92832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_968
timestamp 1679585382
transform 1 0 93504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_975
timestamp 1679585382
transform 1 0 94176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_982
timestamp 1679585382
transform 1 0 94848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_989
timestamp 1679585382
transform 1 0 95520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_996
timestamp 1679585382
transform 1 0 96192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1003
timestamp 1679585382
transform 1 0 96864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1010
timestamp 1679585382
transform 1 0 97536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1017
timestamp 1679585382
transform 1 0 98208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_1024
timestamp 1679581501
transform 1 0 98880 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_1028
timestamp 1677583258
transform 1 0 99264 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679585382
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679585382
transform 1 0 1632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679585382
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_25
timestamp 1679585382
transform 1 0 2976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_32
timestamp 1679585382
transform 1 0 3648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_39
timestamp 1679585382
transform 1 0 4320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_46
timestamp 1679585382
transform 1 0 4992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_53
timestamp 1679585382
transform 1 0 5664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_60
timestamp 1679585382
transform 1 0 6336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_67
timestamp 1679585382
transform 1 0 7008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_74
timestamp 1679585382
transform 1 0 7680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_81
timestamp 1679585382
transform 1 0 8352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_88
timestamp 1679585382
transform 1 0 9024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_120
timestamp 1679585382
transform 1 0 12096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_127
timestamp 1679585382
transform 1 0 12768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_134
timestamp 1679585382
transform 1 0 13440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_141
timestamp 1679585382
transform 1 0 14112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_148
timestamp 1679585382
transform 1 0 14784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_155
timestamp 1679585382
transform 1 0 15456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_162
timestamp 1679585382
transform 1 0 16128 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_169
timestamp 1679585382
transform 1 0 16800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_176
timestamp 1679585382
transform 1 0 17472 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_183
timestamp 1679585382
transform 1 0 18144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_190
timestamp 1679585382
transform 1 0 18816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_197
timestamp 1679585382
transform 1 0 19488 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_204
timestamp 1679585382
transform 1 0 20160 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_211
timestamp 1679585382
transform 1 0 20832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_218
timestamp 1679585382
transform 1 0 21504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_225
timestamp 1679585382
transform 1 0 22176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_232
timestamp 1679585382
transform 1 0 22848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_239
timestamp 1679585382
transform 1 0 23520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_246
timestamp 1679585382
transform 1 0 24192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_253
timestamp 1679585382
transform 1 0 24864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_260
timestamp 1679585382
transform 1 0 25536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_267
timestamp 1679585382
transform 1 0 26208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_274
timestamp 1679585382
transform 1 0 26880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_281
timestamp 1679585382
transform 1 0 27552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_288
timestamp 1679585382
transform 1 0 28224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_295
timestamp 1679585382
transform 1 0 28896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_302
timestamp 1679585382
transform 1 0 29568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_309
timestamp 1679585382
transform 1 0 30240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_316
timestamp 1679585382
transform 1 0 30912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_323
timestamp 1679585382
transform 1 0 31584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_330
timestamp 1679585382
transform 1 0 32256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_337
timestamp 1679585382
transform 1 0 32928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_344
timestamp 1679585382
transform 1 0 33600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_351
timestamp 1679585382
transform 1 0 34272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_358
timestamp 1679585382
transform 1 0 34944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_365
timestamp 1679585382
transform 1 0 35616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_372
timestamp 1679585382
transform 1 0 36288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_379
timestamp 1679585382
transform 1 0 36960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_386
timestamp 1679585382
transform 1 0 37632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_393
timestamp 1679585382
transform 1 0 38304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_400
timestamp 1679585382
transform 1 0 38976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_407
timestamp 1679585382
transform 1 0 39648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_414
timestamp 1679585382
transform 1 0 40320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_421
timestamp 1679585382
transform 1 0 40992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_428
timestamp 1679585382
transform 1 0 41664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_435
timestamp 1679585382
transform 1 0 42336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_442
timestamp 1679585382
transform 1 0 43008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_449
timestamp 1679585382
transform 1 0 43680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_456
timestamp 1679585382
transform 1 0 44352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_463
timestamp 1679585382
transform 1 0 45024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_470
timestamp 1679585382
transform 1 0 45696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_477
timestamp 1679585382
transform 1 0 46368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_484
timestamp 1679585382
transform 1 0 47040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_491
timestamp 1679585382
transform 1 0 47712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_498
timestamp 1679585382
transform 1 0 48384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_505
timestamp 1679585382
transform 1 0 49056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_512
timestamp 1679585382
transform 1 0 49728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_519
timestamp 1679585382
transform 1 0 50400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_526
timestamp 1679585382
transform 1 0 51072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_533
timestamp 1679585382
transform 1 0 51744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_540
timestamp 1679585382
transform 1 0 52416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_547
timestamp 1679585382
transform 1 0 53088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_554
timestamp 1679585382
transform 1 0 53760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_561
timestamp 1679585382
transform 1 0 54432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_568
timestamp 1679585382
transform 1 0 55104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_575
timestamp 1679585382
transform 1 0 55776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_582
timestamp 1679585382
transform 1 0 56448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_589
timestamp 1679585382
transform 1 0 57120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_596
timestamp 1679585382
transform 1 0 57792 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_603
timestamp 1679585382
transform 1 0 58464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_610
timestamp 1679585382
transform 1 0 59136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_617
timestamp 1679585382
transform 1 0 59808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_624
timestamp 1679585382
transform 1 0 60480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_631
timestamp 1679585382
transform 1 0 61152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_638
timestamp 1679585382
transform 1 0 61824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_645
timestamp 1679585382
transform 1 0 62496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_652
timestamp 1679585382
transform 1 0 63168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_659
timestamp 1679585382
transform 1 0 63840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_666
timestamp 1679585382
transform 1 0 64512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_673
timestamp 1679585382
transform 1 0 65184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_680
timestamp 1679585382
transform 1 0 65856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_687
timestamp 1679585382
transform 1 0 66528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_694
timestamp 1679585382
transform 1 0 67200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_701
timestamp 1679585382
transform 1 0 67872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_708
timestamp 1679585382
transform 1 0 68544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_715
timestamp 1679585382
transform 1 0 69216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_722
timestamp 1679585382
transform 1 0 69888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_729
timestamp 1679585382
transform 1 0 70560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_736
timestamp 1679585382
transform 1 0 71232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_743
timestamp 1679585382
transform 1 0 71904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_750
timestamp 1679585382
transform 1 0 72576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_757
timestamp 1679585382
transform 1 0 73248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_764
timestamp 1679585382
transform 1 0 73920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_771
timestamp 1679585382
transform 1 0 74592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_778
timestamp 1679585382
transform 1 0 75264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_785
timestamp 1679585382
transform 1 0 75936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_792
timestamp 1679585382
transform 1 0 76608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_799
timestamp 1679585382
transform 1 0 77280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_806
timestamp 1679585382
transform 1 0 77952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_813
timestamp 1679585382
transform 1 0 78624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_820
timestamp 1679585382
transform 1 0 79296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_827
timestamp 1679585382
transform 1 0 79968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_834
timestamp 1679585382
transform 1 0 80640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_841
timestamp 1679585382
transform 1 0 81312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_848
timestamp 1679585382
transform 1 0 81984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_855
timestamp 1679585382
transform 1 0 82656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_862
timestamp 1679585382
transform 1 0 83328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_869
timestamp 1679585382
transform 1 0 84000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_876
timestamp 1679585382
transform 1 0 84672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_883
timestamp 1679585382
transform 1 0 85344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_890
timestamp 1679585382
transform 1 0 86016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_897
timestamp 1679585382
transform 1 0 86688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_904
timestamp 1679585382
transform 1 0 87360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_911
timestamp 1679585382
transform 1 0 88032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_918
timestamp 1679585382
transform 1 0 88704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_925
timestamp 1679585382
transform 1 0 89376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_932
timestamp 1679585382
transform 1 0 90048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_939
timestamp 1679585382
transform 1 0 90720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_946
timestamp 1679585382
transform 1 0 91392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_953
timestamp 1679585382
transform 1 0 92064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_960
timestamp 1679585382
transform 1 0 92736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_967
timestamp 1679585382
transform 1 0 93408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_974
timestamp 1679585382
transform 1 0 94080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_981
timestamp 1679585382
transform 1 0 94752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_988
timestamp 1679585382
transform 1 0 95424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_995
timestamp 1679585382
transform 1 0 96096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1002
timestamp 1679585382
transform 1 0 96768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1009
timestamp 1679585382
transform 1 0 97440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1016
timestamp 1679585382
transform 1 0 98112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_1023
timestamp 1679581501
transform 1 0 98784 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_1027
timestamp 1677583704
transform 1 0 99168 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679585382
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_11
timestamp 1679585382
transform 1 0 1632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_18
timestamp 1679581501
transform 1 0 2304 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_22
timestamp 1677583704
transform 1 0 2688 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_37
timestamp 1679585382
transform 1 0 4128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_44
timestamp 1679585382
transform 1 0 4800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_51
timestamp 1679585382
transform 1 0 5472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_58
timestamp 1679585382
transform 1 0 6144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_65
timestamp 1679585382
transform 1 0 6816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_72
timestamp 1679585382
transform 1 0 7488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_79
timestamp 1679585382
transform 1 0 8160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_86
timestamp 1679585382
transform 1 0 8832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_93
timestamp 1679581501
transform 1 0 9504 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_97
timestamp 1677583704
transform 1 0 9888 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_104
timestamp 1679585382
transform 1 0 10560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_111
timestamp 1679585382
transform 1 0 11232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_118
timestamp 1679585382
transform 1 0 11904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_125
timestamp 1679585382
transform 1 0 12576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_132
timestamp 1679585382
transform 1 0 13248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_139
timestamp 1679585382
transform 1 0 13920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_146
timestamp 1679585382
transform 1 0 14592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_153
timestamp 1679585382
transform 1 0 15264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_160
timestamp 1679585382
transform 1 0 15936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_167
timestamp 1679585382
transform 1 0 16608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_174
timestamp 1679585382
transform 1 0 17280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_181
timestamp 1679585382
transform 1 0 17952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_188
timestamp 1679585382
transform 1 0 18624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_195
timestamp 1679585382
transform 1 0 19296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_202
timestamp 1679585382
transform 1 0 19968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_209
timestamp 1679585382
transform 1 0 20640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_216
timestamp 1679585382
transform 1 0 21312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_223
timestamp 1679585382
transform 1 0 21984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_230
timestamp 1679585382
transform 1 0 22656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_237
timestamp 1679585382
transform 1 0 23328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_244
timestamp 1679585382
transform 1 0 24000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_251
timestamp 1679585382
transform 1 0 24672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_258
timestamp 1679585382
transform 1 0 25344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_265
timestamp 1679585382
transform 1 0 26016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_272
timestamp 1679585382
transform 1 0 26688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_279
timestamp 1679585382
transform 1 0 27360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_286
timestamp 1679585382
transform 1 0 28032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_293
timestamp 1679585382
transform 1 0 28704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_300
timestamp 1679585382
transform 1 0 29376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_307
timestamp 1679585382
transform 1 0 30048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_314
timestamp 1679585382
transform 1 0 30720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_321
timestamp 1679585382
transform 1 0 31392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_328
timestamp 1679585382
transform 1 0 32064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_335
timestamp 1679585382
transform 1 0 32736 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_342
timestamp 1679585382
transform 1 0 33408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_349
timestamp 1679585382
transform 1 0 34080 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_356
timestamp 1679585382
transform 1 0 34752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_363
timestamp 1679585382
transform 1 0 35424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_370
timestamp 1679585382
transform 1 0 36096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_377
timestamp 1679585382
transform 1 0 36768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_384
timestamp 1679585382
transform 1 0 37440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_391
timestamp 1679585382
transform 1 0 38112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_398
timestamp 1679585382
transform 1 0 38784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_405
timestamp 1679585382
transform 1 0 39456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_412
timestamp 1679585382
transform 1 0 40128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_419
timestamp 1679585382
transform 1 0 40800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_426
timestamp 1679585382
transform 1 0 41472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_433
timestamp 1679585382
transform 1 0 42144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_440
timestamp 1679585382
transform 1 0 42816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_447
timestamp 1679585382
transform 1 0 43488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_454
timestamp 1679585382
transform 1 0 44160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_461
timestamp 1679585382
transform 1 0 44832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_468
timestamp 1679585382
transform 1 0 45504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_475
timestamp 1679585382
transform 1 0 46176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_482
timestamp 1679585382
transform 1 0 46848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_489
timestamp 1679585382
transform 1 0 47520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_496
timestamp 1679585382
transform 1 0 48192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_503
timestamp 1679585382
transform 1 0 48864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_510
timestamp 1679585382
transform 1 0 49536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_517
timestamp 1679585382
transform 1 0 50208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_524
timestamp 1679585382
transform 1 0 50880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_531
timestamp 1679585382
transform 1 0 51552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_538
timestamp 1679585382
transform 1 0 52224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_545
timestamp 1679585382
transform 1 0 52896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_552
timestamp 1679585382
transform 1 0 53568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_559
timestamp 1679585382
transform 1 0 54240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_566
timestamp 1679585382
transform 1 0 54912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_573
timestamp 1679585382
transform 1 0 55584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_580
timestamp 1679585382
transform 1 0 56256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_587
timestamp 1679585382
transform 1 0 56928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_594
timestamp 1679585382
transform 1 0 57600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_601
timestamp 1679585382
transform 1 0 58272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_608
timestamp 1679585382
transform 1 0 58944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_615
timestamp 1679585382
transform 1 0 59616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_622
timestamp 1679585382
transform 1 0 60288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_629
timestamp 1679585382
transform 1 0 60960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_636
timestamp 1679585382
transform 1 0 61632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_643
timestamp 1679585382
transform 1 0 62304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_650
timestamp 1679585382
transform 1 0 62976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_657
timestamp 1679585382
transform 1 0 63648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_664
timestamp 1679585382
transform 1 0 64320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_671
timestamp 1679585382
transform 1 0 64992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_678
timestamp 1679585382
transform 1 0 65664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_685
timestamp 1679585382
transform 1 0 66336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_692
timestamp 1679585382
transform 1 0 67008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_699
timestamp 1679585382
transform 1 0 67680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_706
timestamp 1679585382
transform 1 0 68352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_713
timestamp 1679585382
transform 1 0 69024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_720
timestamp 1679585382
transform 1 0 69696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_727
timestamp 1679585382
transform 1 0 70368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_734
timestamp 1679585382
transform 1 0 71040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_741
timestamp 1679585382
transform 1 0 71712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_748
timestamp 1679585382
transform 1 0 72384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_755
timestamp 1679585382
transform 1 0 73056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_762
timestamp 1679585382
transform 1 0 73728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_769
timestamp 1679585382
transform 1 0 74400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_776
timestamp 1679585382
transform 1 0 75072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_783
timestamp 1679585382
transform 1 0 75744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_790
timestamp 1679585382
transform 1 0 76416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_797
timestamp 1679585382
transform 1 0 77088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_804
timestamp 1679585382
transform 1 0 77760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_811
timestamp 1679585382
transform 1 0 78432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_818
timestamp 1679585382
transform 1 0 79104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_825
timestamp 1679585382
transform 1 0 79776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_832
timestamp 1679585382
transform 1 0 80448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_839
timestamp 1679585382
transform 1 0 81120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_846
timestamp 1679585382
transform 1 0 81792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_853
timestamp 1679585382
transform 1 0 82464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_860
timestamp 1679585382
transform 1 0 83136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_867
timestamp 1679585382
transform 1 0 83808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_874
timestamp 1679585382
transform 1 0 84480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_881
timestamp 1679585382
transform 1 0 85152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_888
timestamp 1679585382
transform 1 0 85824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_895
timestamp 1679585382
transform 1 0 86496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_902
timestamp 1679585382
transform 1 0 87168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_909
timestamp 1679585382
transform 1 0 87840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_916
timestamp 1679585382
transform 1 0 88512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_923
timestamp 1679585382
transform 1 0 89184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_930
timestamp 1679585382
transform 1 0 89856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_937
timestamp 1679585382
transform 1 0 90528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_944
timestamp 1679585382
transform 1 0 91200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_951
timestamp 1679585382
transform 1 0 91872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_958
timestamp 1679585382
transform 1 0 92544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_965
timestamp 1679585382
transform 1 0 93216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_972
timestamp 1679585382
transform 1 0 93888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_979
timestamp 1679585382
transform 1 0 94560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_986
timestamp 1679585382
transform 1 0 95232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_993
timestamp 1679585382
transform 1 0 95904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1000
timestamp 1679585382
transform 1 0 96576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1007
timestamp 1679585382
transform 1 0 97248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1014
timestamp 1679585382
transform 1 0 97920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1021
timestamp 1679585382
transform 1 0 98592 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_1028
timestamp 1677583258
transform 1 0 99264 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679585382
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679585382
transform 1 0 1248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_14
timestamp 1679585382
transform 1 0 1920 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_21
timestamp 1677583258
transform 1 0 2592 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_49
timestamp 1679585382
transform 1 0 5280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_56
timestamp 1679585382
transform 1 0 5952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_63
timestamp 1679585382
transform 1 0 6624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_70
timestamp 1679585382
transform 1 0 7296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_77
timestamp 1679585382
transform 1 0 7968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_84
timestamp 1679585382
transform 1 0 8640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_91
timestamp 1679585382
transform 1 0 9312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_98
timestamp 1679585382
transform 1 0 9984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_105
timestamp 1679581501
transform 1 0 10656 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_114
timestamp 1679585382
transform 1 0 11520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_121
timestamp 1679585382
transform 1 0 12192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_128
timestamp 1679581501
transform 1 0 12864 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_132
timestamp 1677583704
transform 1 0 13248 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_143
timestamp 1679585382
transform 1 0 14304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_150
timestamp 1679585382
transform 1 0 14976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_157
timestamp 1679585382
transform 1 0 15648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_164
timestamp 1679585382
transform 1 0 16320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_171
timestamp 1679585382
transform 1 0 16992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_178
timestamp 1679585382
transform 1 0 17664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_185
timestamp 1679585382
transform 1 0 18336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_192
timestamp 1679585382
transform 1 0 19008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_199
timestamp 1679585382
transform 1 0 19680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_206
timestamp 1679585382
transform 1 0 20352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_213
timestamp 1679585382
transform 1 0 21024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_220
timestamp 1679585382
transform 1 0 21696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_227
timestamp 1679585382
transform 1 0 22368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_234
timestamp 1679585382
transform 1 0 23040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_241
timestamp 1679585382
transform 1 0 23712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_248
timestamp 1679585382
transform 1 0 24384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_255
timestamp 1679585382
transform 1 0 25056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_262
timestamp 1679585382
transform 1 0 25728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_269
timestamp 1679585382
transform 1 0 26400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_276
timestamp 1679585382
transform 1 0 27072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_283
timestamp 1679585382
transform 1 0 27744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_290
timestamp 1679585382
transform 1 0 28416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_297
timestamp 1679585382
transform 1 0 29088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_304
timestamp 1679585382
transform 1 0 29760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_311
timestamp 1679585382
transform 1 0 30432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_318
timestamp 1679585382
transform 1 0 31104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_325
timestamp 1679585382
transform 1 0 31776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_332
timestamp 1679585382
transform 1 0 32448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_339
timestamp 1679585382
transform 1 0 33120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_346
timestamp 1679585382
transform 1 0 33792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_353
timestamp 1679585382
transform 1 0 34464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_360
timestamp 1679585382
transform 1 0 35136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_367
timestamp 1679585382
transform 1 0 35808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_374
timestamp 1679585382
transform 1 0 36480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_381
timestamp 1679585382
transform 1 0 37152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_388
timestamp 1679585382
transform 1 0 37824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_395
timestamp 1679585382
transform 1 0 38496 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_402
timestamp 1679585382
transform 1 0 39168 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_409
timestamp 1679585382
transform 1 0 39840 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_416
timestamp 1679585382
transform 1 0 40512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_423
timestamp 1679585382
transform 1 0 41184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_430
timestamp 1679585382
transform 1 0 41856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_437
timestamp 1679585382
transform 1 0 42528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_444
timestamp 1679585382
transform 1 0 43200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_451
timestamp 1679585382
transform 1 0 43872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_458
timestamp 1679585382
transform 1 0 44544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_465
timestamp 1679585382
transform 1 0 45216 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_472
timestamp 1679585382
transform 1 0 45888 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_479
timestamp 1679585382
transform 1 0 46560 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_486
timestamp 1679585382
transform 1 0 47232 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_493
timestamp 1679585382
transform 1 0 47904 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_500
timestamp 1679585382
transform 1 0 48576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_507
timestamp 1679585382
transform 1 0 49248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_514
timestamp 1679585382
transform 1 0 49920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_521
timestamp 1679585382
transform 1 0 50592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_528
timestamp 1679585382
transform 1 0 51264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_535
timestamp 1679585382
transform 1 0 51936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_542
timestamp 1679585382
transform 1 0 52608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_549
timestamp 1679585382
transform 1 0 53280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_556
timestamp 1679585382
transform 1 0 53952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_563
timestamp 1679585382
transform 1 0 54624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_570
timestamp 1679585382
transform 1 0 55296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_577
timestamp 1679585382
transform 1 0 55968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_584
timestamp 1679585382
transform 1 0 56640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_591
timestamp 1679585382
transform 1 0 57312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_598
timestamp 1679585382
transform 1 0 57984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_605
timestamp 1679585382
transform 1 0 58656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_612
timestamp 1679585382
transform 1 0 59328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_619
timestamp 1679585382
transform 1 0 60000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_626
timestamp 1679585382
transform 1 0 60672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_633
timestamp 1679585382
transform 1 0 61344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_640
timestamp 1679585382
transform 1 0 62016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_647
timestamp 1679585382
transform 1 0 62688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_654
timestamp 1679585382
transform 1 0 63360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_661
timestamp 1679585382
transform 1 0 64032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_668
timestamp 1679585382
transform 1 0 64704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_675
timestamp 1679585382
transform 1 0 65376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_682
timestamp 1679585382
transform 1 0 66048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_689
timestamp 1679585382
transform 1 0 66720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_696
timestamp 1679585382
transform 1 0 67392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_703
timestamp 1679585382
transform 1 0 68064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_710
timestamp 1679585382
transform 1 0 68736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_717
timestamp 1679585382
transform 1 0 69408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_724
timestamp 1679585382
transform 1 0 70080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_731
timestamp 1679585382
transform 1 0 70752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_738
timestamp 1679585382
transform 1 0 71424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_745
timestamp 1679585382
transform 1 0 72096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_752
timestamp 1679585382
transform 1 0 72768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_759
timestamp 1679585382
transform 1 0 73440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_766
timestamp 1679585382
transform 1 0 74112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_773
timestamp 1679585382
transform 1 0 74784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_780
timestamp 1679585382
transform 1 0 75456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_787
timestamp 1679585382
transform 1 0 76128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_794
timestamp 1679585382
transform 1 0 76800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_801
timestamp 1679585382
transform 1 0 77472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_808
timestamp 1679585382
transform 1 0 78144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_815
timestamp 1679585382
transform 1 0 78816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_822
timestamp 1679585382
transform 1 0 79488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_829
timestamp 1679585382
transform 1 0 80160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_836
timestamp 1679585382
transform 1 0 80832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_843
timestamp 1679585382
transform 1 0 81504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_850
timestamp 1679585382
transform 1 0 82176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_857
timestamp 1679585382
transform 1 0 82848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_864
timestamp 1679585382
transform 1 0 83520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_871
timestamp 1679585382
transform 1 0 84192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_878
timestamp 1679585382
transform 1 0 84864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_885
timestamp 1679585382
transform 1 0 85536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_892
timestamp 1679585382
transform 1 0 86208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_899
timestamp 1679585382
transform 1 0 86880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_906
timestamp 1679585382
transform 1 0 87552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_913
timestamp 1679585382
transform 1 0 88224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_920
timestamp 1679585382
transform 1 0 88896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_927
timestamp 1679585382
transform 1 0 89568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_934
timestamp 1679585382
transform 1 0 90240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_941
timestamp 1679585382
transform 1 0 90912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_948
timestamp 1679585382
transform 1 0 91584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_955
timestamp 1679585382
transform 1 0 92256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_962
timestamp 1679585382
transform 1 0 92928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_969
timestamp 1679585382
transform 1 0 93600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_976
timestamp 1679585382
transform 1 0 94272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_983
timestamp 1679585382
transform 1 0 94944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_990
timestamp 1679585382
transform 1 0 95616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_997
timestamp 1679585382
transform 1 0 96288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1004
timestamp 1679585382
transform 1 0 96960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1011
timestamp 1679585382
transform 1 0 97632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1018
timestamp 1679585382
transform 1 0 98304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_1025
timestamp 1679581501
transform 1 0 98976 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_4
timestamp 1679585382
transform 1 0 960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_11
timestamp 1679585382
transform 1 0 1632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_18
timestamp 1679585382
transform 1 0 2304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_25
timestamp 1679585382
transform 1 0 2976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_32
timestamp 1679585382
transform 1 0 3648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_39
timestamp 1679585382
transform 1 0 4320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_46
timestamp 1679585382
transform 1 0 4992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_53
timestamp 1679585382
transform 1 0 5664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_60
timestamp 1679585382
transform 1 0 6336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_67
timestamp 1679585382
transform 1 0 7008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_74
timestamp 1679585382
transform 1 0 7680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_81
timestamp 1679585382
transform 1 0 8352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_88
timestamp 1679585382
transform 1 0 9024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_95
timestamp 1679585382
transform 1 0 9696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_102
timestamp 1679585382
transform 1 0 10368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_109
timestamp 1679585382
transform 1 0 11040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_116
timestamp 1679585382
transform 1 0 11712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_123
timestamp 1679585382
transform 1 0 12384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_157
timestamp 1679585382
transform 1 0 15648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_164
timestamp 1679585382
transform 1 0 16320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_171
timestamp 1679585382
transform 1 0 16992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_178
timestamp 1679585382
transform 1 0 17664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_185
timestamp 1679585382
transform 1 0 18336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_192
timestamp 1679585382
transform 1 0 19008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_199
timestamp 1679585382
transform 1 0 19680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_206
timestamp 1679585382
transform 1 0 20352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_213
timestamp 1679585382
transform 1 0 21024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_220
timestamp 1679585382
transform 1 0 21696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_227
timestamp 1679585382
transform 1 0 22368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_234
timestamp 1679585382
transform 1 0 23040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_241
timestamp 1679585382
transform 1 0 23712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_248
timestamp 1679585382
transform 1 0 24384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_255
timestamp 1679585382
transform 1 0 25056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_262
timestamp 1679585382
transform 1 0 25728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_269
timestamp 1679585382
transform 1 0 26400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_276
timestamp 1679585382
transform 1 0 27072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_283
timestamp 1679585382
transform 1 0 27744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_290
timestamp 1679585382
transform 1 0 28416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_297
timestamp 1679585382
transform 1 0 29088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_304
timestamp 1679585382
transform 1 0 29760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_311
timestamp 1679585382
transform 1 0 30432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_318
timestamp 1679585382
transform 1 0 31104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_325
timestamp 1679585382
transform 1 0 31776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_332
timestamp 1679585382
transform 1 0 32448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_339
timestamp 1679585382
transform 1 0 33120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_346
timestamp 1679585382
transform 1 0 33792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_353
timestamp 1679585382
transform 1 0 34464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_360
timestamp 1679585382
transform 1 0 35136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_367
timestamp 1679585382
transform 1 0 35808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_374
timestamp 1679585382
transform 1 0 36480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_381
timestamp 1679585382
transform 1 0 37152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_388
timestamp 1679585382
transform 1 0 37824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_395
timestamp 1679585382
transform 1 0 38496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_402
timestamp 1679585382
transform 1 0 39168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_409
timestamp 1679585382
transform 1 0 39840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_416
timestamp 1679585382
transform 1 0 40512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_423
timestamp 1679585382
transform 1 0 41184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_430
timestamp 1679585382
transform 1 0 41856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_437
timestamp 1679585382
transform 1 0 42528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_444
timestamp 1679585382
transform 1 0 43200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_451
timestamp 1679585382
transform 1 0 43872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_458
timestamp 1679585382
transform 1 0 44544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_465
timestamp 1679585382
transform 1 0 45216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_472
timestamp 1679585382
transform 1 0 45888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_479
timestamp 1679585382
transform 1 0 46560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_486
timestamp 1679585382
transform 1 0 47232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_493
timestamp 1679585382
transform 1 0 47904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_500
timestamp 1679585382
transform 1 0 48576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_507
timestamp 1679585382
transform 1 0 49248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_514
timestamp 1679585382
transform 1 0 49920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_521
timestamp 1679585382
transform 1 0 50592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_528
timestamp 1679585382
transform 1 0 51264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_535
timestamp 1679585382
transform 1 0 51936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_542
timestamp 1679585382
transform 1 0 52608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_549
timestamp 1679585382
transform 1 0 53280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_556
timestamp 1679585382
transform 1 0 53952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_563
timestamp 1679585382
transform 1 0 54624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_570
timestamp 1679585382
transform 1 0 55296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_577
timestamp 1679585382
transform 1 0 55968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_584
timestamp 1679585382
transform 1 0 56640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_591
timestamp 1679585382
transform 1 0 57312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_598
timestamp 1679585382
transform 1 0 57984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_605
timestamp 1679585382
transform 1 0 58656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_612
timestamp 1679585382
transform 1 0 59328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_619
timestamp 1679585382
transform 1 0 60000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_626
timestamp 1679585382
transform 1 0 60672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_633
timestamp 1679585382
transform 1 0 61344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_640
timestamp 1679585382
transform 1 0 62016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_647
timestamp 1679585382
transform 1 0 62688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_654
timestamp 1679585382
transform 1 0 63360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_661
timestamp 1679585382
transform 1 0 64032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_668
timestamp 1679585382
transform 1 0 64704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_675
timestamp 1679585382
transform 1 0 65376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_682
timestamp 1679585382
transform 1 0 66048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_689
timestamp 1679585382
transform 1 0 66720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_696
timestamp 1679585382
transform 1 0 67392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_703
timestamp 1679585382
transform 1 0 68064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_710
timestamp 1679585382
transform 1 0 68736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_717
timestamp 1679585382
transform 1 0 69408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_724
timestamp 1679585382
transform 1 0 70080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_731
timestamp 1679585382
transform 1 0 70752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_738
timestamp 1679585382
transform 1 0 71424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_745
timestamp 1679585382
transform 1 0 72096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_752
timestamp 1679585382
transform 1 0 72768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_759
timestamp 1679585382
transform 1 0 73440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_766
timestamp 1679585382
transform 1 0 74112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_773
timestamp 1679585382
transform 1 0 74784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_780
timestamp 1679585382
transform 1 0 75456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_787
timestamp 1679585382
transform 1 0 76128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_794
timestamp 1679585382
transform 1 0 76800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_801
timestamp 1679585382
transform 1 0 77472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_808
timestamp 1679585382
transform 1 0 78144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_815
timestamp 1679585382
transform 1 0 78816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_822
timestamp 1679585382
transform 1 0 79488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_829
timestamp 1679585382
transform 1 0 80160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_836
timestamp 1679585382
transform 1 0 80832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_843
timestamp 1679585382
transform 1 0 81504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_850
timestamp 1679585382
transform 1 0 82176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_857
timestamp 1679585382
transform 1 0 82848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_864
timestamp 1679585382
transform 1 0 83520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_871
timestamp 1679585382
transform 1 0 84192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_878
timestamp 1679585382
transform 1 0 84864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_885
timestamp 1679585382
transform 1 0 85536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_892
timestamp 1679585382
transform 1 0 86208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_899
timestamp 1679585382
transform 1 0 86880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_906
timestamp 1679585382
transform 1 0 87552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_913
timestamp 1679585382
transform 1 0 88224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_920
timestamp 1679585382
transform 1 0 88896 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_927
timestamp 1679585382
transform 1 0 89568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_934
timestamp 1679585382
transform 1 0 90240 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_941
timestamp 1679585382
transform 1 0 90912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_948
timestamp 1679585382
transform 1 0 91584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_955
timestamp 1679585382
transform 1 0 92256 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_962
timestamp 1679585382
transform 1 0 92928 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_969
timestamp 1679585382
transform 1 0 93600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_976
timestamp 1679585382
transform 1 0 94272 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_983
timestamp 1679585382
transform 1 0 94944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_990
timestamp 1679585382
transform 1 0 95616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_997
timestamp 1679585382
transform 1 0 96288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1004
timestamp 1679585382
transform 1 0 96960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1011
timestamp 1679585382
transform 1 0 97632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1018
timestamp 1679585382
transform 1 0 98304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_1025
timestamp 1679581501
transform 1 0 98976 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_4
timestamp 1679585382
transform 1 0 960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_11
timestamp 1679585382
transform 1 0 1632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679585382
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_25
timestamp 1679585382
transform 1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_32
timestamp 1679585382
transform 1 0 3648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_39
timestamp 1679585382
transform 1 0 4320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_46
timestamp 1679585382
transform 1 0 4992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_53
timestamp 1679585382
transform 1 0 5664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_60
timestamp 1679585382
transform 1 0 6336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_67
timestamp 1679585382
transform 1 0 7008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_74
timestamp 1679585382
transform 1 0 7680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_81
timestamp 1679581501
transform 1 0 8352 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_85
timestamp 1677583258
transform 1 0 8736 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_111
timestamp 1679585382
transform 1 0 11232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_118
timestamp 1679585382
transform 1 0 11904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_125
timestamp 1679585382
transform 1 0 12576 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_132
timestamp 1677583704
transform 1 0 13248 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_134
timestamp 1677583258
transform 1 0 13440 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_139
timestamp 1679585382
transform 1 0 13920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_146
timestamp 1679585382
transform 1 0 14592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_153
timestamp 1679585382
transform 1 0 15264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_160
timestamp 1679585382
transform 1 0 15936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_167
timestamp 1679585382
transform 1 0 16608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_174
timestamp 1679585382
transform 1 0 17280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_181
timestamp 1679585382
transform 1 0 17952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_188
timestamp 1679585382
transform 1 0 18624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_195
timestamp 1679585382
transform 1 0 19296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_202
timestamp 1679585382
transform 1 0 19968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_209
timestamp 1679585382
transform 1 0 20640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_216
timestamp 1679585382
transform 1 0 21312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_223
timestamp 1679585382
transform 1 0 21984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_230
timestamp 1679585382
transform 1 0 22656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_237
timestamp 1679585382
transform 1 0 23328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_244
timestamp 1679585382
transform 1 0 24000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_251
timestamp 1679585382
transform 1 0 24672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_258
timestamp 1679585382
transform 1 0 25344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_265
timestamp 1679585382
transform 1 0 26016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_272
timestamp 1679585382
transform 1 0 26688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_279
timestamp 1679585382
transform 1 0 27360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_286
timestamp 1679585382
transform 1 0 28032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_293
timestamp 1679585382
transform 1 0 28704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_300
timestamp 1679585382
transform 1 0 29376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_307
timestamp 1679585382
transform 1 0 30048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_314
timestamp 1679585382
transform 1 0 30720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_321
timestamp 1679585382
transform 1 0 31392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_328
timestamp 1679585382
transform 1 0 32064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_335
timestamp 1679585382
transform 1 0 32736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_342
timestamp 1679585382
transform 1 0 33408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_349
timestamp 1679585382
transform 1 0 34080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_356
timestamp 1679585382
transform 1 0 34752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_363
timestamp 1679585382
transform 1 0 35424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_370
timestamp 1679585382
transform 1 0 36096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_377
timestamp 1679585382
transform 1 0 36768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_384
timestamp 1679585382
transform 1 0 37440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_391
timestamp 1679585382
transform 1 0 38112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_398
timestamp 1679585382
transform 1 0 38784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_405
timestamp 1679585382
transform 1 0 39456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_412
timestamp 1679585382
transform 1 0 40128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_419
timestamp 1679585382
transform 1 0 40800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_426
timestamp 1679585382
transform 1 0 41472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_433
timestamp 1679585382
transform 1 0 42144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_440
timestamp 1679585382
transform 1 0 42816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_447
timestamp 1679585382
transform 1 0 43488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_454
timestamp 1679585382
transform 1 0 44160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_461
timestamp 1679585382
transform 1 0 44832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_468
timestamp 1679585382
transform 1 0 45504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_475
timestamp 1679585382
transform 1 0 46176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_482
timestamp 1679585382
transform 1 0 46848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_489
timestamp 1679585382
transform 1 0 47520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_496
timestamp 1679585382
transform 1 0 48192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_503
timestamp 1679585382
transform 1 0 48864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_510
timestamp 1679585382
transform 1 0 49536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_517
timestamp 1679585382
transform 1 0 50208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_524
timestamp 1679585382
transform 1 0 50880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_531
timestamp 1679585382
transform 1 0 51552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_538
timestamp 1679585382
transform 1 0 52224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_545
timestamp 1679585382
transform 1 0 52896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_552
timestamp 1679585382
transform 1 0 53568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_559
timestamp 1679585382
transform 1 0 54240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_566
timestamp 1679585382
transform 1 0 54912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_573
timestamp 1679585382
transform 1 0 55584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_580
timestamp 1679585382
transform 1 0 56256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_587
timestamp 1679585382
transform 1 0 56928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_594
timestamp 1679585382
transform 1 0 57600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_601
timestamp 1679585382
transform 1 0 58272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_608
timestamp 1679585382
transform 1 0 58944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_615
timestamp 1679585382
transform 1 0 59616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_622
timestamp 1679585382
transform 1 0 60288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_629
timestamp 1679585382
transform 1 0 60960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_636
timestamp 1679585382
transform 1 0 61632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_643
timestamp 1679585382
transform 1 0 62304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_650
timestamp 1679585382
transform 1 0 62976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_657
timestamp 1679585382
transform 1 0 63648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_664
timestamp 1679585382
transform 1 0 64320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_671
timestamp 1679585382
transform 1 0 64992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_678
timestamp 1679585382
transform 1 0 65664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_685
timestamp 1679585382
transform 1 0 66336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_692
timestamp 1679585382
transform 1 0 67008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_699
timestamp 1679585382
transform 1 0 67680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_706
timestamp 1679585382
transform 1 0 68352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_713
timestamp 1679585382
transform 1 0 69024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_720
timestamp 1679585382
transform 1 0 69696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_727
timestamp 1679585382
transform 1 0 70368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_734
timestamp 1679585382
transform 1 0 71040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_741
timestamp 1679585382
transform 1 0 71712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_748
timestamp 1679585382
transform 1 0 72384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_755
timestamp 1679585382
transform 1 0 73056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_762
timestamp 1679585382
transform 1 0 73728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_769
timestamp 1679585382
transform 1 0 74400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_776
timestamp 1679585382
transform 1 0 75072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_783
timestamp 1679585382
transform 1 0 75744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_790
timestamp 1679585382
transform 1 0 76416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_797
timestamp 1679585382
transform 1 0 77088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_804
timestamp 1679585382
transform 1 0 77760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_811
timestamp 1679585382
transform 1 0 78432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_818
timestamp 1679585382
transform 1 0 79104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_825
timestamp 1679585382
transform 1 0 79776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_832
timestamp 1679585382
transform 1 0 80448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_839
timestamp 1679585382
transform 1 0 81120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_846
timestamp 1679585382
transform 1 0 81792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_853
timestamp 1679585382
transform 1 0 82464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_860
timestamp 1679585382
transform 1 0 83136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_867
timestamp 1679585382
transform 1 0 83808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_874
timestamp 1679585382
transform 1 0 84480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_881
timestamp 1679585382
transform 1 0 85152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_888
timestamp 1679585382
transform 1 0 85824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_895
timestamp 1679585382
transform 1 0 86496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_902
timestamp 1679585382
transform 1 0 87168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_909
timestamp 1679585382
transform 1 0 87840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_916
timestamp 1679585382
transform 1 0 88512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_923
timestamp 1679585382
transform 1 0 89184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_930
timestamp 1679585382
transform 1 0 89856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_937
timestamp 1679585382
transform 1 0 90528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_944
timestamp 1679585382
transform 1 0 91200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_951
timestamp 1679585382
transform 1 0 91872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_958
timestamp 1679585382
transform 1 0 92544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_965
timestamp 1679585382
transform 1 0 93216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_972
timestamp 1679585382
transform 1 0 93888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_979
timestamp 1679585382
transform 1 0 94560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_986
timestamp 1679585382
transform 1 0 95232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_993
timestamp 1679585382
transform 1 0 95904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1000
timestamp 1679585382
transform 1 0 96576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1007
timestamp 1679585382
transform 1 0 97248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1014
timestamp 1679585382
transform 1 0 97920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1021
timestamp 1679585382
transform 1 0 98592 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_1028
timestamp 1677583258
transform 1 0 99264 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679585382
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679585382
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679585382
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679585382
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679585382
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679585382
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679585382
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679585382
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679585382
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679585382
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679585382
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_91
timestamp 1679585382
transform 1 0 9312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_98
timestamp 1679585382
transform 1 0 9984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_105
timestamp 1679585382
transform 1 0 10656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_112
timestamp 1679585382
transform 1 0 11328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_119
timestamp 1679585382
transform 1 0 12000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_126
timestamp 1679585382
transform 1 0 12672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_133
timestamp 1679585382
transform 1 0 13344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_140
timestamp 1679585382
transform 1 0 14016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_147
timestamp 1679585382
transform 1 0 14688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_154
timestamp 1679585382
transform 1 0 15360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_161
timestamp 1679585382
transform 1 0 16032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_168
timestamp 1679585382
transform 1 0 16704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_175
timestamp 1679585382
transform 1 0 17376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_182
timestamp 1679585382
transform 1 0 18048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_189
timestamp 1679585382
transform 1 0 18720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_196
timestamp 1679585382
transform 1 0 19392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_203
timestamp 1679585382
transform 1 0 20064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_210
timestamp 1679585382
transform 1 0 20736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_217
timestamp 1679585382
transform 1 0 21408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_224
timestamp 1679585382
transform 1 0 22080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_231
timestamp 1679585382
transform 1 0 22752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_238
timestamp 1679585382
transform 1 0 23424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_245
timestamp 1679585382
transform 1 0 24096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_252
timestamp 1679585382
transform 1 0 24768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_259
timestamp 1679585382
transform 1 0 25440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_266
timestamp 1679585382
transform 1 0 26112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_273
timestamp 1679585382
transform 1 0 26784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_280
timestamp 1679585382
transform 1 0 27456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_287
timestamp 1679585382
transform 1 0 28128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_294
timestamp 1679585382
transform 1 0 28800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_301
timestamp 1679585382
transform 1 0 29472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_308
timestamp 1679585382
transform 1 0 30144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_315
timestamp 1679585382
transform 1 0 30816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_322
timestamp 1679585382
transform 1 0 31488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_329
timestamp 1679585382
transform 1 0 32160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_336
timestamp 1679585382
transform 1 0 32832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_343
timestamp 1679585382
transform 1 0 33504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_350
timestamp 1679585382
transform 1 0 34176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_357
timestamp 1679585382
transform 1 0 34848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_364
timestamp 1679585382
transform 1 0 35520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_371
timestamp 1679585382
transform 1 0 36192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_378
timestamp 1679585382
transform 1 0 36864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_385
timestamp 1679585382
transform 1 0 37536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_392
timestamp 1679585382
transform 1 0 38208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_399
timestamp 1679585382
transform 1 0 38880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_406
timestamp 1679585382
transform 1 0 39552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_413
timestamp 1679585382
transform 1 0 40224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_420
timestamp 1679585382
transform 1 0 40896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_427
timestamp 1679585382
transform 1 0 41568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_434
timestamp 1679585382
transform 1 0 42240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_441
timestamp 1679585382
transform 1 0 42912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_448
timestamp 1679585382
transform 1 0 43584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_455
timestamp 1679585382
transform 1 0 44256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_462
timestamp 1679585382
transform 1 0 44928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_469
timestamp 1679585382
transform 1 0 45600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_476
timestamp 1679585382
transform 1 0 46272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_483
timestamp 1679585382
transform 1 0 46944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_490
timestamp 1679585382
transform 1 0 47616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_497
timestamp 1679585382
transform 1 0 48288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_504
timestamp 1679585382
transform 1 0 48960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_511
timestamp 1679585382
transform 1 0 49632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_518
timestamp 1679585382
transform 1 0 50304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_525
timestamp 1679585382
transform 1 0 50976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_532
timestamp 1679585382
transform 1 0 51648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_539
timestamp 1679585382
transform 1 0 52320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_546
timestamp 1679585382
transform 1 0 52992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_553
timestamp 1679585382
transform 1 0 53664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_560
timestamp 1679585382
transform 1 0 54336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_567
timestamp 1679585382
transform 1 0 55008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_574
timestamp 1679585382
transform 1 0 55680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_581
timestamp 1679585382
transform 1 0 56352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_588
timestamp 1679585382
transform 1 0 57024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_595
timestamp 1679585382
transform 1 0 57696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_602
timestamp 1679585382
transform 1 0 58368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_609
timestamp 1679585382
transform 1 0 59040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_616
timestamp 1679585382
transform 1 0 59712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_623
timestamp 1679585382
transform 1 0 60384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_630
timestamp 1679585382
transform 1 0 61056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_637
timestamp 1679585382
transform 1 0 61728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_644
timestamp 1679585382
transform 1 0 62400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_651
timestamp 1679585382
transform 1 0 63072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_658
timestamp 1679585382
transform 1 0 63744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_665
timestamp 1679585382
transform 1 0 64416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_672
timestamp 1679585382
transform 1 0 65088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_679
timestamp 1679585382
transform 1 0 65760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_686
timestamp 1679585382
transform 1 0 66432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_693
timestamp 1679585382
transform 1 0 67104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_700
timestamp 1679585382
transform 1 0 67776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_707
timestamp 1679585382
transform 1 0 68448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_714
timestamp 1679585382
transform 1 0 69120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_721
timestamp 1679585382
transform 1 0 69792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_728
timestamp 1679585382
transform 1 0 70464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_735
timestamp 1679585382
transform 1 0 71136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_742
timestamp 1679585382
transform 1 0 71808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_749
timestamp 1679585382
transform 1 0 72480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_756
timestamp 1679585382
transform 1 0 73152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_763
timestamp 1679585382
transform 1 0 73824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_770
timestamp 1679585382
transform 1 0 74496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_777
timestamp 1679585382
transform 1 0 75168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_784
timestamp 1679585382
transform 1 0 75840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_791
timestamp 1679585382
transform 1 0 76512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_798
timestamp 1679585382
transform 1 0 77184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_805
timestamp 1679585382
transform 1 0 77856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_812
timestamp 1679585382
transform 1 0 78528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_819
timestamp 1679585382
transform 1 0 79200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_826
timestamp 1679585382
transform 1 0 79872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_833
timestamp 1679585382
transform 1 0 80544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_840
timestamp 1679585382
transform 1 0 81216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_847
timestamp 1679585382
transform 1 0 81888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_854
timestamp 1679585382
transform 1 0 82560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_861
timestamp 1679585382
transform 1 0 83232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_868
timestamp 1679585382
transform 1 0 83904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_875
timestamp 1679585382
transform 1 0 84576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_882
timestamp 1679585382
transform 1 0 85248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_889
timestamp 1679585382
transform 1 0 85920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_896
timestamp 1679585382
transform 1 0 86592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_903
timestamp 1679585382
transform 1 0 87264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_910
timestamp 1679585382
transform 1 0 87936 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_917
timestamp 1679585382
transform 1 0 88608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_924
timestamp 1679585382
transform 1 0 89280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_931
timestamp 1679585382
transform 1 0 89952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_938
timestamp 1679585382
transform 1 0 90624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_945
timestamp 1679585382
transform 1 0 91296 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_952
timestamp 1679585382
transform 1 0 91968 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_959
timestamp 1679585382
transform 1 0 92640 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_966
timestamp 1679585382
transform 1 0 93312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_973
timestamp 1679585382
transform 1 0 93984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_980
timestamp 1679585382
transform 1 0 94656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_987
timestamp 1679585382
transform 1 0 95328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_994
timestamp 1679585382
transform 1 0 96000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1001
timestamp 1679585382
transform 1 0 96672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1008
timestamp 1679585382
transform 1 0 97344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1015
timestamp 1679585382
transform 1 0 98016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1022
timestamp 1679585382
transform 1 0 98688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679585382
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679585382
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679585382
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_25
timestamp 1679585382
transform 1 0 2976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_32
timestamp 1679585382
transform 1 0 3648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_39
timestamp 1679585382
transform 1 0 4320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_46
timestamp 1679585382
transform 1 0 4992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_53
timestamp 1679585382
transform 1 0 5664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_60
timestamp 1679585382
transform 1 0 6336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_67
timestamp 1679585382
transform 1 0 7008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_87
timestamp 1679581501
transform 1 0 8928 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_91
timestamp 1677583258
transform 1 0 9312 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_101
timestamp 1679585382
transform 1 0 10272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_108
timestamp 1679585382
transform 1 0 10944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_115
timestamp 1679585382
transform 1 0 11616 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_122
timestamp 1679585382
transform 1 0 12288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_129
timestamp 1679585382
transform 1 0 12960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_136
timestamp 1679585382
transform 1 0 13632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_143
timestamp 1679585382
transform 1 0 14304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_150
timestamp 1679585382
transform 1 0 14976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_157
timestamp 1679585382
transform 1 0 15648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_164
timestamp 1679585382
transform 1 0 16320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_171
timestamp 1679585382
transform 1 0 16992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_178
timestamp 1679585382
transform 1 0 17664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_185
timestamp 1679585382
transform 1 0 18336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_192
timestamp 1679585382
transform 1 0 19008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_199
timestamp 1679585382
transform 1 0 19680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_206
timestamp 1679585382
transform 1 0 20352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_213
timestamp 1679585382
transform 1 0 21024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_220
timestamp 1679585382
transform 1 0 21696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_227
timestamp 1679585382
transform 1 0 22368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_234
timestamp 1679585382
transform 1 0 23040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_241
timestamp 1679585382
transform 1 0 23712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_248
timestamp 1679585382
transform 1 0 24384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_255
timestamp 1679585382
transform 1 0 25056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_262
timestamp 1679585382
transform 1 0 25728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_269
timestamp 1679585382
transform 1 0 26400 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_276
timestamp 1679585382
transform 1 0 27072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_283
timestamp 1679585382
transform 1 0 27744 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_290
timestamp 1679585382
transform 1 0 28416 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_297
timestamp 1679585382
transform 1 0 29088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_304
timestamp 1679585382
transform 1 0 29760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_311
timestamp 1679585382
transform 1 0 30432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_318
timestamp 1679585382
transform 1 0 31104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_325
timestamp 1679585382
transform 1 0 31776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_332
timestamp 1679585382
transform 1 0 32448 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_339
timestamp 1679585382
transform 1 0 33120 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_346
timestamp 1679585382
transform 1 0 33792 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_353
timestamp 1679585382
transform 1 0 34464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_360
timestamp 1679585382
transform 1 0 35136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_367
timestamp 1679585382
transform 1 0 35808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_374
timestamp 1679585382
transform 1 0 36480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_381
timestamp 1679585382
transform 1 0 37152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_388
timestamp 1679585382
transform 1 0 37824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_395
timestamp 1679585382
transform 1 0 38496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_402
timestamp 1679585382
transform 1 0 39168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_409
timestamp 1679585382
transform 1 0 39840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_416
timestamp 1679585382
transform 1 0 40512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_423
timestamp 1679585382
transform 1 0 41184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_430
timestamp 1679585382
transform 1 0 41856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_437
timestamp 1679585382
transform 1 0 42528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_444
timestamp 1679585382
transform 1 0 43200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_451
timestamp 1679585382
transform 1 0 43872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_458
timestamp 1679585382
transform 1 0 44544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_465
timestamp 1679585382
transform 1 0 45216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_472
timestamp 1679585382
transform 1 0 45888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_479
timestamp 1679585382
transform 1 0 46560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_486
timestamp 1679585382
transform 1 0 47232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_493
timestamp 1679585382
transform 1 0 47904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_500
timestamp 1679585382
transform 1 0 48576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_507
timestamp 1679585382
transform 1 0 49248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_514
timestamp 1679585382
transform 1 0 49920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_521
timestamp 1679585382
transform 1 0 50592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_528
timestamp 1679585382
transform 1 0 51264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_535
timestamp 1679585382
transform 1 0 51936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_542
timestamp 1679585382
transform 1 0 52608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_549
timestamp 1679585382
transform 1 0 53280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_556
timestamp 1679585382
transform 1 0 53952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_563
timestamp 1679585382
transform 1 0 54624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_570
timestamp 1679585382
transform 1 0 55296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_577
timestamp 1679585382
transform 1 0 55968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_584
timestamp 1679585382
transform 1 0 56640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_591
timestamp 1679585382
transform 1 0 57312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_598
timestamp 1679585382
transform 1 0 57984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_605
timestamp 1679585382
transform 1 0 58656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_612
timestamp 1679585382
transform 1 0 59328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_619
timestamp 1679585382
transform 1 0 60000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_626
timestamp 1679585382
transform 1 0 60672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_633
timestamp 1679585382
transform 1 0 61344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_640
timestamp 1679585382
transform 1 0 62016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_647
timestamp 1679585382
transform 1 0 62688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_654
timestamp 1679585382
transform 1 0 63360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_661
timestamp 1679585382
transform 1 0 64032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_668
timestamp 1679585382
transform 1 0 64704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_675
timestamp 1679585382
transform 1 0 65376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_682
timestamp 1679585382
transform 1 0 66048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_689
timestamp 1679585382
transform 1 0 66720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_696
timestamp 1679585382
transform 1 0 67392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_703
timestamp 1679585382
transform 1 0 68064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_710
timestamp 1679585382
transform 1 0 68736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_717
timestamp 1679585382
transform 1 0 69408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_724
timestamp 1679585382
transform 1 0 70080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_731
timestamp 1679585382
transform 1 0 70752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_738
timestamp 1679585382
transform 1 0 71424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_745
timestamp 1679585382
transform 1 0 72096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_752
timestamp 1679585382
transform 1 0 72768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_759
timestamp 1679585382
transform 1 0 73440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_766
timestamp 1679585382
transform 1 0 74112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_773
timestamp 1679585382
transform 1 0 74784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_780
timestamp 1679585382
transform 1 0 75456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_787
timestamp 1679585382
transform 1 0 76128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_794
timestamp 1679585382
transform 1 0 76800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_801
timestamp 1679585382
transform 1 0 77472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_808
timestamp 1679585382
transform 1 0 78144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_815
timestamp 1679585382
transform 1 0 78816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_822
timestamp 1679585382
transform 1 0 79488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_829
timestamp 1679585382
transform 1 0 80160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_836
timestamp 1679585382
transform 1 0 80832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_843
timestamp 1679585382
transform 1 0 81504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_850
timestamp 1679585382
transform 1 0 82176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_857
timestamp 1679585382
transform 1 0 82848 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_864
timestamp 1679585382
transform 1 0 83520 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_871
timestamp 1679585382
transform 1 0 84192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_878
timestamp 1679585382
transform 1 0 84864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_885
timestamp 1679585382
transform 1 0 85536 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_892
timestamp 1679585382
transform 1 0 86208 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_899
timestamp 1679585382
transform 1 0 86880 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_906
timestamp 1679585382
transform 1 0 87552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_913
timestamp 1679585382
transform 1 0 88224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_920
timestamp 1679585382
transform 1 0 88896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_927
timestamp 1679585382
transform 1 0 89568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_934
timestamp 1679585382
transform 1 0 90240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_941
timestamp 1679585382
transform 1 0 90912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_948
timestamp 1679585382
transform 1 0 91584 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_955
timestamp 1679585382
transform 1 0 92256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_962
timestamp 1679585382
transform 1 0 92928 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_969
timestamp 1679585382
transform 1 0 93600 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_976
timestamp 1679585382
transform 1 0 94272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_983
timestamp 1679585382
transform 1 0 94944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_990
timestamp 1679585382
transform 1 0 95616 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_997
timestamp 1679585382
transform 1 0 96288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1004
timestamp 1679585382
transform 1 0 96960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1011
timestamp 1679585382
transform 1 0 97632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1018
timestamp 1679585382
transform 1 0 98304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_1025
timestamp 1679581501
transform 1 0 98976 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679585382
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679585382
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679585382
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679585382
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_32
timestamp 1679585382
transform 1 0 3648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_39
timestamp 1679585382
transform 1 0 4320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679585382
transform 1 0 4992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_53
timestamp 1679585382
transform 1 0 5664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_60
timestamp 1679585382
transform 1 0 6336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_67
timestamp 1679581501
transform 1 0 7008 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_71
timestamp 1677583704
transform 1 0 7392 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_100
timestamp 1679585382
transform 1 0 10176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_107
timestamp 1679585382
transform 1 0 10848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_114
timestamp 1679585382
transform 1 0 11520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_121
timestamp 1679585382
transform 1 0 12192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_128
timestamp 1679585382
transform 1 0 12864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_135
timestamp 1679585382
transform 1 0 13536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_142
timestamp 1679585382
transform 1 0 14208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_149
timestamp 1679585382
transform 1 0 14880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_156
timestamp 1679585382
transform 1 0 15552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_163
timestamp 1679585382
transform 1 0 16224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_170
timestamp 1679585382
transform 1 0 16896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_177
timestamp 1679585382
transform 1 0 17568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_184
timestamp 1679585382
transform 1 0 18240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_191
timestamp 1679585382
transform 1 0 18912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_198
timestamp 1679585382
transform 1 0 19584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_205
timestamp 1679585382
transform 1 0 20256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_212
timestamp 1679585382
transform 1 0 20928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_219
timestamp 1679585382
transform 1 0 21600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_226
timestamp 1679585382
transform 1 0 22272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_233
timestamp 1679585382
transform 1 0 22944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_240
timestamp 1679585382
transform 1 0 23616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_247
timestamp 1679585382
transform 1 0 24288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_254
timestamp 1679585382
transform 1 0 24960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_261
timestamp 1679585382
transform 1 0 25632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_268
timestamp 1679585382
transform 1 0 26304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_275
timestamp 1679585382
transform 1 0 26976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_282
timestamp 1679585382
transform 1 0 27648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_289
timestamp 1679585382
transform 1 0 28320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_296
timestamp 1679585382
transform 1 0 28992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_303
timestamp 1679585382
transform 1 0 29664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_310
timestamp 1679585382
transform 1 0 30336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_317
timestamp 1679585382
transform 1 0 31008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_324
timestamp 1679585382
transform 1 0 31680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_331
timestamp 1679585382
transform 1 0 32352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_338
timestamp 1679585382
transform 1 0 33024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_345
timestamp 1679585382
transform 1 0 33696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_352
timestamp 1679585382
transform 1 0 34368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_359
timestamp 1679585382
transform 1 0 35040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_366
timestamp 1679585382
transform 1 0 35712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_373
timestamp 1679585382
transform 1 0 36384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_380
timestamp 1679585382
transform 1 0 37056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_387
timestamp 1679585382
transform 1 0 37728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_394
timestamp 1679585382
transform 1 0 38400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_401
timestamp 1679585382
transform 1 0 39072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_408
timestamp 1679585382
transform 1 0 39744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_415
timestamp 1679585382
transform 1 0 40416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_422
timestamp 1679585382
transform 1 0 41088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_429
timestamp 1679585382
transform 1 0 41760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_436
timestamp 1679585382
transform 1 0 42432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_443
timestamp 1679585382
transform 1 0 43104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_450
timestamp 1679585382
transform 1 0 43776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_457
timestamp 1679585382
transform 1 0 44448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_464
timestamp 1679585382
transform 1 0 45120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_471
timestamp 1679585382
transform 1 0 45792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_478
timestamp 1679585382
transform 1 0 46464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_485
timestamp 1679585382
transform 1 0 47136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_492
timestamp 1679585382
transform 1 0 47808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_499
timestamp 1679585382
transform 1 0 48480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_506
timestamp 1679585382
transform 1 0 49152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_513
timestamp 1679585382
transform 1 0 49824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_520
timestamp 1679585382
transform 1 0 50496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_527
timestamp 1679585382
transform 1 0 51168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_534
timestamp 1679585382
transform 1 0 51840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_541
timestamp 1679585382
transform 1 0 52512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_548
timestamp 1679585382
transform 1 0 53184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_555
timestamp 1679585382
transform 1 0 53856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_562
timestamp 1679585382
transform 1 0 54528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_569
timestamp 1679585382
transform 1 0 55200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_576
timestamp 1679585382
transform 1 0 55872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_583
timestamp 1679585382
transform 1 0 56544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_590
timestamp 1679585382
transform 1 0 57216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_597
timestamp 1679585382
transform 1 0 57888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_604
timestamp 1679585382
transform 1 0 58560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_611
timestamp 1679585382
transform 1 0 59232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_618
timestamp 1679585382
transform 1 0 59904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_625
timestamp 1679585382
transform 1 0 60576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_632
timestamp 1679585382
transform 1 0 61248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_639
timestamp 1679585382
transform 1 0 61920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_646
timestamp 1679585382
transform 1 0 62592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_653
timestamp 1679585382
transform 1 0 63264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_660
timestamp 1679585382
transform 1 0 63936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_667
timestamp 1679585382
transform 1 0 64608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_674
timestamp 1679585382
transform 1 0 65280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_681
timestamp 1679585382
transform 1 0 65952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_688
timestamp 1679585382
transform 1 0 66624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_695
timestamp 1679585382
transform 1 0 67296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_702
timestamp 1679585382
transform 1 0 67968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_709
timestamp 1679585382
transform 1 0 68640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_716
timestamp 1679585382
transform 1 0 69312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_723
timestamp 1679585382
transform 1 0 69984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_730
timestamp 1679585382
transform 1 0 70656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_737
timestamp 1679585382
transform 1 0 71328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_744
timestamp 1679585382
transform 1 0 72000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_751
timestamp 1679585382
transform 1 0 72672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_758
timestamp 1679585382
transform 1 0 73344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_765
timestamp 1679585382
transform 1 0 74016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_772
timestamp 1679585382
transform 1 0 74688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_779
timestamp 1679585382
transform 1 0 75360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_786
timestamp 1679585382
transform 1 0 76032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_793
timestamp 1679585382
transform 1 0 76704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_800
timestamp 1679585382
transform 1 0 77376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_807
timestamp 1679585382
transform 1 0 78048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_814
timestamp 1679585382
transform 1 0 78720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_821
timestamp 1679585382
transform 1 0 79392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_828
timestamp 1679585382
transform 1 0 80064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_835
timestamp 1679585382
transform 1 0 80736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_842
timestamp 1679585382
transform 1 0 81408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_849
timestamp 1679585382
transform 1 0 82080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_856
timestamp 1679585382
transform 1 0 82752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_863
timestamp 1679585382
transform 1 0 83424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_870
timestamp 1679585382
transform 1 0 84096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_877
timestamp 1679585382
transform 1 0 84768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_884
timestamp 1679585382
transform 1 0 85440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_891
timestamp 1679585382
transform 1 0 86112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_898
timestamp 1679585382
transform 1 0 86784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_905
timestamp 1679585382
transform 1 0 87456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_912
timestamp 1679585382
transform 1 0 88128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_919
timestamp 1679585382
transform 1 0 88800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_926
timestamp 1679585382
transform 1 0 89472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_933
timestamp 1679585382
transform 1 0 90144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_940
timestamp 1679585382
transform 1 0 90816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_947
timestamp 1679585382
transform 1 0 91488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_954
timestamp 1679585382
transform 1 0 92160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_961
timestamp 1679585382
transform 1 0 92832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_968
timestamp 1679585382
transform 1 0 93504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_975
timestamp 1679585382
transform 1 0 94176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_982
timestamp 1679585382
transform 1 0 94848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_989
timestamp 1679585382
transform 1 0 95520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_996
timestamp 1679585382
transform 1 0 96192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1003
timestamp 1679585382
transform 1 0 96864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1010
timestamp 1679585382
transform 1 0 97536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1017
timestamp 1679585382
transform 1 0 98208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_1024
timestamp 1679581501
transform 1 0 98880 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_1028
timestamp 1677583258
transform 1 0 99264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679585382
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_11
timestamp 1679585382
transform 1 0 1632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_18
timestamp 1679585382
transform 1 0 2304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_25
timestamp 1679585382
transform 1 0 2976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_32
timestamp 1679585382
transform 1 0 3648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_39
timestamp 1679585382
transform 1 0 4320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_46
timestamp 1679585382
transform 1 0 4992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_53
timestamp 1679585382
transform 1 0 5664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_60
timestamp 1679585382
transform 1 0 6336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_67
timestamp 1679585382
transform 1 0 7008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_74
timestamp 1679585382
transform 1 0 7680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_81
timestamp 1679585382
transform 1 0 8352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_88
timestamp 1679585382
transform 1 0 9024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_95
timestamp 1679585382
transform 1 0 9696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_102
timestamp 1679585382
transform 1 0 10368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_109
timestamp 1679585382
transform 1 0 11040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_116
timestamp 1679585382
transform 1 0 11712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_123
timestamp 1679585382
transform 1 0 12384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_130
timestamp 1679585382
transform 1 0 13056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_137
timestamp 1679585382
transform 1 0 13728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_144
timestamp 1679585382
transform 1 0 14400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_151
timestamp 1679585382
transform 1 0 15072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_158
timestamp 1679585382
transform 1 0 15744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_165
timestamp 1679585382
transform 1 0 16416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_172
timestamp 1679585382
transform 1 0 17088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_179
timestamp 1679585382
transform 1 0 17760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_186
timestamp 1679585382
transform 1 0 18432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_193
timestamp 1679585382
transform 1 0 19104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_200
timestamp 1679585382
transform 1 0 19776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_207
timestamp 1679585382
transform 1 0 20448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_214
timestamp 1679585382
transform 1 0 21120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_221
timestamp 1679585382
transform 1 0 21792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_228
timestamp 1679585382
transform 1 0 22464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_235
timestamp 1679585382
transform 1 0 23136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_242
timestamp 1679585382
transform 1 0 23808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_249
timestamp 1679585382
transform 1 0 24480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_256
timestamp 1679585382
transform 1 0 25152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_263
timestamp 1679585382
transform 1 0 25824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_270
timestamp 1679585382
transform 1 0 26496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_277
timestamp 1679585382
transform 1 0 27168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_284
timestamp 1679585382
transform 1 0 27840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_291
timestamp 1679585382
transform 1 0 28512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_298
timestamp 1679585382
transform 1 0 29184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_305
timestamp 1679585382
transform 1 0 29856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_312
timestamp 1679585382
transform 1 0 30528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_319
timestamp 1679585382
transform 1 0 31200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_326
timestamp 1679585382
transform 1 0 31872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_333
timestamp 1679585382
transform 1 0 32544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_340
timestamp 1679585382
transform 1 0 33216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_347
timestamp 1679585382
transform 1 0 33888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_354
timestamp 1679585382
transform 1 0 34560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_361
timestamp 1679585382
transform 1 0 35232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_368
timestamp 1679585382
transform 1 0 35904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_375
timestamp 1679585382
transform 1 0 36576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_382
timestamp 1679585382
transform 1 0 37248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_389
timestamp 1679585382
transform 1 0 37920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_396
timestamp 1679585382
transform 1 0 38592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_403
timestamp 1679585382
transform 1 0 39264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_410
timestamp 1679585382
transform 1 0 39936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_417
timestamp 1679585382
transform 1 0 40608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_424
timestamp 1679585382
transform 1 0 41280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_431
timestamp 1679585382
transform 1 0 41952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_438
timestamp 1679585382
transform 1 0 42624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_445
timestamp 1679585382
transform 1 0 43296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_452
timestamp 1679585382
transform 1 0 43968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_459
timestamp 1679585382
transform 1 0 44640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_466
timestamp 1679585382
transform 1 0 45312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_473
timestamp 1679585382
transform 1 0 45984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_480
timestamp 1679585382
transform 1 0 46656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_487
timestamp 1679585382
transform 1 0 47328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_494
timestamp 1679585382
transform 1 0 48000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_501
timestamp 1679585382
transform 1 0 48672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_508
timestamp 1679585382
transform 1 0 49344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_515
timestamp 1679585382
transform 1 0 50016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_522
timestamp 1679585382
transform 1 0 50688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_529
timestamp 1679585382
transform 1 0 51360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_536
timestamp 1679585382
transform 1 0 52032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_543
timestamp 1679585382
transform 1 0 52704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_550
timestamp 1679585382
transform 1 0 53376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_557
timestamp 1679585382
transform 1 0 54048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_564
timestamp 1679585382
transform 1 0 54720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_571
timestamp 1679585382
transform 1 0 55392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_578
timestamp 1679585382
transform 1 0 56064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_585
timestamp 1679585382
transform 1 0 56736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_592
timestamp 1679585382
transform 1 0 57408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_599
timestamp 1679585382
transform 1 0 58080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_606
timestamp 1679585382
transform 1 0 58752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_613
timestamp 1679585382
transform 1 0 59424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_620
timestamp 1679585382
transform 1 0 60096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_627
timestamp 1679585382
transform 1 0 60768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_634
timestamp 1679585382
transform 1 0 61440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_641
timestamp 1679585382
transform 1 0 62112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_648
timestamp 1679585382
transform 1 0 62784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_655
timestamp 1679585382
transform 1 0 63456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_662
timestamp 1679585382
transform 1 0 64128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_669
timestamp 1679585382
transform 1 0 64800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_676
timestamp 1679585382
transform 1 0 65472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_683
timestamp 1679585382
transform 1 0 66144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_690
timestamp 1679585382
transform 1 0 66816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_697
timestamp 1679585382
transform 1 0 67488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_704
timestamp 1679585382
transform 1 0 68160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_711
timestamp 1679585382
transform 1 0 68832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_718
timestamp 1679585382
transform 1 0 69504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_725
timestamp 1679585382
transform 1 0 70176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_732
timestamp 1679585382
transform 1 0 70848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_739
timestamp 1679585382
transform 1 0 71520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_746
timestamp 1679585382
transform 1 0 72192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_753
timestamp 1679585382
transform 1 0 72864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_760
timestamp 1679585382
transform 1 0 73536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_767
timestamp 1679585382
transform 1 0 74208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_774
timestamp 1679585382
transform 1 0 74880 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_781
timestamp 1679585382
transform 1 0 75552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_788
timestamp 1679585382
transform 1 0 76224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_795
timestamp 1679585382
transform 1 0 76896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_802
timestamp 1679585382
transform 1 0 77568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_809
timestamp 1679585382
transform 1 0 78240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_816
timestamp 1679585382
transform 1 0 78912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_823
timestamp 1679585382
transform 1 0 79584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_830
timestamp 1679585382
transform 1 0 80256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_837
timestamp 1679585382
transform 1 0 80928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_844
timestamp 1679585382
transform 1 0 81600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_851
timestamp 1679585382
transform 1 0 82272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_858
timestamp 1679585382
transform 1 0 82944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_865
timestamp 1679585382
transform 1 0 83616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_872
timestamp 1679585382
transform 1 0 84288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_879
timestamp 1679585382
transform 1 0 84960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_886
timestamp 1679585382
transform 1 0 85632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_893
timestamp 1679585382
transform 1 0 86304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_900
timestamp 1679585382
transform 1 0 86976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_907
timestamp 1679585382
transform 1 0 87648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_914
timestamp 1679585382
transform 1 0 88320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_921
timestamp 1679585382
transform 1 0 88992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_928
timestamp 1679585382
transform 1 0 89664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_935
timestamp 1679585382
transform 1 0 90336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_942
timestamp 1679585382
transform 1 0 91008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_949
timestamp 1679585382
transform 1 0 91680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_956
timestamp 1679585382
transform 1 0 92352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_963
timestamp 1679585382
transform 1 0 93024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_970
timestamp 1679585382
transform 1 0 93696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_977
timestamp 1679585382
transform 1 0 94368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_984
timestamp 1679585382
transform 1 0 95040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_991
timestamp 1679585382
transform 1 0 95712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_998
timestamp 1679585382
transform 1 0 96384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1005
timestamp 1679585382
transform 1 0 97056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1012
timestamp 1679585382
transform 1 0 97728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1019
timestamp 1679585382
transform 1 0 98400 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_1026
timestamp 1677583704
transform 1 0 99072 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_1028
timestamp 1677583258
transform 1 0 99264 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679585382
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679585382
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679585382
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679585382
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679585382
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679585382
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679585382
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679585382
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_60
timestamp 1679585382
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_67
timestamp 1679585382
transform 1 0 7008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_74
timestamp 1679585382
transform 1 0 7680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_81
timestamp 1679585382
transform 1 0 8352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_88
timestamp 1679585382
transform 1 0 9024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_95
timestamp 1679585382
transform 1 0 9696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_102
timestamp 1679585382
transform 1 0 10368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_109
timestamp 1679585382
transform 1 0 11040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_116
timestamp 1679585382
transform 1 0 11712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_123
timestamp 1679585382
transform 1 0 12384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_130
timestamp 1679585382
transform 1 0 13056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_137
timestamp 1679585382
transform 1 0 13728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_144
timestamp 1679585382
transform 1 0 14400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_151
timestamp 1679585382
transform 1 0 15072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_158
timestamp 1679585382
transform 1 0 15744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_165
timestamp 1679585382
transform 1 0 16416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_172
timestamp 1679585382
transform 1 0 17088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_179
timestamp 1679585382
transform 1 0 17760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_186
timestamp 1679585382
transform 1 0 18432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_193
timestamp 1679585382
transform 1 0 19104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_200
timestamp 1679585382
transform 1 0 19776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_207
timestamp 1679585382
transform 1 0 20448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_214
timestamp 1679585382
transform 1 0 21120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_221
timestamp 1679585382
transform 1 0 21792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_228
timestamp 1679585382
transform 1 0 22464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_235
timestamp 1679585382
transform 1 0 23136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_242
timestamp 1679585382
transform 1 0 23808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_249
timestamp 1679585382
transform 1 0 24480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_256
timestamp 1679585382
transform 1 0 25152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_263
timestamp 1679585382
transform 1 0 25824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_270
timestamp 1679585382
transform 1 0 26496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_277
timestamp 1679585382
transform 1 0 27168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_284
timestamp 1679585382
transform 1 0 27840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_291
timestamp 1679585382
transform 1 0 28512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_298
timestamp 1679585382
transform 1 0 29184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_305
timestamp 1679585382
transform 1 0 29856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_312
timestamp 1679585382
transform 1 0 30528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_319
timestamp 1679585382
transform 1 0 31200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_326
timestamp 1679585382
transform 1 0 31872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_333
timestamp 1679585382
transform 1 0 32544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_340
timestamp 1679585382
transform 1 0 33216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_347
timestamp 1679585382
transform 1 0 33888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_354
timestamp 1679585382
transform 1 0 34560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_361
timestamp 1679585382
transform 1 0 35232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_368
timestamp 1679585382
transform 1 0 35904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_375
timestamp 1679585382
transform 1 0 36576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_382
timestamp 1679585382
transform 1 0 37248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_389
timestamp 1679585382
transform 1 0 37920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_396
timestamp 1679585382
transform 1 0 38592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_403
timestamp 1679585382
transform 1 0 39264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_410
timestamp 1679585382
transform 1 0 39936 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_417
timestamp 1679585382
transform 1 0 40608 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_424
timestamp 1679585382
transform 1 0 41280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_431
timestamp 1679585382
transform 1 0 41952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_438
timestamp 1679585382
transform 1 0 42624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_445
timestamp 1679585382
transform 1 0 43296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_452
timestamp 1679585382
transform 1 0 43968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_459
timestamp 1679585382
transform 1 0 44640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_466
timestamp 1679585382
transform 1 0 45312 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_473
timestamp 1679585382
transform 1 0 45984 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_480
timestamp 1679585382
transform 1 0 46656 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_487
timestamp 1679585382
transform 1 0 47328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_494
timestamp 1679585382
transform 1 0 48000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_501
timestamp 1679585382
transform 1 0 48672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_508
timestamp 1679585382
transform 1 0 49344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_515
timestamp 1679585382
transform 1 0 50016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_522
timestamp 1679585382
transform 1 0 50688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_529
timestamp 1679585382
transform 1 0 51360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_536
timestamp 1679585382
transform 1 0 52032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_543
timestamp 1679585382
transform 1 0 52704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_550
timestamp 1679585382
transform 1 0 53376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_557
timestamp 1679585382
transform 1 0 54048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_564
timestamp 1679585382
transform 1 0 54720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_571
timestamp 1679585382
transform 1 0 55392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_578
timestamp 1679585382
transform 1 0 56064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_585
timestamp 1679585382
transform 1 0 56736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_592
timestamp 1679585382
transform 1 0 57408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_599
timestamp 1679585382
transform 1 0 58080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_606
timestamp 1679585382
transform 1 0 58752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_613
timestamp 1679585382
transform 1 0 59424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_620
timestamp 1679585382
transform 1 0 60096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_627
timestamp 1679585382
transform 1 0 60768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_634
timestamp 1679585382
transform 1 0 61440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_641
timestamp 1679585382
transform 1 0 62112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_648
timestamp 1679585382
transform 1 0 62784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_655
timestamp 1679585382
transform 1 0 63456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_662
timestamp 1679585382
transform 1 0 64128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_669
timestamp 1679585382
transform 1 0 64800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_676
timestamp 1679585382
transform 1 0 65472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_683
timestamp 1679585382
transform 1 0 66144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_690
timestamp 1679585382
transform 1 0 66816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_697
timestamp 1679585382
transform 1 0 67488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_704
timestamp 1679585382
transform 1 0 68160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_711
timestamp 1679585382
transform 1 0 68832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_718
timestamp 1679585382
transform 1 0 69504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_725
timestamp 1679585382
transform 1 0 70176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_732
timestamp 1679585382
transform 1 0 70848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_739
timestamp 1679585382
transform 1 0 71520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_746
timestamp 1679585382
transform 1 0 72192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_753
timestamp 1679585382
transform 1 0 72864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_760
timestamp 1679585382
transform 1 0 73536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_767
timestamp 1679585382
transform 1 0 74208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_774
timestamp 1679585382
transform 1 0 74880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_781
timestamp 1679585382
transform 1 0 75552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_788
timestamp 1679585382
transform 1 0 76224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_795
timestamp 1679585382
transform 1 0 76896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_802
timestamp 1679585382
transform 1 0 77568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_809
timestamp 1679585382
transform 1 0 78240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_816
timestamp 1679585382
transform 1 0 78912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_823
timestamp 1679585382
transform 1 0 79584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_830
timestamp 1679585382
transform 1 0 80256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_837
timestamp 1679585382
transform 1 0 80928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_844
timestamp 1679585382
transform 1 0 81600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_851
timestamp 1679585382
transform 1 0 82272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_858
timestamp 1679585382
transform 1 0 82944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_865
timestamp 1679585382
transform 1 0 83616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_872
timestamp 1679585382
transform 1 0 84288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_879
timestamp 1679585382
transform 1 0 84960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_886
timestamp 1679585382
transform 1 0 85632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_893
timestamp 1679585382
transform 1 0 86304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_900
timestamp 1679585382
transform 1 0 86976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_907
timestamp 1679585382
transform 1 0 87648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_914
timestamp 1679585382
transform 1 0 88320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_921
timestamp 1679585382
transform 1 0 88992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_928
timestamp 1679585382
transform 1 0 89664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_935
timestamp 1679585382
transform 1 0 90336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_942
timestamp 1679585382
transform 1 0 91008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_949
timestamp 1679585382
transform 1 0 91680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_956
timestamp 1679585382
transform 1 0 92352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_963
timestamp 1679585382
transform 1 0 93024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_970
timestamp 1679585382
transform 1 0 93696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_977
timestamp 1679585382
transform 1 0 94368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_984
timestamp 1679585382
transform 1 0 95040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_991
timestamp 1679585382
transform 1 0 95712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_998
timestamp 1679585382
transform 1 0 96384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1005
timestamp 1679585382
transform 1 0 97056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1012
timestamp 1679585382
transform 1 0 97728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1019
timestamp 1679585382
transform 1 0 98400 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_1026
timestamp 1677583704
transform 1 0 99072 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_1028
timestamp 1677583258
transform 1 0 99264 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679585382
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679585382
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679585382
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679585382
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679585382
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_39
timestamp 1679585382
transform 1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_46
timestamp 1679585382
transform 1 0 4992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_53
timestamp 1679585382
transform 1 0 5664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_60
timestamp 1679585382
transform 1 0 6336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_67
timestamp 1679585382
transform 1 0 7008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_74
timestamp 1679585382
transform 1 0 7680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_81
timestamp 1679585382
transform 1 0 8352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_88
timestamp 1679585382
transform 1 0 9024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_95
timestamp 1679585382
transform 1 0 9696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_102
timestamp 1679585382
transform 1 0 10368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_109
timestamp 1679585382
transform 1 0 11040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_116
timestamp 1679585382
transform 1 0 11712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_123
timestamp 1679585382
transform 1 0 12384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_130
timestamp 1679585382
transform 1 0 13056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_137
timestamp 1679585382
transform 1 0 13728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_144
timestamp 1679585382
transform 1 0 14400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_151
timestamp 1679585382
transform 1 0 15072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_158
timestamp 1679585382
transform 1 0 15744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_165
timestamp 1679585382
transform 1 0 16416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_172
timestamp 1679585382
transform 1 0 17088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_179
timestamp 1679585382
transform 1 0 17760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_186
timestamp 1679585382
transform 1 0 18432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_193
timestamp 1679585382
transform 1 0 19104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_200
timestamp 1679585382
transform 1 0 19776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_207
timestamp 1679585382
transform 1 0 20448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_214
timestamp 1679585382
transform 1 0 21120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_221
timestamp 1679585382
transform 1 0 21792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_228
timestamp 1679585382
transform 1 0 22464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_235
timestamp 1679585382
transform 1 0 23136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_242
timestamp 1679585382
transform 1 0 23808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_249
timestamp 1679585382
transform 1 0 24480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_256
timestamp 1679585382
transform 1 0 25152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_263
timestamp 1679585382
transform 1 0 25824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_270
timestamp 1679585382
transform 1 0 26496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_277
timestamp 1679585382
transform 1 0 27168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_284
timestamp 1679585382
transform 1 0 27840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_291
timestamp 1679585382
transform 1 0 28512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_298
timestamp 1679585382
transform 1 0 29184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_305
timestamp 1679585382
transform 1 0 29856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_312
timestamp 1679585382
transform 1 0 30528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_319
timestamp 1679585382
transform 1 0 31200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_326
timestamp 1679585382
transform 1 0 31872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_333
timestamp 1679585382
transform 1 0 32544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_340
timestamp 1679585382
transform 1 0 33216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_347
timestamp 1679585382
transform 1 0 33888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_354
timestamp 1679585382
transform 1 0 34560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_361
timestamp 1679585382
transform 1 0 35232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_368
timestamp 1679585382
transform 1 0 35904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_375
timestamp 1679585382
transform 1 0 36576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_382
timestamp 1679585382
transform 1 0 37248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_389
timestamp 1679585382
transform 1 0 37920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_396
timestamp 1679585382
transform 1 0 38592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_403
timestamp 1679585382
transform 1 0 39264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_410
timestamp 1679585382
transform 1 0 39936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_417
timestamp 1679585382
transform 1 0 40608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_424
timestamp 1679585382
transform 1 0 41280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_431
timestamp 1679585382
transform 1 0 41952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_438
timestamp 1679585382
transform 1 0 42624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_445
timestamp 1679585382
transform 1 0 43296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_452
timestamp 1679585382
transform 1 0 43968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_459
timestamp 1679585382
transform 1 0 44640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_466
timestamp 1679585382
transform 1 0 45312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_473
timestamp 1679585382
transform 1 0 45984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_480
timestamp 1679585382
transform 1 0 46656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_487
timestamp 1679585382
transform 1 0 47328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_494
timestamp 1679585382
transform 1 0 48000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_501
timestamp 1679585382
transform 1 0 48672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_508
timestamp 1679585382
transform 1 0 49344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_515
timestamp 1679585382
transform 1 0 50016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_522
timestamp 1679585382
transform 1 0 50688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_529
timestamp 1679585382
transform 1 0 51360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_536
timestamp 1679585382
transform 1 0 52032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_543
timestamp 1679585382
transform 1 0 52704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_550
timestamp 1679585382
transform 1 0 53376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_557
timestamp 1679585382
transform 1 0 54048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_564
timestamp 1679585382
transform 1 0 54720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_571
timestamp 1679585382
transform 1 0 55392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_578
timestamp 1679585382
transform 1 0 56064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_585
timestamp 1679585382
transform 1 0 56736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_592
timestamp 1679585382
transform 1 0 57408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_599
timestamp 1679585382
transform 1 0 58080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_606
timestamp 1679585382
transform 1 0 58752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_613
timestamp 1679585382
transform 1 0 59424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_620
timestamp 1679585382
transform 1 0 60096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_627
timestamp 1679585382
transform 1 0 60768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_634
timestamp 1679585382
transform 1 0 61440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_641
timestamp 1679585382
transform 1 0 62112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_648
timestamp 1679585382
transform 1 0 62784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_655
timestamp 1679585382
transform 1 0 63456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_662
timestamp 1679585382
transform 1 0 64128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_669
timestamp 1679585382
transform 1 0 64800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_676
timestamp 1679585382
transform 1 0 65472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_683
timestamp 1679585382
transform 1 0 66144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_690
timestamp 1679585382
transform 1 0 66816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_697
timestamp 1679585382
transform 1 0 67488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_704
timestamp 1679585382
transform 1 0 68160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_711
timestamp 1679585382
transform 1 0 68832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_718
timestamp 1679585382
transform 1 0 69504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_725
timestamp 1679585382
transform 1 0 70176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_732
timestamp 1679585382
transform 1 0 70848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_739
timestamp 1679585382
transform 1 0 71520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_746
timestamp 1679585382
transform 1 0 72192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_753
timestamp 1679585382
transform 1 0 72864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_760
timestamp 1679585382
transform 1 0 73536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_767
timestamp 1679585382
transform 1 0 74208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_774
timestamp 1679585382
transform 1 0 74880 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_781
timestamp 1679585382
transform 1 0 75552 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_788
timestamp 1679585382
transform 1 0 76224 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_795
timestamp 1679585382
transform 1 0 76896 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_802
timestamp 1679585382
transform 1 0 77568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_809
timestamp 1679585382
transform 1 0 78240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_816
timestamp 1679585382
transform 1 0 78912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_823
timestamp 1679585382
transform 1 0 79584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_830
timestamp 1679585382
transform 1 0 80256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_837
timestamp 1679585382
transform 1 0 80928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_844
timestamp 1679585382
transform 1 0 81600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_851
timestamp 1679585382
transform 1 0 82272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_858
timestamp 1679585382
transform 1 0 82944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_865
timestamp 1679585382
transform 1 0 83616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_872
timestamp 1679585382
transform 1 0 84288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_879
timestamp 1679585382
transform 1 0 84960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_886
timestamp 1679585382
transform 1 0 85632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_893
timestamp 1679585382
transform 1 0 86304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_900
timestamp 1679585382
transform 1 0 86976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_907
timestamp 1679585382
transform 1 0 87648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_914
timestamp 1679585382
transform 1 0 88320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_921
timestamp 1679585382
transform 1 0 88992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_928
timestamp 1679585382
transform 1 0 89664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_935
timestamp 1679585382
transform 1 0 90336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_942
timestamp 1679585382
transform 1 0 91008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_949
timestamp 1679585382
transform 1 0 91680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_956
timestamp 1679585382
transform 1 0 92352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_963
timestamp 1679585382
transform 1 0 93024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_970
timestamp 1679585382
transform 1 0 93696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_977
timestamp 1679585382
transform 1 0 94368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_984
timestamp 1679585382
transform 1 0 95040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_991
timestamp 1679585382
transform 1 0 95712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_998
timestamp 1679585382
transform 1 0 96384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1005
timestamp 1679585382
transform 1 0 97056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1012
timestamp 1679585382
transform 1 0 97728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1019
timestamp 1679585382
transform 1 0 98400 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_1026
timestamp 1677583704
transform 1 0 99072 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_1028
timestamp 1677583258
transform 1 0 99264 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679585382
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679585382
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_18
timestamp 1677583704
transform 1 0 2304 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_25
timestamp 1677583704
transform 1 0 2976 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679585382
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_39
timestamp 1679585382
transform 1 0 4320 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_46
timestamp 1677583258
transform 1 0 4992 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_60
timestamp 1679585382
transform 1 0 6336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1679585382
transform 1 0 7008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_74
timestamp 1679585382
transform 1 0 7680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_81
timestamp 1679585382
transform 1 0 8352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679585382
transform 1 0 9024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_95
timestamp 1679585382
transform 1 0 9696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_102
timestamp 1679585382
transform 1 0 10368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_109
timestamp 1679585382
transform 1 0 11040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_116
timestamp 1679585382
transform 1 0 11712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_123
timestamp 1679585382
transform 1 0 12384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_130
timestamp 1679585382
transform 1 0 13056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_137
timestamp 1679585382
transform 1 0 13728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_144
timestamp 1679585382
transform 1 0 14400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_151
timestamp 1679585382
transform 1 0 15072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_158
timestamp 1679585382
transform 1 0 15744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1679585382
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_172
timestamp 1679585382
transform 1 0 17088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_179
timestamp 1679585382
transform 1 0 17760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1679585382
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_193
timestamp 1679585382
transform 1 0 19104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_200
timestamp 1679585382
transform 1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_207
timestamp 1679585382
transform 1 0 20448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_214
timestamp 1679585382
transform 1 0 21120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_221
timestamp 1679585382
transform 1 0 21792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_228
timestamp 1679585382
transform 1 0 22464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_235
timestamp 1679585382
transform 1 0 23136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_242
timestamp 1679585382
transform 1 0 23808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_249
timestamp 1679585382
transform 1 0 24480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_256
timestamp 1679585382
transform 1 0 25152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_263
timestamp 1679585382
transform 1 0 25824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_270
timestamp 1679585382
transform 1 0 26496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_277
timestamp 1679585382
transform 1 0 27168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_284
timestamp 1679585382
transform 1 0 27840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_291
timestamp 1679585382
transform 1 0 28512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_298
timestamp 1679585382
transform 1 0 29184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_305
timestamp 1679585382
transform 1 0 29856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_312
timestamp 1679585382
transform 1 0 30528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_319
timestamp 1679585382
transform 1 0 31200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_326
timestamp 1679585382
transform 1 0 31872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_333
timestamp 1679585382
transform 1 0 32544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_340
timestamp 1679585382
transform 1 0 33216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_347
timestamp 1679585382
transform 1 0 33888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_354
timestamp 1679585382
transform 1 0 34560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_361
timestamp 1679585382
transform 1 0 35232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_368
timestamp 1679585382
transform 1 0 35904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_375
timestamp 1679585382
transform 1 0 36576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_382
timestamp 1679585382
transform 1 0 37248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_389
timestamp 1679585382
transform 1 0 37920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_396
timestamp 1679585382
transform 1 0 38592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_403
timestamp 1679585382
transform 1 0 39264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_410
timestamp 1679585382
transform 1 0 39936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_417
timestamp 1679585382
transform 1 0 40608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_424
timestamp 1679585382
transform 1 0 41280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_431
timestamp 1679585382
transform 1 0 41952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_438
timestamp 1679585382
transform 1 0 42624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_445
timestamp 1679585382
transform 1 0 43296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_452
timestamp 1679585382
transform 1 0 43968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_459
timestamp 1679585382
transform 1 0 44640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_466
timestamp 1679585382
transform 1 0 45312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_473
timestamp 1679585382
transform 1 0 45984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_480
timestamp 1679585382
transform 1 0 46656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_487
timestamp 1679585382
transform 1 0 47328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_494
timestamp 1679585382
transform 1 0 48000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_501
timestamp 1679585382
transform 1 0 48672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_508
timestamp 1679585382
transform 1 0 49344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_515
timestamp 1679585382
transform 1 0 50016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_522
timestamp 1679585382
transform 1 0 50688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_529
timestamp 1679585382
transform 1 0 51360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_536
timestamp 1679585382
transform 1 0 52032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_543
timestamp 1679585382
transform 1 0 52704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_550
timestamp 1679585382
transform 1 0 53376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_557
timestamp 1679585382
transform 1 0 54048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_564
timestamp 1679585382
transform 1 0 54720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_571
timestamp 1679585382
transform 1 0 55392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_578
timestamp 1679585382
transform 1 0 56064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_585
timestamp 1679585382
transform 1 0 56736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_592
timestamp 1679585382
transform 1 0 57408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_599
timestamp 1679585382
transform 1 0 58080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_606
timestamp 1679585382
transform 1 0 58752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_613
timestamp 1679585382
transform 1 0 59424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_620
timestamp 1679585382
transform 1 0 60096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_627
timestamp 1679585382
transform 1 0 60768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_634
timestamp 1679585382
transform 1 0 61440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_641
timestamp 1679585382
transform 1 0 62112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_648
timestamp 1679585382
transform 1 0 62784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_655
timestamp 1679585382
transform 1 0 63456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_662
timestamp 1679585382
transform 1 0 64128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_669
timestamp 1679585382
transform 1 0 64800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_676
timestamp 1679585382
transform 1 0 65472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_683
timestamp 1679585382
transform 1 0 66144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_690
timestamp 1679585382
transform 1 0 66816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_697
timestamp 1679585382
transform 1 0 67488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_704
timestamp 1679585382
transform 1 0 68160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_711
timestamp 1679585382
transform 1 0 68832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_718
timestamp 1679585382
transform 1 0 69504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_725
timestamp 1679585382
transform 1 0 70176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_732
timestamp 1679585382
transform 1 0 70848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_739
timestamp 1679585382
transform 1 0 71520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_746
timestamp 1679585382
transform 1 0 72192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_753
timestamp 1679585382
transform 1 0 72864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_760
timestamp 1679585382
transform 1 0 73536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_767
timestamp 1679585382
transform 1 0 74208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_774
timestamp 1679585382
transform 1 0 74880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_781
timestamp 1679585382
transform 1 0 75552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_788
timestamp 1679585382
transform 1 0 76224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_795
timestamp 1679585382
transform 1 0 76896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_802
timestamp 1679585382
transform 1 0 77568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_809
timestamp 1679585382
transform 1 0 78240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_816
timestamp 1679585382
transform 1 0 78912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_823
timestamp 1679585382
transform 1 0 79584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_830
timestamp 1679585382
transform 1 0 80256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_837
timestamp 1679585382
transform 1 0 80928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_844
timestamp 1679585382
transform 1 0 81600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_851
timestamp 1679585382
transform 1 0 82272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_858
timestamp 1679585382
transform 1 0 82944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_865
timestamp 1679585382
transform 1 0 83616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_872
timestamp 1679585382
transform 1 0 84288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_879
timestamp 1679585382
transform 1 0 84960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_886
timestamp 1679585382
transform 1 0 85632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_893
timestamp 1679585382
transform 1 0 86304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_900
timestamp 1679585382
transform 1 0 86976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_907
timestamp 1679585382
transform 1 0 87648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_914
timestamp 1679585382
transform 1 0 88320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_921
timestamp 1679585382
transform 1 0 88992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_928
timestamp 1679585382
transform 1 0 89664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_935
timestamp 1679585382
transform 1 0 90336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_942
timestamp 1679585382
transform 1 0 91008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_949
timestamp 1679585382
transform 1 0 91680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_956
timestamp 1679585382
transform 1 0 92352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_963
timestamp 1679585382
transform 1 0 93024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_970
timestamp 1679585382
transform 1 0 93696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_977
timestamp 1679585382
transform 1 0 94368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_984
timestamp 1679585382
transform 1 0 95040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_991
timestamp 1679585382
transform 1 0 95712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_998
timestamp 1679585382
transform 1 0 96384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1005
timestamp 1679585382
transform 1 0 97056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1012
timestamp 1679585382
transform 1 0 97728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1019
timestamp 1679585382
transform 1 0 98400 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_1026
timestamp 1677583704
transform 1 0 99072 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_1028
timestamp 1677583258
transform 1 0 99264 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679585382
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679585382
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679585382
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679585382
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679585382
transform 1 0 3264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679585382
transform 1 0 3936 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_42
timestamp 1677583704
transform 1 0 4608 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_44
timestamp 1677583258
transform 1 0 4800 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_72
timestamp 1679585382
transform 1 0 7488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_79
timestamp 1679585382
transform 1 0 8160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_86
timestamp 1679585382
transform 1 0 8832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_93
timestamp 1679585382
transform 1 0 9504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_100
timestamp 1679585382
transform 1 0 10176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_107
timestamp 1679585382
transform 1 0 10848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_114
timestamp 1679585382
transform 1 0 11520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_121
timestamp 1679585382
transform 1 0 12192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_128
timestamp 1679585382
transform 1 0 12864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_135
timestamp 1679585382
transform 1 0 13536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_142
timestamp 1679585382
transform 1 0 14208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_149
timestamp 1679585382
transform 1 0 14880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_156
timestamp 1679585382
transform 1 0 15552 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_163
timestamp 1679585382
transform 1 0 16224 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_170
timestamp 1679585382
transform 1 0 16896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_177
timestamp 1679585382
transform 1 0 17568 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_184
timestamp 1679585382
transform 1 0 18240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_191
timestamp 1679585382
transform 1 0 18912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_198
timestamp 1679585382
transform 1 0 19584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_205
timestamp 1679585382
transform 1 0 20256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_212
timestamp 1679585382
transform 1 0 20928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_219
timestamp 1679585382
transform 1 0 21600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_226
timestamp 1679585382
transform 1 0 22272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_233
timestamp 1679585382
transform 1 0 22944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_240
timestamp 1679585382
transform 1 0 23616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_247
timestamp 1679585382
transform 1 0 24288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_254
timestamp 1679585382
transform 1 0 24960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_261
timestamp 1679585382
transform 1 0 25632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_268
timestamp 1679585382
transform 1 0 26304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_275
timestamp 1679585382
transform 1 0 26976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_282
timestamp 1679585382
transform 1 0 27648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_289
timestamp 1679585382
transform 1 0 28320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_296
timestamp 1679585382
transform 1 0 28992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_303
timestamp 1679585382
transform 1 0 29664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_310
timestamp 1679585382
transform 1 0 30336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_317
timestamp 1679585382
transform 1 0 31008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_324
timestamp 1679585382
transform 1 0 31680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_331
timestamp 1679585382
transform 1 0 32352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_338
timestamp 1679585382
transform 1 0 33024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_345
timestamp 1679585382
transform 1 0 33696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_352
timestamp 1679585382
transform 1 0 34368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_359
timestamp 1679585382
transform 1 0 35040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_366
timestamp 1679585382
transform 1 0 35712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_373
timestamp 1679585382
transform 1 0 36384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_380
timestamp 1679585382
transform 1 0 37056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_387
timestamp 1679585382
transform 1 0 37728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_394
timestamp 1679585382
transform 1 0 38400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_401
timestamp 1679585382
transform 1 0 39072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_408
timestamp 1679585382
transform 1 0 39744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_415
timestamp 1679585382
transform 1 0 40416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_422
timestamp 1679585382
transform 1 0 41088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_429
timestamp 1679585382
transform 1 0 41760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_436
timestamp 1679585382
transform 1 0 42432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_443
timestamp 1679585382
transform 1 0 43104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_450
timestamp 1679585382
transform 1 0 43776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_457
timestamp 1679585382
transform 1 0 44448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_464
timestamp 1679585382
transform 1 0 45120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_471
timestamp 1679585382
transform 1 0 45792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_478
timestamp 1679585382
transform 1 0 46464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_485
timestamp 1679585382
transform 1 0 47136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_492
timestamp 1679585382
transform 1 0 47808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_499
timestamp 1679585382
transform 1 0 48480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_506
timestamp 1679585382
transform 1 0 49152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_513
timestamp 1679585382
transform 1 0 49824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_520
timestamp 1679585382
transform 1 0 50496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_527
timestamp 1679585382
transform 1 0 51168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_534
timestamp 1679585382
transform 1 0 51840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_541
timestamp 1679585382
transform 1 0 52512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_548
timestamp 1679585382
transform 1 0 53184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_555
timestamp 1679585382
transform 1 0 53856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_562
timestamp 1679585382
transform 1 0 54528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_569
timestamp 1679585382
transform 1 0 55200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_576
timestamp 1679585382
transform 1 0 55872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_583
timestamp 1679585382
transform 1 0 56544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_590
timestamp 1679585382
transform 1 0 57216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_597
timestamp 1679585382
transform 1 0 57888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_604
timestamp 1679585382
transform 1 0 58560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_611
timestamp 1679585382
transform 1 0 59232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_618
timestamp 1679585382
transform 1 0 59904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_625
timestamp 1679585382
transform 1 0 60576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_632
timestamp 1679585382
transform 1 0 61248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_639
timestamp 1679585382
transform 1 0 61920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_646
timestamp 1679585382
transform 1 0 62592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_653
timestamp 1679585382
transform 1 0 63264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_660
timestamp 1679585382
transform 1 0 63936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_667
timestamp 1679585382
transform 1 0 64608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_674
timestamp 1679585382
transform 1 0 65280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_681
timestamp 1679585382
transform 1 0 65952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_688
timestamp 1679585382
transform 1 0 66624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_695
timestamp 1679585382
transform 1 0 67296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_702
timestamp 1679585382
transform 1 0 67968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_709
timestamp 1679585382
transform 1 0 68640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_716
timestamp 1679585382
transform 1 0 69312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_723
timestamp 1679585382
transform 1 0 69984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_730
timestamp 1679585382
transform 1 0 70656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_737
timestamp 1679585382
transform 1 0 71328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_744
timestamp 1679585382
transform 1 0 72000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_751
timestamp 1679585382
transform 1 0 72672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_758
timestamp 1679585382
transform 1 0 73344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_765
timestamp 1679585382
transform 1 0 74016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_772
timestamp 1679585382
transform 1 0 74688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_779
timestamp 1679585382
transform 1 0 75360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_786
timestamp 1679585382
transform 1 0 76032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_793
timestamp 1679585382
transform 1 0 76704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_800
timestamp 1679585382
transform 1 0 77376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_807
timestamp 1679585382
transform 1 0 78048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_814
timestamp 1679585382
transform 1 0 78720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_821
timestamp 1679585382
transform 1 0 79392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_828
timestamp 1679585382
transform 1 0 80064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_835
timestamp 1679585382
transform 1 0 80736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_842
timestamp 1679585382
transform 1 0 81408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_849
timestamp 1679585382
transform 1 0 82080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_856
timestamp 1679585382
transform 1 0 82752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_863
timestamp 1679585382
transform 1 0 83424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_870
timestamp 1679585382
transform 1 0 84096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_877
timestamp 1679585382
transform 1 0 84768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_884
timestamp 1679585382
transform 1 0 85440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_891
timestamp 1679585382
transform 1 0 86112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_898
timestamp 1679585382
transform 1 0 86784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_905
timestamp 1679585382
transform 1 0 87456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_912
timestamp 1679585382
transform 1 0 88128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_919
timestamp 1679585382
transform 1 0 88800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_926
timestamp 1679585382
transform 1 0 89472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_933
timestamp 1679585382
transform 1 0 90144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_940
timestamp 1679585382
transform 1 0 90816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_947
timestamp 1679585382
transform 1 0 91488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_954
timestamp 1679585382
transform 1 0 92160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_961
timestamp 1679585382
transform 1 0 92832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_968
timestamp 1679585382
transform 1 0 93504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_975
timestamp 1679585382
transform 1 0 94176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_982
timestamp 1679585382
transform 1 0 94848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_989
timestamp 1679585382
transform 1 0 95520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_996
timestamp 1679585382
transform 1 0 96192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1003
timestamp 1679585382
transform 1 0 96864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1010
timestamp 1679585382
transform 1 0 97536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1017
timestamp 1679585382
transform 1 0 98208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_1024
timestamp 1679581501
transform 1 0 98880 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_1028
timestamp 1677583258
transform 1 0 99264 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679585382
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679585382
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679585382
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_25
timestamp 1679585382
transform 1 0 2976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_32
timestamp 1679585382
transform 1 0 3648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_39
timestamp 1679585382
transform 1 0 4320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679585382
transform 1 0 4992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679585382
transform 1 0 5664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679585382
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_67
timestamp 1679585382
transform 1 0 7008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_74
timestamp 1679585382
transform 1 0 7680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_81
timestamp 1679585382
transform 1 0 8352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679585382
transform 1 0 9024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_95
timestamp 1679585382
transform 1 0 9696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_102
timestamp 1679585382
transform 1 0 10368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_109
timestamp 1679585382
transform 1 0 11040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_116
timestamp 1679585382
transform 1 0 11712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_123
timestamp 1679585382
transform 1 0 12384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_130
timestamp 1679585382
transform 1 0 13056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_137
timestamp 1679585382
transform 1 0 13728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_144
timestamp 1679585382
transform 1 0 14400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_151
timestamp 1679585382
transform 1 0 15072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_158
timestamp 1679585382
transform 1 0 15744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_165
timestamp 1679585382
transform 1 0 16416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_172
timestamp 1679585382
transform 1 0 17088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_179
timestamp 1679585382
transform 1 0 17760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_186
timestamp 1679585382
transform 1 0 18432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_193
timestamp 1679585382
transform 1 0 19104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_200
timestamp 1679585382
transform 1 0 19776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_207
timestamp 1679585382
transform 1 0 20448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_214
timestamp 1679585382
transform 1 0 21120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_221
timestamp 1679585382
transform 1 0 21792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_228
timestamp 1679585382
transform 1 0 22464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_235
timestamp 1679585382
transform 1 0 23136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_242
timestamp 1679585382
transform 1 0 23808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_249
timestamp 1679585382
transform 1 0 24480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_256
timestamp 1679585382
transform 1 0 25152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_263
timestamp 1679585382
transform 1 0 25824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_270
timestamp 1679585382
transform 1 0 26496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_277
timestamp 1679585382
transform 1 0 27168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_284
timestamp 1679585382
transform 1 0 27840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_291
timestamp 1679585382
transform 1 0 28512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_298
timestamp 1679585382
transform 1 0 29184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_305
timestamp 1679585382
transform 1 0 29856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_312
timestamp 1679585382
transform 1 0 30528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_319
timestamp 1679585382
transform 1 0 31200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_326
timestamp 1679585382
transform 1 0 31872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_333
timestamp 1679585382
transform 1 0 32544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_340
timestamp 1679585382
transform 1 0 33216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_347
timestamp 1679585382
transform 1 0 33888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_354
timestamp 1679585382
transform 1 0 34560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_361
timestamp 1679585382
transform 1 0 35232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_368
timestamp 1679585382
transform 1 0 35904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_375
timestamp 1679585382
transform 1 0 36576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_382
timestamp 1679585382
transform 1 0 37248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_389
timestamp 1679585382
transform 1 0 37920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_396
timestamp 1679585382
transform 1 0 38592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_403
timestamp 1679585382
transform 1 0 39264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_410
timestamp 1679585382
transform 1 0 39936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_417
timestamp 1679585382
transform 1 0 40608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_424
timestamp 1679585382
transform 1 0 41280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_431
timestamp 1679585382
transform 1 0 41952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_438
timestamp 1679585382
transform 1 0 42624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_445
timestamp 1679585382
transform 1 0 43296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_452
timestamp 1679585382
transform 1 0 43968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_459
timestamp 1679585382
transform 1 0 44640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_466
timestamp 1679585382
transform 1 0 45312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_473
timestamp 1679585382
transform 1 0 45984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_480
timestamp 1679585382
transform 1 0 46656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_487
timestamp 1679585382
transform 1 0 47328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_494
timestamp 1679585382
transform 1 0 48000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_501
timestamp 1679585382
transform 1 0 48672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_508
timestamp 1679585382
transform 1 0 49344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_515
timestamp 1679585382
transform 1 0 50016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_522
timestamp 1679585382
transform 1 0 50688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_529
timestamp 1679585382
transform 1 0 51360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_536
timestamp 1679585382
transform 1 0 52032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_543
timestamp 1679585382
transform 1 0 52704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_550
timestamp 1679585382
transform 1 0 53376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_557
timestamp 1679585382
transform 1 0 54048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_564
timestamp 1679585382
transform 1 0 54720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_571
timestamp 1679585382
transform 1 0 55392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_578
timestamp 1679585382
transform 1 0 56064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_585
timestamp 1679585382
transform 1 0 56736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_592
timestamp 1679585382
transform 1 0 57408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_599
timestamp 1679585382
transform 1 0 58080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_606
timestamp 1679585382
transform 1 0 58752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_613
timestamp 1679585382
transform 1 0 59424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_620
timestamp 1679585382
transform 1 0 60096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_627
timestamp 1679585382
transform 1 0 60768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_634
timestamp 1679585382
transform 1 0 61440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_641
timestamp 1679585382
transform 1 0 62112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_648
timestamp 1679585382
transform 1 0 62784 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_655
timestamp 1679585382
transform 1 0 63456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_662
timestamp 1679585382
transform 1 0 64128 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_669
timestamp 1679585382
transform 1 0 64800 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_676
timestamp 1679585382
transform 1 0 65472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_683
timestamp 1679585382
transform 1 0 66144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_690
timestamp 1679585382
transform 1 0 66816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_697
timestamp 1679585382
transform 1 0 67488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_704
timestamp 1679585382
transform 1 0 68160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_711
timestamp 1679585382
transform 1 0 68832 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_718
timestamp 1679585382
transform 1 0 69504 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_725
timestamp 1679585382
transform 1 0 70176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_732
timestamp 1679585382
transform 1 0 70848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_739
timestamp 1679585382
transform 1 0 71520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_746
timestamp 1679585382
transform 1 0 72192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_753
timestamp 1679585382
transform 1 0 72864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_760
timestamp 1679585382
transform 1 0 73536 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_767
timestamp 1679585382
transform 1 0 74208 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_774
timestamp 1679585382
transform 1 0 74880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_781
timestamp 1679585382
transform 1 0 75552 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_788
timestamp 1679585382
transform 1 0 76224 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_795
timestamp 1679585382
transform 1 0 76896 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_802
timestamp 1679585382
transform 1 0 77568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_809
timestamp 1679585382
transform 1 0 78240 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_816
timestamp 1679585382
transform 1 0 78912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_823
timestamp 1679585382
transform 1 0 79584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_830
timestamp 1679585382
transform 1 0 80256 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_837
timestamp 1679585382
transform 1 0 80928 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_844
timestamp 1679585382
transform 1 0 81600 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_851
timestamp 1679585382
transform 1 0 82272 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_858
timestamp 1679585382
transform 1 0 82944 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_865
timestamp 1679585382
transform 1 0 83616 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_872
timestamp 1679585382
transform 1 0 84288 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_879
timestamp 1679585382
transform 1 0 84960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_886
timestamp 1679585382
transform 1 0 85632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_893
timestamp 1679585382
transform 1 0 86304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_900
timestamp 1679585382
transform 1 0 86976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_907
timestamp 1679585382
transform 1 0 87648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_914
timestamp 1679585382
transform 1 0 88320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_921
timestamp 1679585382
transform 1 0 88992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_928
timestamp 1679585382
transform 1 0 89664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_935
timestamp 1679585382
transform 1 0 90336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_942
timestamp 1679585382
transform 1 0 91008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_949
timestamp 1679585382
transform 1 0 91680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_956
timestamp 1679585382
transform 1 0 92352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_963
timestamp 1679585382
transform 1 0 93024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_970
timestamp 1679585382
transform 1 0 93696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_977
timestamp 1679585382
transform 1 0 94368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_984
timestamp 1679585382
transform 1 0 95040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_991
timestamp 1679585382
transform 1 0 95712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_998
timestamp 1679585382
transform 1 0 96384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1005
timestamp 1679585382
transform 1 0 97056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1012
timestamp 1679585382
transform 1 0 97728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1019
timestamp 1679585382
transform 1 0 98400 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_1026
timestamp 1677583704
transform 1 0 99072 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_1028
timestamp 1677583258
transform 1 0 99264 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_4
timestamp 1679585382
transform 1 0 960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_11
timestamp 1679585382
transform 1 0 1632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_18
timestamp 1679585382
transform 1 0 2304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_25
timestamp 1679585382
transform 1 0 2976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_32
timestamp 1679585382
transform 1 0 3648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_39
timestamp 1679585382
transform 1 0 4320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_46
timestamp 1679585382
transform 1 0 4992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_53
timestamp 1679585382
transform 1 0 5664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_60
timestamp 1679585382
transform 1 0 6336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_67
timestamp 1679585382
transform 1 0 7008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_74
timestamp 1679585382
transform 1 0 7680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_81
timestamp 1679585382
transform 1 0 8352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_88
timestamp 1679585382
transform 1 0 9024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_95
timestamp 1679585382
transform 1 0 9696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_102
timestamp 1679585382
transform 1 0 10368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_109
timestamp 1679585382
transform 1 0 11040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_116
timestamp 1679585382
transform 1 0 11712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_123
timestamp 1679585382
transform 1 0 12384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_130
timestamp 1679585382
transform 1 0 13056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_137
timestamp 1679585382
transform 1 0 13728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_144
timestamp 1679585382
transform 1 0 14400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_151
timestamp 1679585382
transform 1 0 15072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_158
timestamp 1679585382
transform 1 0 15744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_165
timestamp 1679585382
transform 1 0 16416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_172
timestamp 1679585382
transform 1 0 17088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_179
timestamp 1679585382
transform 1 0 17760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_186
timestamp 1679585382
transform 1 0 18432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_193
timestamp 1679585382
transform 1 0 19104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_200
timestamp 1679585382
transform 1 0 19776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_207
timestamp 1679585382
transform 1 0 20448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_214
timestamp 1679585382
transform 1 0 21120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_221
timestamp 1679585382
transform 1 0 21792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_228
timestamp 1679585382
transform 1 0 22464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_235
timestamp 1679585382
transform 1 0 23136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_242
timestamp 1679585382
transform 1 0 23808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_249
timestamp 1679585382
transform 1 0 24480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_256
timestamp 1679585382
transform 1 0 25152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_263
timestamp 1679585382
transform 1 0 25824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_270
timestamp 1679585382
transform 1 0 26496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_277
timestamp 1679585382
transform 1 0 27168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_284
timestamp 1679585382
transform 1 0 27840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_291
timestamp 1679585382
transform 1 0 28512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_298
timestamp 1679585382
transform 1 0 29184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_305
timestamp 1679585382
transform 1 0 29856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_312
timestamp 1679585382
transform 1 0 30528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_319
timestamp 1679585382
transform 1 0 31200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_326
timestamp 1679585382
transform 1 0 31872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_333
timestamp 1679585382
transform 1 0 32544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_340
timestamp 1679585382
transform 1 0 33216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_347
timestamp 1679585382
transform 1 0 33888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_354
timestamp 1679585382
transform 1 0 34560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_361
timestamp 1679585382
transform 1 0 35232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_368
timestamp 1679585382
transform 1 0 35904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_375
timestamp 1679585382
transform 1 0 36576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_382
timestamp 1679585382
transform 1 0 37248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_389
timestamp 1679585382
transform 1 0 37920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_396
timestamp 1679585382
transform 1 0 38592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_403
timestamp 1679585382
transform 1 0 39264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_410
timestamp 1679585382
transform 1 0 39936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_417
timestamp 1679585382
transform 1 0 40608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_424
timestamp 1679585382
transform 1 0 41280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_431
timestamp 1679585382
transform 1 0 41952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_438
timestamp 1679585382
transform 1 0 42624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_445
timestamp 1679585382
transform 1 0 43296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_452
timestamp 1679585382
transform 1 0 43968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_459
timestamp 1679585382
transform 1 0 44640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_466
timestamp 1679585382
transform 1 0 45312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_473
timestamp 1679585382
transform 1 0 45984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_480
timestamp 1679585382
transform 1 0 46656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_487
timestamp 1679585382
transform 1 0 47328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_494
timestamp 1679585382
transform 1 0 48000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_501
timestamp 1679585382
transform 1 0 48672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_508
timestamp 1679585382
transform 1 0 49344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_515
timestamp 1679585382
transform 1 0 50016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_522
timestamp 1679585382
transform 1 0 50688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_529
timestamp 1679585382
transform 1 0 51360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_536
timestamp 1679585382
transform 1 0 52032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_543
timestamp 1679585382
transform 1 0 52704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_550
timestamp 1679585382
transform 1 0 53376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_557
timestamp 1679585382
transform 1 0 54048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_564
timestamp 1679585382
transform 1 0 54720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_571
timestamp 1679585382
transform 1 0 55392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_578
timestamp 1679585382
transform 1 0 56064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_585
timestamp 1679585382
transform 1 0 56736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_592
timestamp 1679585382
transform 1 0 57408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_599
timestamp 1679585382
transform 1 0 58080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_606
timestamp 1679585382
transform 1 0 58752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_613
timestamp 1679585382
transform 1 0 59424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_620
timestamp 1679585382
transform 1 0 60096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_627
timestamp 1679585382
transform 1 0 60768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_634
timestamp 1679585382
transform 1 0 61440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_641
timestamp 1679585382
transform 1 0 62112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_648
timestamp 1679585382
transform 1 0 62784 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_655
timestamp 1679585382
transform 1 0 63456 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_662
timestamp 1679585382
transform 1 0 64128 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_669
timestamp 1679585382
transform 1 0 64800 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_676
timestamp 1679585382
transform 1 0 65472 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_683
timestamp 1679585382
transform 1 0 66144 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_690
timestamp 1679585382
transform 1 0 66816 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_697
timestamp 1679585382
transform 1 0 67488 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_704
timestamp 1679585382
transform 1 0 68160 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_711
timestamp 1679585382
transform 1 0 68832 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_718
timestamp 1679585382
transform 1 0 69504 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_725
timestamp 1679585382
transform 1 0 70176 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_732
timestamp 1679585382
transform 1 0 70848 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_739
timestamp 1679585382
transform 1 0 71520 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_746
timestamp 1679585382
transform 1 0 72192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_753
timestamp 1679585382
transform 1 0 72864 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_760
timestamp 1679585382
transform 1 0 73536 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_767
timestamp 1679585382
transform 1 0 74208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_774
timestamp 1679585382
transform 1 0 74880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_781
timestamp 1679585382
transform 1 0 75552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_788
timestamp 1679585382
transform 1 0 76224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_795
timestamp 1679585382
transform 1 0 76896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_802
timestamp 1679585382
transform 1 0 77568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_809
timestamp 1679585382
transform 1 0 78240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_816
timestamp 1679585382
transform 1 0 78912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_823
timestamp 1679585382
transform 1 0 79584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_830
timestamp 1679585382
transform 1 0 80256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_837
timestamp 1679585382
transform 1 0 80928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_844
timestamp 1679585382
transform 1 0 81600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_851
timestamp 1679585382
transform 1 0 82272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_858
timestamp 1679585382
transform 1 0 82944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_865
timestamp 1679585382
transform 1 0 83616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_872
timestamp 1679585382
transform 1 0 84288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_879
timestamp 1679585382
transform 1 0 84960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_886
timestamp 1679585382
transform 1 0 85632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_893
timestamp 1679585382
transform 1 0 86304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_900
timestamp 1679585382
transform 1 0 86976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_907
timestamp 1679585382
transform 1 0 87648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_914
timestamp 1679585382
transform 1 0 88320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_921
timestamp 1679585382
transform 1 0 88992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_928
timestamp 1679585382
transform 1 0 89664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_935
timestamp 1679585382
transform 1 0 90336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_942
timestamp 1679585382
transform 1 0 91008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_949
timestamp 1679585382
transform 1 0 91680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_956
timestamp 1679585382
transform 1 0 92352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_963
timestamp 1679585382
transform 1 0 93024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_970
timestamp 1679585382
transform 1 0 93696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_977
timestamp 1679585382
transform 1 0 94368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_984
timestamp 1679585382
transform 1 0 95040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_991
timestamp 1679585382
transform 1 0 95712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_998
timestamp 1679585382
transform 1 0 96384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1005
timestamp 1679585382
transform 1 0 97056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1012
timestamp 1679585382
transform 1 0 97728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1019
timestamp 1679585382
transform 1 0 98400 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_1026
timestamp 1677583704
transform 1 0 99072 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_1028
timestamp 1677583258
transform 1 0 99264 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679585382
transform 1 0 576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_7
timestamp 1679585382
transform 1 0 1248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1679585382
transform 1 0 1920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_21
timestamp 1679585382
transform 1 0 2592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_28
timestamp 1679585382
transform 1 0 3264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_35
timestamp 1679585382
transform 1 0 3936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_42
timestamp 1679585382
transform 1 0 4608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_49
timestamp 1679585382
transform 1 0 5280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_56
timestamp 1679585382
transform 1 0 5952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_63
timestamp 1679585382
transform 1 0 6624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_70
timestamp 1679585382
transform 1 0 7296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_77
timestamp 1679585382
transform 1 0 7968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_84
timestamp 1679585382
transform 1 0 8640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_91
timestamp 1679585382
transform 1 0 9312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_98
timestamp 1679585382
transform 1 0 9984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_105
timestamp 1679585382
transform 1 0 10656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_112
timestamp 1679585382
transform 1 0 11328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_119
timestamp 1679585382
transform 1 0 12000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_126
timestamp 1679585382
transform 1 0 12672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_133
timestamp 1679585382
transform 1 0 13344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_140
timestamp 1679585382
transform 1 0 14016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_147
timestamp 1679585382
transform 1 0 14688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_154
timestamp 1679585382
transform 1 0 15360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_161
timestamp 1679585382
transform 1 0 16032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_168
timestamp 1679585382
transform 1 0 16704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_175
timestamp 1679585382
transform 1 0 17376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_182
timestamp 1679585382
transform 1 0 18048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_189
timestamp 1679585382
transform 1 0 18720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_196
timestamp 1679585382
transform 1 0 19392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_203
timestamp 1679585382
transform 1 0 20064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_210
timestamp 1679585382
transform 1 0 20736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_217
timestamp 1679585382
transform 1 0 21408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_224
timestamp 1679585382
transform 1 0 22080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_231
timestamp 1679585382
transform 1 0 22752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_238
timestamp 1679585382
transform 1 0 23424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_245
timestamp 1679585382
transform 1 0 24096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_252
timestamp 1679585382
transform 1 0 24768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_259
timestamp 1679585382
transform 1 0 25440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_266
timestamp 1679585382
transform 1 0 26112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_273
timestamp 1679585382
transform 1 0 26784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_280
timestamp 1679585382
transform 1 0 27456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_287
timestamp 1679585382
transform 1 0 28128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_294
timestamp 1679585382
transform 1 0 28800 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_301
timestamp 1679585382
transform 1 0 29472 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_308
timestamp 1679585382
transform 1 0 30144 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_315
timestamp 1679585382
transform 1 0 30816 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_322
timestamp 1679585382
transform 1 0 31488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_329
timestamp 1679585382
transform 1 0 32160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_336
timestamp 1679585382
transform 1 0 32832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_343
timestamp 1679585382
transform 1 0 33504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_350
timestamp 1679585382
transform 1 0 34176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_357
timestamp 1679585382
transform 1 0 34848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_364
timestamp 1679585382
transform 1 0 35520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_371
timestamp 1679585382
transform 1 0 36192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_378
timestamp 1679585382
transform 1 0 36864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_385
timestamp 1679585382
transform 1 0 37536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_392
timestamp 1679585382
transform 1 0 38208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_399
timestamp 1679585382
transform 1 0 38880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_406
timestamp 1679585382
transform 1 0 39552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_413
timestamp 1679585382
transform 1 0 40224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_420
timestamp 1679585382
transform 1 0 40896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_427
timestamp 1679585382
transform 1 0 41568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_434
timestamp 1679585382
transform 1 0 42240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_441
timestamp 1679585382
transform 1 0 42912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_448
timestamp 1679585382
transform 1 0 43584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_455
timestamp 1679585382
transform 1 0 44256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_462
timestamp 1679585382
transform 1 0 44928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_469
timestamp 1679585382
transform 1 0 45600 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_476
timestamp 1679585382
transform 1 0 46272 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_483
timestamp 1679585382
transform 1 0 46944 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_490
timestamp 1679585382
transform 1 0 47616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_497
timestamp 1679585382
transform 1 0 48288 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_504
timestamp 1679585382
transform 1 0 48960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_511
timestamp 1679585382
transform 1 0 49632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_518
timestamp 1679585382
transform 1 0 50304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_525
timestamp 1679585382
transform 1 0 50976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_532
timestamp 1679585382
transform 1 0 51648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_539
timestamp 1679585382
transform 1 0 52320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_546
timestamp 1679585382
transform 1 0 52992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_553
timestamp 1679585382
transform 1 0 53664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_560
timestamp 1679585382
transform 1 0 54336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_567
timestamp 1679585382
transform 1 0 55008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_574
timestamp 1679585382
transform 1 0 55680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_581
timestamp 1679585382
transform 1 0 56352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_588
timestamp 1679585382
transform 1 0 57024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_595
timestamp 1679585382
transform 1 0 57696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_602
timestamp 1679585382
transform 1 0 58368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_609
timestamp 1679585382
transform 1 0 59040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_616
timestamp 1679585382
transform 1 0 59712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_623
timestamp 1679585382
transform 1 0 60384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_630
timestamp 1679585382
transform 1 0 61056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_637
timestamp 1679585382
transform 1 0 61728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_644
timestamp 1679585382
transform 1 0 62400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_651
timestamp 1679585382
transform 1 0 63072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_658
timestamp 1679585382
transform 1 0 63744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_665
timestamp 1679585382
transform 1 0 64416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_672
timestamp 1679585382
transform 1 0 65088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_679
timestamp 1679585382
transform 1 0 65760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_686
timestamp 1679585382
transform 1 0 66432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_693
timestamp 1679585382
transform 1 0 67104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_700
timestamp 1679585382
transform 1 0 67776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_707
timestamp 1679585382
transform 1 0 68448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_714
timestamp 1679585382
transform 1 0 69120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_721
timestamp 1679585382
transform 1 0 69792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_728
timestamp 1679585382
transform 1 0 70464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_735
timestamp 1679585382
transform 1 0 71136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_742
timestamp 1679585382
transform 1 0 71808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_749
timestamp 1679585382
transform 1 0 72480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_756
timestamp 1679585382
transform 1 0 73152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_763
timestamp 1679585382
transform 1 0 73824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_770
timestamp 1679585382
transform 1 0 74496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_777
timestamp 1679585382
transform 1 0 75168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_784
timestamp 1679585382
transform 1 0 75840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_791
timestamp 1679585382
transform 1 0 76512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_798
timestamp 1679585382
transform 1 0 77184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_805
timestamp 1679585382
transform 1 0 77856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_812
timestamp 1679585382
transform 1 0 78528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_819
timestamp 1679585382
transform 1 0 79200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_826
timestamp 1679585382
transform 1 0 79872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_833
timestamp 1679585382
transform 1 0 80544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_840
timestamp 1679585382
transform 1 0 81216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_847
timestamp 1679585382
transform 1 0 81888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_854
timestamp 1679585382
transform 1 0 82560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_861
timestamp 1679585382
transform 1 0 83232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_868
timestamp 1679585382
transform 1 0 83904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_875
timestamp 1679585382
transform 1 0 84576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_882
timestamp 1679585382
transform 1 0 85248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_889
timestamp 1679585382
transform 1 0 85920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_896
timestamp 1679585382
transform 1 0 86592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_903
timestamp 1679585382
transform 1 0 87264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_910
timestamp 1679585382
transform 1 0 87936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_917
timestamp 1679585382
transform 1 0 88608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_924
timestamp 1679585382
transform 1 0 89280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_931
timestamp 1679585382
transform 1 0 89952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_938
timestamp 1679585382
transform 1 0 90624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_945
timestamp 1679585382
transform 1 0 91296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_952
timestamp 1679585382
transform 1 0 91968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_959
timestamp 1679585382
transform 1 0 92640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_966
timestamp 1679585382
transform 1 0 93312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_973
timestamp 1679585382
transform 1 0 93984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_980
timestamp 1679585382
transform 1 0 94656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_987
timestamp 1679585382
transform 1 0 95328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_994
timestamp 1679585382
transform 1 0 96000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1001
timestamp 1679585382
transform 1 0 96672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1008
timestamp 1679585382
transform 1 0 97344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1015
timestamp 1679585382
transform 1 0 98016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1022
timestamp 1679585382
transform 1 0 98688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1679585382
transform 1 0 576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1679585382
transform 1 0 1248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1679585382
transform 1 0 1920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_21
timestamp 1679585382
transform 1 0 2592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_28
timestamp 1679585382
transform 1 0 3264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_35
timestamp 1679585382
transform 1 0 3936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_42
timestamp 1679585382
transform 1 0 4608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_49
timestamp 1679585382
transform 1 0 5280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_56
timestamp 1679585382
transform 1 0 5952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_63
timestamp 1679585382
transform 1 0 6624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_70
timestamp 1679585382
transform 1 0 7296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_77
timestamp 1679585382
transform 1 0 7968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_84
timestamp 1679585382
transform 1 0 8640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_91
timestamp 1679585382
transform 1 0 9312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_98
timestamp 1679585382
transform 1 0 9984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_105
timestamp 1679585382
transform 1 0 10656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_112
timestamp 1679585382
transform 1 0 11328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_119
timestamp 1679585382
transform 1 0 12000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_126
timestamp 1679585382
transform 1 0 12672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_133
timestamp 1679585382
transform 1 0 13344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_140
timestamp 1679585382
transform 1 0 14016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_147
timestamp 1679585382
transform 1 0 14688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_154
timestamp 1679585382
transform 1 0 15360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_161
timestamp 1679585382
transform 1 0 16032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_168
timestamp 1679585382
transform 1 0 16704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_175
timestamp 1679585382
transform 1 0 17376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_182
timestamp 1679585382
transform 1 0 18048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_189
timestamp 1679585382
transform 1 0 18720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_196
timestamp 1679585382
transform 1 0 19392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_203
timestamp 1679585382
transform 1 0 20064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_210
timestamp 1679585382
transform 1 0 20736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_217
timestamp 1679585382
transform 1 0 21408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_224
timestamp 1679585382
transform 1 0 22080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_231
timestamp 1679585382
transform 1 0 22752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_238
timestamp 1679585382
transform 1 0 23424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_245
timestamp 1679585382
transform 1 0 24096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_252
timestamp 1679585382
transform 1 0 24768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_259
timestamp 1679585382
transform 1 0 25440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_266
timestamp 1679585382
transform 1 0 26112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_273
timestamp 1679585382
transform 1 0 26784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_280
timestamp 1679585382
transform 1 0 27456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_287
timestamp 1679585382
transform 1 0 28128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_294
timestamp 1679585382
transform 1 0 28800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_301
timestamp 1679585382
transform 1 0 29472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_308
timestamp 1679585382
transform 1 0 30144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_315
timestamp 1679585382
transform 1 0 30816 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_322
timestamp 1679585382
transform 1 0 31488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_329
timestamp 1679585382
transform 1 0 32160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_336
timestamp 1679585382
transform 1 0 32832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_343
timestamp 1679585382
transform 1 0 33504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_350
timestamp 1679585382
transform 1 0 34176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_357
timestamp 1679585382
transform 1 0 34848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_364
timestamp 1679585382
transform 1 0 35520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_371
timestamp 1679585382
transform 1 0 36192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_378
timestamp 1679585382
transform 1 0 36864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_385
timestamp 1679585382
transform 1 0 37536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_392
timestamp 1679585382
transform 1 0 38208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_399
timestamp 1679585382
transform 1 0 38880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_406
timestamp 1679585382
transform 1 0 39552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_413
timestamp 1679585382
transform 1 0 40224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_420
timestamp 1679585382
transform 1 0 40896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_427
timestamp 1679585382
transform 1 0 41568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_434
timestamp 1679585382
transform 1 0 42240 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_441
timestamp 1679585382
transform 1 0 42912 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_448
timestamp 1679585382
transform 1 0 43584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_455
timestamp 1679585382
transform 1 0 44256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_462
timestamp 1679585382
transform 1 0 44928 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_469
timestamp 1679585382
transform 1 0 45600 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_476
timestamp 1679585382
transform 1 0 46272 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_483
timestamp 1679585382
transform 1 0 46944 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_490
timestamp 1679585382
transform 1 0 47616 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_497
timestamp 1679585382
transform 1 0 48288 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_504
timestamp 1679585382
transform 1 0 48960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_511
timestamp 1679585382
transform 1 0 49632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_518
timestamp 1679585382
transform 1 0 50304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_525
timestamp 1679585382
transform 1 0 50976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_532
timestamp 1679585382
transform 1 0 51648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_539
timestamp 1679585382
transform 1 0 52320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_546
timestamp 1679585382
transform 1 0 52992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_553
timestamp 1679585382
transform 1 0 53664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_560
timestamp 1679585382
transform 1 0 54336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_567
timestamp 1679585382
transform 1 0 55008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_574
timestamp 1679585382
transform 1 0 55680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_581
timestamp 1679585382
transform 1 0 56352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_588
timestamp 1679585382
transform 1 0 57024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_595
timestamp 1679585382
transform 1 0 57696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_602
timestamp 1679585382
transform 1 0 58368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_609
timestamp 1679585382
transform 1 0 59040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_616
timestamp 1679585382
transform 1 0 59712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_623
timestamp 1679585382
transform 1 0 60384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_630
timestamp 1679585382
transform 1 0 61056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_637
timestamp 1679585382
transform 1 0 61728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_644
timestamp 1679585382
transform 1 0 62400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_651
timestamp 1679585382
transform 1 0 63072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_658
timestamp 1679585382
transform 1 0 63744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_665
timestamp 1679585382
transform 1 0 64416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_672
timestamp 1679585382
transform 1 0 65088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_679
timestamp 1679585382
transform 1 0 65760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_686
timestamp 1679585382
transform 1 0 66432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_693
timestamp 1679585382
transform 1 0 67104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_700
timestamp 1679585382
transform 1 0 67776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_707
timestamp 1679585382
transform 1 0 68448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_714
timestamp 1679585382
transform 1 0 69120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_721
timestamp 1679585382
transform 1 0 69792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_728
timestamp 1679585382
transform 1 0 70464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_735
timestamp 1679585382
transform 1 0 71136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_742
timestamp 1679585382
transform 1 0 71808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_749
timestamp 1679585382
transform 1 0 72480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_756
timestamp 1679585382
transform 1 0 73152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_763
timestamp 1679585382
transform 1 0 73824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_770
timestamp 1679585382
transform 1 0 74496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_777
timestamp 1679585382
transform 1 0 75168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_784
timestamp 1679585382
transform 1 0 75840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_791
timestamp 1679585382
transform 1 0 76512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_798
timestamp 1679585382
transform 1 0 77184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_805
timestamp 1679585382
transform 1 0 77856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_812
timestamp 1679585382
transform 1 0 78528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_819
timestamp 1679585382
transform 1 0 79200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_826
timestamp 1679585382
transform 1 0 79872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_833
timestamp 1679585382
transform 1 0 80544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_840
timestamp 1679585382
transform 1 0 81216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_847
timestamp 1679585382
transform 1 0 81888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_854
timestamp 1679585382
transform 1 0 82560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_861
timestamp 1679585382
transform 1 0 83232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_868
timestamp 1679585382
transform 1 0 83904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_875
timestamp 1679585382
transform 1 0 84576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_882
timestamp 1679585382
transform 1 0 85248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_889
timestamp 1679585382
transform 1 0 85920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_896
timestamp 1679585382
transform 1 0 86592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_903
timestamp 1679585382
transform 1 0 87264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_910
timestamp 1679585382
transform 1 0 87936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_917
timestamp 1679585382
transform 1 0 88608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_924
timestamp 1679585382
transform 1 0 89280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_931
timestamp 1679585382
transform 1 0 89952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_938
timestamp 1679585382
transform 1 0 90624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_945
timestamp 1679585382
transform 1 0 91296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_952
timestamp 1679585382
transform 1 0 91968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_959
timestamp 1679585382
transform 1 0 92640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_966
timestamp 1679585382
transform 1 0 93312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_973
timestamp 1679585382
transform 1 0 93984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_980
timestamp 1679585382
transform 1 0 94656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_987
timestamp 1679585382
transform 1 0 95328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_994
timestamp 1679585382
transform 1 0 96000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1001
timestamp 1679585382
transform 1 0 96672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1008
timestamp 1679585382
transform 1 0 97344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1015
timestamp 1679585382
transform 1 0 98016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1022
timestamp 1679585382
transform 1 0 98688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679585382
transform 1 0 576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_7
timestamp 1679585382
transform 1 0 1248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_14
timestamp 1679585382
transform 1 0 1920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_21
timestamp 1679585382
transform 1 0 2592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_28
timestamp 1679585382
transform 1 0 3264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_35
timestamp 1679585382
transform 1 0 3936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_42
timestamp 1679585382
transform 1 0 4608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_49
timestamp 1679585382
transform 1 0 5280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_56
timestamp 1679585382
transform 1 0 5952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_63
timestamp 1679585382
transform 1 0 6624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_70
timestamp 1679585382
transform 1 0 7296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_77
timestamp 1679585382
transform 1 0 7968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_84
timestamp 1679585382
transform 1 0 8640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_91
timestamp 1679585382
transform 1 0 9312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_98
timestamp 1679585382
transform 1 0 9984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_105
timestamp 1679585382
transform 1 0 10656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_112
timestamp 1679585382
transform 1 0 11328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_119
timestamp 1679585382
transform 1 0 12000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_126
timestamp 1679585382
transform 1 0 12672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_133
timestamp 1679585382
transform 1 0 13344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_140
timestamp 1679585382
transform 1 0 14016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_147
timestamp 1679585382
transform 1 0 14688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_154
timestamp 1679585382
transform 1 0 15360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_161
timestamp 1679585382
transform 1 0 16032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_168
timestamp 1679585382
transform 1 0 16704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_175
timestamp 1679585382
transform 1 0 17376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_182
timestamp 1679585382
transform 1 0 18048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_189
timestamp 1679585382
transform 1 0 18720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_196
timestamp 1679585382
transform 1 0 19392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_203
timestamp 1679585382
transform 1 0 20064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_210
timestamp 1679585382
transform 1 0 20736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_217
timestamp 1679585382
transform 1 0 21408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_224
timestamp 1679585382
transform 1 0 22080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_231
timestamp 1679585382
transform 1 0 22752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_238
timestamp 1679585382
transform 1 0 23424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_245
timestamp 1679585382
transform 1 0 24096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_252
timestamp 1679585382
transform 1 0 24768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_259
timestamp 1679585382
transform 1 0 25440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_266
timestamp 1679585382
transform 1 0 26112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_273
timestamp 1679585382
transform 1 0 26784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_280
timestamp 1679585382
transform 1 0 27456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_287
timestamp 1679585382
transform 1 0 28128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_294
timestamp 1679585382
transform 1 0 28800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_301
timestamp 1679585382
transform 1 0 29472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_308
timestamp 1679585382
transform 1 0 30144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_315
timestamp 1679585382
transform 1 0 30816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_322
timestamp 1679585382
transform 1 0 31488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_329
timestamp 1679585382
transform 1 0 32160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_336
timestamp 1679585382
transform 1 0 32832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_343
timestamp 1679585382
transform 1 0 33504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_350
timestamp 1679585382
transform 1 0 34176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_357
timestamp 1679585382
transform 1 0 34848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_364
timestamp 1679585382
transform 1 0 35520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_371
timestamp 1679585382
transform 1 0 36192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_378
timestamp 1679585382
transform 1 0 36864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_385
timestamp 1679585382
transform 1 0 37536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_392
timestamp 1679585382
transform 1 0 38208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_399
timestamp 1679585382
transform 1 0 38880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_406
timestamp 1679585382
transform 1 0 39552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_413
timestamp 1679585382
transform 1 0 40224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_420
timestamp 1679585382
transform 1 0 40896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_427
timestamp 1679585382
transform 1 0 41568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_434
timestamp 1679585382
transform 1 0 42240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_441
timestamp 1679585382
transform 1 0 42912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_448
timestamp 1679585382
transform 1 0 43584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_455
timestamp 1679585382
transform 1 0 44256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_462
timestamp 1679585382
transform 1 0 44928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_469
timestamp 1679585382
transform 1 0 45600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_476
timestamp 1679585382
transform 1 0 46272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_483
timestamp 1679585382
transform 1 0 46944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_490
timestamp 1679585382
transform 1 0 47616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_497
timestamp 1679585382
transform 1 0 48288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_504
timestamp 1679585382
transform 1 0 48960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_511
timestamp 1679585382
transform 1 0 49632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_518
timestamp 1679585382
transform 1 0 50304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_525
timestamp 1679585382
transform 1 0 50976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_532
timestamp 1679585382
transform 1 0 51648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_539
timestamp 1679585382
transform 1 0 52320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_546
timestamp 1679585382
transform 1 0 52992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_553
timestamp 1679585382
transform 1 0 53664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_560
timestamp 1679585382
transform 1 0 54336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_567
timestamp 1679585382
transform 1 0 55008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_574
timestamp 1679585382
transform 1 0 55680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_581
timestamp 1679585382
transform 1 0 56352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_588
timestamp 1679585382
transform 1 0 57024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_595
timestamp 1679585382
transform 1 0 57696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_602
timestamp 1679585382
transform 1 0 58368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_609
timestamp 1679585382
transform 1 0 59040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_616
timestamp 1679585382
transform 1 0 59712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_623
timestamp 1679585382
transform 1 0 60384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_630
timestamp 1679585382
transform 1 0 61056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_637
timestamp 1679585382
transform 1 0 61728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_644
timestamp 1679585382
transform 1 0 62400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_651
timestamp 1679585382
transform 1 0 63072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_658
timestamp 1679585382
transform 1 0 63744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_665
timestamp 1679585382
transform 1 0 64416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_672
timestamp 1679585382
transform 1 0 65088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_679
timestamp 1679585382
transform 1 0 65760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_686
timestamp 1679585382
transform 1 0 66432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_693
timestamp 1679585382
transform 1 0 67104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_700
timestamp 1679585382
transform 1 0 67776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_707
timestamp 1679585382
transform 1 0 68448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_714
timestamp 1679585382
transform 1 0 69120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_721
timestamp 1679585382
transform 1 0 69792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_728
timestamp 1679585382
transform 1 0 70464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_735
timestamp 1679585382
transform 1 0 71136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_742
timestamp 1679585382
transform 1 0 71808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_749
timestamp 1679585382
transform 1 0 72480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_756
timestamp 1679585382
transform 1 0 73152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_763
timestamp 1679585382
transform 1 0 73824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_770
timestamp 1679585382
transform 1 0 74496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_777
timestamp 1679585382
transform 1 0 75168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_784
timestamp 1679585382
transform 1 0 75840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_791
timestamp 1679585382
transform 1 0 76512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_798
timestamp 1679585382
transform 1 0 77184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_805
timestamp 1679585382
transform 1 0 77856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_812
timestamp 1679585382
transform 1 0 78528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_819
timestamp 1679585382
transform 1 0 79200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_826
timestamp 1679585382
transform 1 0 79872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_833
timestamp 1679585382
transform 1 0 80544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_840
timestamp 1679585382
transform 1 0 81216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_847
timestamp 1679585382
transform 1 0 81888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_854
timestamp 1679585382
transform 1 0 82560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_861
timestamp 1679585382
transform 1 0 83232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_868
timestamp 1679585382
transform 1 0 83904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_875
timestamp 1679585382
transform 1 0 84576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_882
timestamp 1679585382
transform 1 0 85248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_889
timestamp 1679585382
transform 1 0 85920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_896
timestamp 1679585382
transform 1 0 86592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_903
timestamp 1679585382
transform 1 0 87264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_910
timestamp 1679585382
transform 1 0 87936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_917
timestamp 1679585382
transform 1 0 88608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_924
timestamp 1679585382
transform 1 0 89280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_931
timestamp 1679585382
transform 1 0 89952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_938
timestamp 1679585382
transform 1 0 90624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_945
timestamp 1679585382
transform 1 0 91296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_952
timestamp 1679585382
transform 1 0 91968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_959
timestamp 1679585382
transform 1 0 92640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_966
timestamp 1679585382
transform 1 0 93312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_973
timestamp 1679585382
transform 1 0 93984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_980
timestamp 1679585382
transform 1 0 94656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_987
timestamp 1679585382
transform 1 0 95328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_994
timestamp 1679585382
transform 1 0 96000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1001
timestamp 1679585382
transform 1 0 96672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1008
timestamp 1679585382
transform 1 0 97344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1015
timestamp 1679585382
transform 1 0 98016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1022
timestamp 1679585382
transform 1 0 98688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679585382
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679585382
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679585382
transform 1 0 1920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679585382
transform 1 0 2592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_28
timestamp 1679585382
transform 1 0 3264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_35
timestamp 1679585382
transform 1 0 3936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_42
timestamp 1679585382
transform 1 0 4608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_49
timestamp 1679585382
transform 1 0 5280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_56
timestamp 1679585382
transform 1 0 5952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_63
timestamp 1679585382
transform 1 0 6624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_70
timestamp 1679585382
transform 1 0 7296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_77
timestamp 1679585382
transform 1 0 7968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_84
timestamp 1679585382
transform 1 0 8640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_91
timestamp 1679585382
transform 1 0 9312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_98
timestamp 1679585382
transform 1 0 9984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_105
timestamp 1679585382
transform 1 0 10656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_112
timestamp 1679585382
transform 1 0 11328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_119
timestamp 1679585382
transform 1 0 12000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_126
timestamp 1679585382
transform 1 0 12672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_133
timestamp 1679585382
transform 1 0 13344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_140
timestamp 1679585382
transform 1 0 14016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_147
timestamp 1679585382
transform 1 0 14688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_154
timestamp 1679585382
transform 1 0 15360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_161
timestamp 1679585382
transform 1 0 16032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_168
timestamp 1679585382
transform 1 0 16704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_175
timestamp 1679585382
transform 1 0 17376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_182
timestamp 1679585382
transform 1 0 18048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_189
timestamp 1679585382
transform 1 0 18720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_196
timestamp 1679585382
transform 1 0 19392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_203
timestamp 1679585382
transform 1 0 20064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_210
timestamp 1679585382
transform 1 0 20736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_217
timestamp 1679585382
transform 1 0 21408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_224
timestamp 1679585382
transform 1 0 22080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_231
timestamp 1679585382
transform 1 0 22752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_238
timestamp 1679585382
transform 1 0 23424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_245
timestamp 1679585382
transform 1 0 24096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_252
timestamp 1679585382
transform 1 0 24768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_259
timestamp 1679585382
transform 1 0 25440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_266
timestamp 1679585382
transform 1 0 26112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_273
timestamp 1679585382
transform 1 0 26784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_280
timestamp 1679585382
transform 1 0 27456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_287
timestamp 1679585382
transform 1 0 28128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_294
timestamp 1679585382
transform 1 0 28800 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_301
timestamp 1679585382
transform 1 0 29472 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_308
timestamp 1679585382
transform 1 0 30144 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_315
timestamp 1679585382
transform 1 0 30816 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_322
timestamp 1679585382
transform 1 0 31488 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_329
timestamp 1679585382
transform 1 0 32160 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_336
timestamp 1679585382
transform 1 0 32832 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_343
timestamp 1679585382
transform 1 0 33504 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_350
timestamp 1679585382
transform 1 0 34176 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_357
timestamp 1679585382
transform 1 0 34848 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_364
timestamp 1679585382
transform 1 0 35520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_371
timestamp 1679585382
transform 1 0 36192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_378
timestamp 1679585382
transform 1 0 36864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_385
timestamp 1679585382
transform 1 0 37536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_392
timestamp 1679585382
transform 1 0 38208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_399
timestamp 1679585382
transform 1 0 38880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_406
timestamp 1679585382
transform 1 0 39552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_413
timestamp 1679585382
transform 1 0 40224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_420
timestamp 1679585382
transform 1 0 40896 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_427
timestamp 1679585382
transform 1 0 41568 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_434
timestamp 1679585382
transform 1 0 42240 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_441
timestamp 1679585382
transform 1 0 42912 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_448
timestamp 1679585382
transform 1 0 43584 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_455
timestamp 1679585382
transform 1 0 44256 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_462
timestamp 1679585382
transform 1 0 44928 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_469
timestamp 1679585382
transform 1 0 45600 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_476
timestamp 1679585382
transform 1 0 46272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_483
timestamp 1679585382
transform 1 0 46944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_490
timestamp 1679585382
transform 1 0 47616 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_497
timestamp 1679585382
transform 1 0 48288 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_504
timestamp 1679585382
transform 1 0 48960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_511
timestamp 1679585382
transform 1 0 49632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_518
timestamp 1679585382
transform 1 0 50304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_525
timestamp 1679585382
transform 1 0 50976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_532
timestamp 1679585382
transform 1 0 51648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_539
timestamp 1679585382
transform 1 0 52320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_546
timestamp 1679585382
transform 1 0 52992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_553
timestamp 1679585382
transform 1 0 53664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_560
timestamp 1679585382
transform 1 0 54336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_567
timestamp 1679585382
transform 1 0 55008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_574
timestamp 1679585382
transform 1 0 55680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_581
timestamp 1679585382
transform 1 0 56352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_588
timestamp 1679585382
transform 1 0 57024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_595
timestamp 1679585382
transform 1 0 57696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_602
timestamp 1679585382
transform 1 0 58368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_609
timestamp 1679585382
transform 1 0 59040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_616
timestamp 1679585382
transform 1 0 59712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_623
timestamp 1679585382
transform 1 0 60384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_630
timestamp 1679585382
transform 1 0 61056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_637
timestamp 1679585382
transform 1 0 61728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_644
timestamp 1679585382
transform 1 0 62400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_651
timestamp 1679585382
transform 1 0 63072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_658
timestamp 1679585382
transform 1 0 63744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_665
timestamp 1679585382
transform 1 0 64416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_672
timestamp 1679585382
transform 1 0 65088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_679
timestamp 1679585382
transform 1 0 65760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_686
timestamp 1679585382
transform 1 0 66432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_693
timestamp 1679585382
transform 1 0 67104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_700
timestamp 1679585382
transform 1 0 67776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_707
timestamp 1679585382
transform 1 0 68448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_714
timestamp 1679585382
transform 1 0 69120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_721
timestamp 1679585382
transform 1 0 69792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_728
timestamp 1679585382
transform 1 0 70464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_735
timestamp 1679585382
transform 1 0 71136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_742
timestamp 1679585382
transform 1 0 71808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_749
timestamp 1679585382
transform 1 0 72480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_756
timestamp 1679585382
transform 1 0 73152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_763
timestamp 1679585382
transform 1 0 73824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_770
timestamp 1679585382
transform 1 0 74496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_777
timestamp 1679585382
transform 1 0 75168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_784
timestamp 1679585382
transform 1 0 75840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_791
timestamp 1679585382
transform 1 0 76512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_798
timestamp 1679585382
transform 1 0 77184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_805
timestamp 1679585382
transform 1 0 77856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_812
timestamp 1679585382
transform 1 0 78528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_819
timestamp 1679585382
transform 1 0 79200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_826
timestamp 1679585382
transform 1 0 79872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_833
timestamp 1679585382
transform 1 0 80544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_840
timestamp 1679585382
transform 1 0 81216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_847
timestamp 1679585382
transform 1 0 81888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_854
timestamp 1679585382
transform 1 0 82560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_861
timestamp 1679585382
transform 1 0 83232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_868
timestamp 1679585382
transform 1 0 83904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_875
timestamp 1679585382
transform 1 0 84576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_882
timestamp 1679585382
transform 1 0 85248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_889
timestamp 1679585382
transform 1 0 85920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_896
timestamp 1679585382
transform 1 0 86592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_903
timestamp 1679585382
transform 1 0 87264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_910
timestamp 1679585382
transform 1 0 87936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_917
timestamp 1679585382
transform 1 0 88608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_924
timestamp 1679585382
transform 1 0 89280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_931
timestamp 1679585382
transform 1 0 89952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_938
timestamp 1679585382
transform 1 0 90624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_945
timestamp 1679585382
transform 1 0 91296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_952
timestamp 1679585382
transform 1 0 91968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_959
timestamp 1679585382
transform 1 0 92640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_966
timestamp 1679585382
transform 1 0 93312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_973
timestamp 1679585382
transform 1 0 93984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_980
timestamp 1679585382
transform 1 0 94656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_987
timestamp 1679585382
transform 1 0 95328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_994
timestamp 1679585382
transform 1 0 96000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1001
timestamp 1679585382
transform 1 0 96672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1008
timestamp 1679585382
transform 1 0 97344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1015
timestamp 1679585382
transform 1 0 98016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1022
timestamp 1679585382
transform 1 0 98688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679585382
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679585382
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679585382
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679585382
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679585382
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679585382
transform 1 0 3936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679585382
transform 1 0 4608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679585382
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679585382
transform 1 0 5952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679585382
transform 1 0 6624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679585382
transform 1 0 7296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679585382
transform 1 0 7968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679585382
transform 1 0 8640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679585382
transform 1 0 9312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679585382
transform 1 0 9984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_105
timestamp 1679585382
transform 1 0 10656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679585382
transform 1 0 11328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679585382
transform 1 0 12000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679585382
transform 1 0 12672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679585382
transform 1 0 13344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679585382
transform 1 0 14016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679585382
transform 1 0 14688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679585382
transform 1 0 15360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679585382
transform 1 0 16032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679585382
transform 1 0 16704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679585382
transform 1 0 17376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679585382
transform 1 0 18048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679585382
transform 1 0 18720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679585382
transform 1 0 19392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679585382
transform 1 0 20064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679585382
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679585382
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679585382
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679585382
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679585382
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679585382
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679585382
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679585382
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679585382
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679585382
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679585382
transform 1 0 27456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679585382
transform 1 0 28128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_294
timestamp 1679585382
transform 1 0 28800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_301
timestamp 1679585382
transform 1 0 29472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_308
timestamp 1679585382
transform 1 0 30144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_315
timestamp 1679585382
transform 1 0 30816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_322
timestamp 1679585382
transform 1 0 31488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_329
timestamp 1679585382
transform 1 0 32160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_336
timestamp 1679585382
transform 1 0 32832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_343
timestamp 1679585382
transform 1 0 33504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_350
timestamp 1679585382
transform 1 0 34176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_357
timestamp 1679585382
transform 1 0 34848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_364
timestamp 1679585382
transform 1 0 35520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_371
timestamp 1679585382
transform 1 0 36192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_378
timestamp 1679585382
transform 1 0 36864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_385
timestamp 1679585382
transform 1 0 37536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_392
timestamp 1679585382
transform 1 0 38208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_399
timestamp 1679585382
transform 1 0 38880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_406
timestamp 1679585382
transform 1 0 39552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_413
timestamp 1679585382
transform 1 0 40224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_420
timestamp 1679585382
transform 1 0 40896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_427
timestamp 1679585382
transform 1 0 41568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_434
timestamp 1679585382
transform 1 0 42240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_441
timestamp 1679585382
transform 1 0 42912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_448
timestamp 1679585382
transform 1 0 43584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_455
timestamp 1679585382
transform 1 0 44256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_462
timestamp 1679585382
transform 1 0 44928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_469
timestamp 1679585382
transform 1 0 45600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_476
timestamp 1679585382
transform 1 0 46272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_483
timestamp 1679585382
transform 1 0 46944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_490
timestamp 1679585382
transform 1 0 47616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_497
timestamp 1679585382
transform 1 0 48288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_504
timestamp 1679585382
transform 1 0 48960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_511
timestamp 1679585382
transform 1 0 49632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_518
timestamp 1679585382
transform 1 0 50304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_525
timestamp 1679585382
transform 1 0 50976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_532
timestamp 1679585382
transform 1 0 51648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_539
timestamp 1679585382
transform 1 0 52320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_546
timestamp 1679585382
transform 1 0 52992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_553
timestamp 1679585382
transform 1 0 53664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_560
timestamp 1679585382
transform 1 0 54336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_567
timestamp 1679585382
transform 1 0 55008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_574
timestamp 1679585382
transform 1 0 55680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_581
timestamp 1679585382
transform 1 0 56352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_588
timestamp 1679585382
transform 1 0 57024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_595
timestamp 1679585382
transform 1 0 57696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_602
timestamp 1679585382
transform 1 0 58368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_609
timestamp 1679585382
transform 1 0 59040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_616
timestamp 1679585382
transform 1 0 59712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_623
timestamp 1679585382
transform 1 0 60384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_630
timestamp 1679585382
transform 1 0 61056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_637
timestamp 1679585382
transform 1 0 61728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_644
timestamp 1679585382
transform 1 0 62400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_651
timestamp 1679585382
transform 1 0 63072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_658
timestamp 1679585382
transform 1 0 63744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_665
timestamp 1679585382
transform 1 0 64416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_672
timestamp 1679585382
transform 1 0 65088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_679
timestamp 1679585382
transform 1 0 65760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_686
timestamp 1679585382
transform 1 0 66432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_693
timestamp 1679585382
transform 1 0 67104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_700
timestamp 1679585382
transform 1 0 67776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_707
timestamp 1679585382
transform 1 0 68448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_714
timestamp 1679585382
transform 1 0 69120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_721
timestamp 1679585382
transform 1 0 69792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_728
timestamp 1679585382
transform 1 0 70464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_735
timestamp 1679585382
transform 1 0 71136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_742
timestamp 1679585382
transform 1 0 71808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_749
timestamp 1679585382
transform 1 0 72480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_756
timestamp 1679585382
transform 1 0 73152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_763
timestamp 1679585382
transform 1 0 73824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_770
timestamp 1679585382
transform 1 0 74496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_777
timestamp 1679585382
transform 1 0 75168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_784
timestamp 1679585382
transform 1 0 75840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_791
timestamp 1679585382
transform 1 0 76512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_798
timestamp 1679585382
transform 1 0 77184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_805
timestamp 1679585382
transform 1 0 77856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_812
timestamp 1679585382
transform 1 0 78528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_819
timestamp 1679585382
transform 1 0 79200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_826
timestamp 1679585382
transform 1 0 79872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_833
timestamp 1679585382
transform 1 0 80544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_840
timestamp 1679585382
transform 1 0 81216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_847
timestamp 1679585382
transform 1 0 81888 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_854
timestamp 1679585382
transform 1 0 82560 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_861
timestamp 1679585382
transform 1 0 83232 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_868
timestamp 1679585382
transform 1 0 83904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_875
timestamp 1679585382
transform 1 0 84576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_882
timestamp 1679585382
transform 1 0 85248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_889
timestamp 1679585382
transform 1 0 85920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_896
timestamp 1679585382
transform 1 0 86592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_903
timestamp 1679585382
transform 1 0 87264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_910
timestamp 1679585382
transform 1 0 87936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_917
timestamp 1679585382
transform 1 0 88608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_924
timestamp 1679585382
transform 1 0 89280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_931
timestamp 1679585382
transform 1 0 89952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_938
timestamp 1679585382
transform 1 0 90624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_945
timestamp 1679585382
transform 1 0 91296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_952
timestamp 1679585382
transform 1 0 91968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_959
timestamp 1679585382
transform 1 0 92640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_966
timestamp 1679585382
transform 1 0 93312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_973
timestamp 1679585382
transform 1 0 93984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_980
timestamp 1679585382
transform 1 0 94656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_987
timestamp 1679585382
transform 1 0 95328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_994
timestamp 1679585382
transform 1 0 96000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1001
timestamp 1679585382
transform 1 0 96672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1008
timestamp 1679585382
transform 1 0 97344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1015
timestamp 1679585382
transform 1 0 98016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1022
timestamp 1679585382
transform 1 0 98688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679585382
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679585382
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679585382
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679585382
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679585382
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679585382
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679585382
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679585382
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679585382
transform 1 0 5952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679585382
transform 1 0 6624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679585382
transform 1 0 7296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679585382
transform 1 0 7968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679585382
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679585382
transform 1 0 9312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679585382
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679585382
transform 1 0 10656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679585382
transform 1 0 11328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679585382
transform 1 0 12000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679585382
transform 1 0 12672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679585382
transform 1 0 13344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679585382
transform 1 0 14016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679585382
transform 1 0 14688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679585382
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679585382
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679585382
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679585382
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679585382
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679585382
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679585382
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679585382
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679585382
transform 1 0 20736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679585382
transform 1 0 21408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679585382
transform 1 0 22080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679585382
transform 1 0 22752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679585382
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679585382
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679585382
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679585382
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679585382
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679585382
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679585382
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679585382
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679585382
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679585382
transform 1 0 29472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679585382
transform 1 0 30144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679585382
transform 1 0 30816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679585382
transform 1 0 31488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679585382
transform 1 0 32160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679585382
transform 1 0 32832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679585382
transform 1 0 33504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679585382
transform 1 0 34176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679585382
transform 1 0 34848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679585382
transform 1 0 35520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679585382
transform 1 0 36192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679585382
transform 1 0 36864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_385
timestamp 1679585382
transform 1 0 37536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_392
timestamp 1679585382
transform 1 0 38208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_399
timestamp 1679585382
transform 1 0 38880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_406
timestamp 1679585382
transform 1 0 39552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_413
timestamp 1679585382
transform 1 0 40224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_420
timestamp 1679585382
transform 1 0 40896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_427
timestamp 1679585382
transform 1 0 41568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_434
timestamp 1679585382
transform 1 0 42240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_441
timestamp 1679585382
transform 1 0 42912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_448
timestamp 1679585382
transform 1 0 43584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_455
timestamp 1679585382
transform 1 0 44256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_462
timestamp 1679585382
transform 1 0 44928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_469
timestamp 1679585382
transform 1 0 45600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_476
timestamp 1679585382
transform 1 0 46272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_483
timestamp 1679585382
transform 1 0 46944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_490
timestamp 1679585382
transform 1 0 47616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_497
timestamp 1679585382
transform 1 0 48288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_504
timestamp 1679585382
transform 1 0 48960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_511
timestamp 1679585382
transform 1 0 49632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_518
timestamp 1679585382
transform 1 0 50304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_525
timestamp 1679585382
transform 1 0 50976 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_532
timestamp 1679585382
transform 1 0 51648 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_539
timestamp 1679585382
transform 1 0 52320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_546
timestamp 1679585382
transform 1 0 52992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_553
timestamp 1679585382
transform 1 0 53664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_560
timestamp 1679585382
transform 1 0 54336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_567
timestamp 1679585382
transform 1 0 55008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_574
timestamp 1679585382
transform 1 0 55680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_581
timestamp 1679585382
transform 1 0 56352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_588
timestamp 1679585382
transform 1 0 57024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_595
timestamp 1679585382
transform 1 0 57696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_602
timestamp 1679585382
transform 1 0 58368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_609
timestamp 1679585382
transform 1 0 59040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_616
timestamp 1679585382
transform 1 0 59712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_623
timestamp 1679585382
transform 1 0 60384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_630
timestamp 1679585382
transform 1 0 61056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_637
timestamp 1679585382
transform 1 0 61728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_644
timestamp 1679585382
transform 1 0 62400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_651
timestamp 1679585382
transform 1 0 63072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_658
timestamp 1679585382
transform 1 0 63744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_665
timestamp 1679585382
transform 1 0 64416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_672
timestamp 1679585382
transform 1 0 65088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_679
timestamp 1679585382
transform 1 0 65760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_686
timestamp 1679585382
transform 1 0 66432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_693
timestamp 1679585382
transform 1 0 67104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_700
timestamp 1679585382
transform 1 0 67776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_707
timestamp 1679585382
transform 1 0 68448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_714
timestamp 1679585382
transform 1 0 69120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_721
timestamp 1679585382
transform 1 0 69792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_728
timestamp 1679585382
transform 1 0 70464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_735
timestamp 1679585382
transform 1 0 71136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_742
timestamp 1679585382
transform 1 0 71808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_749
timestamp 1679585382
transform 1 0 72480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_756
timestamp 1679585382
transform 1 0 73152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_763
timestamp 1679585382
transform 1 0 73824 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_770
timestamp 1679585382
transform 1 0 74496 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_777
timestamp 1679585382
transform 1 0 75168 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_784
timestamp 1679585382
transform 1 0 75840 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_791
timestamp 1679585382
transform 1 0 76512 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_798
timestamp 1679585382
transform 1 0 77184 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_805
timestamp 1679585382
transform 1 0 77856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_812
timestamp 1679585382
transform 1 0 78528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_819
timestamp 1679585382
transform 1 0 79200 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_826
timestamp 1679585382
transform 1 0 79872 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_833
timestamp 1679585382
transform 1 0 80544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_840
timestamp 1679585382
transform 1 0 81216 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_847
timestamp 1679585382
transform 1 0 81888 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_854
timestamp 1679585382
transform 1 0 82560 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_861
timestamp 1679585382
transform 1 0 83232 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_868
timestamp 1679585382
transform 1 0 83904 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_875
timestamp 1679585382
transform 1 0 84576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_882
timestamp 1679585382
transform 1 0 85248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_889
timestamp 1679585382
transform 1 0 85920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_896
timestamp 1679585382
transform 1 0 86592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_903
timestamp 1679585382
transform 1 0 87264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_910
timestamp 1679585382
transform 1 0 87936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_917
timestamp 1679585382
transform 1 0 88608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_924
timestamp 1679585382
transform 1 0 89280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_931
timestamp 1679585382
transform 1 0 89952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_938
timestamp 1679585382
transform 1 0 90624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_945
timestamp 1679585382
transform 1 0 91296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_952
timestamp 1679585382
transform 1 0 91968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_959
timestamp 1679585382
transform 1 0 92640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_966
timestamp 1679585382
transform 1 0 93312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_973
timestamp 1679585382
transform 1 0 93984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_980
timestamp 1679585382
transform 1 0 94656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_987
timestamp 1679585382
transform 1 0 95328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_994
timestamp 1679585382
transform 1 0 96000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1001
timestamp 1679585382
transform 1 0 96672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1008
timestamp 1679585382
transform 1 0 97344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1015
timestamp 1679585382
transform 1 0 98016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1022
timestamp 1679585382
transform 1 0 98688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679585382
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679585382
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679585382
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679585382
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679585382
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679585382
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679585382
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679585382
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679585382
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679585382
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679585382
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679585382
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679585382
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679585382
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679585382
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679585382
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679585382
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679585382
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679585382
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679585382
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679585382
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679585382
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679585382
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679585382
transform 1 0 16032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679585382
transform 1 0 16704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679585382
transform 1 0 17376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679585382
transform 1 0 18048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679585382
transform 1 0 18720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679585382
transform 1 0 19392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679585382
transform 1 0 20064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679585382
transform 1 0 20736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679585382
transform 1 0 21408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679585382
transform 1 0 22080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679585382
transform 1 0 22752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679585382
transform 1 0 23424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679585382
transform 1 0 24096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679585382
transform 1 0 24768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679585382
transform 1 0 25440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679585382
transform 1 0 26112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679585382
transform 1 0 26784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679585382
transform 1 0 27456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679585382
transform 1 0 28128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679585382
transform 1 0 28800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679585382
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679585382
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679585382
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679585382
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679585382
transform 1 0 32160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679585382
transform 1 0 32832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679585382
transform 1 0 33504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679585382
transform 1 0 34176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679585382
transform 1 0 34848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679585382
transform 1 0 35520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679585382
transform 1 0 36192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679585382
transform 1 0 36864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679585382
transform 1 0 37536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679585382
transform 1 0 38208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_399
timestamp 1679585382
transform 1 0 38880 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_406
timestamp 1679585382
transform 1 0 39552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_413
timestamp 1679585382
transform 1 0 40224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_420
timestamp 1679585382
transform 1 0 40896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_427
timestamp 1679585382
transform 1 0 41568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_434
timestamp 1679585382
transform 1 0 42240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_441
timestamp 1679585382
transform 1 0 42912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_448
timestamp 1679585382
transform 1 0 43584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_455
timestamp 1679585382
transform 1 0 44256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_462
timestamp 1679585382
transform 1 0 44928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_469
timestamp 1679585382
transform 1 0 45600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_476
timestamp 1679585382
transform 1 0 46272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_483
timestamp 1679585382
transform 1 0 46944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_490
timestamp 1679585382
transform 1 0 47616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_497
timestamp 1679585382
transform 1 0 48288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_504
timestamp 1679585382
transform 1 0 48960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_511
timestamp 1679585382
transform 1 0 49632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_518
timestamp 1679585382
transform 1 0 50304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_525
timestamp 1679585382
transform 1 0 50976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_532
timestamp 1679585382
transform 1 0 51648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_539
timestamp 1679585382
transform 1 0 52320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_546
timestamp 1679585382
transform 1 0 52992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_553
timestamp 1679585382
transform 1 0 53664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_560
timestamp 1679585382
transform 1 0 54336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_567
timestamp 1679585382
transform 1 0 55008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_574
timestamp 1679585382
transform 1 0 55680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_581
timestamp 1679585382
transform 1 0 56352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_588
timestamp 1679585382
transform 1 0 57024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_595
timestamp 1679585382
transform 1 0 57696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_602
timestamp 1679585382
transform 1 0 58368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_609
timestamp 1679585382
transform 1 0 59040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_616
timestamp 1679585382
transform 1 0 59712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_623
timestamp 1679585382
transform 1 0 60384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_630
timestamp 1679585382
transform 1 0 61056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_637
timestamp 1679585382
transform 1 0 61728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_644
timestamp 1679585382
transform 1 0 62400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_651
timestamp 1679585382
transform 1 0 63072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_658
timestamp 1679585382
transform 1 0 63744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_665
timestamp 1679585382
transform 1 0 64416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_672
timestamp 1679585382
transform 1 0 65088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_679
timestamp 1679585382
transform 1 0 65760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_686
timestamp 1679585382
transform 1 0 66432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_693
timestamp 1679585382
transform 1 0 67104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_700
timestamp 1679585382
transform 1 0 67776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_707
timestamp 1679585382
transform 1 0 68448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_714
timestamp 1679585382
transform 1 0 69120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_721
timestamp 1679585382
transform 1 0 69792 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_728
timestamp 1679585382
transform 1 0 70464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_735
timestamp 1679585382
transform 1 0 71136 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_742
timestamp 1679585382
transform 1 0 71808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_749
timestamp 1679585382
transform 1 0 72480 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_756
timestamp 1679585382
transform 1 0 73152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_763
timestamp 1679585382
transform 1 0 73824 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_770
timestamp 1679585382
transform 1 0 74496 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_777
timestamp 1679585382
transform 1 0 75168 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_784
timestamp 1679585382
transform 1 0 75840 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_791
timestamp 1679585382
transform 1 0 76512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_798
timestamp 1679585382
transform 1 0 77184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_805
timestamp 1679585382
transform 1 0 77856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_812
timestamp 1679585382
transform 1 0 78528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_819
timestamp 1679585382
transform 1 0 79200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_826
timestamp 1679585382
transform 1 0 79872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_833
timestamp 1679585382
transform 1 0 80544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_840
timestamp 1679585382
transform 1 0 81216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_847
timestamp 1679585382
transform 1 0 81888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_854
timestamp 1679585382
transform 1 0 82560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_861
timestamp 1679585382
transform 1 0 83232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_868
timestamp 1679585382
transform 1 0 83904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_875
timestamp 1679585382
transform 1 0 84576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_882
timestamp 1679585382
transform 1 0 85248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_889
timestamp 1679585382
transform 1 0 85920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_896
timestamp 1679585382
transform 1 0 86592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_903
timestamp 1679585382
transform 1 0 87264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_910
timestamp 1679585382
transform 1 0 87936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_917
timestamp 1679585382
transform 1 0 88608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_924
timestamp 1679585382
transform 1 0 89280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_931
timestamp 1679585382
transform 1 0 89952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_938
timestamp 1679585382
transform 1 0 90624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_945
timestamp 1679585382
transform 1 0 91296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_952
timestamp 1679585382
transform 1 0 91968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_959
timestamp 1679585382
transform 1 0 92640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_966
timestamp 1679585382
transform 1 0 93312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_973
timestamp 1679585382
transform 1 0 93984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_980
timestamp 1679585382
transform 1 0 94656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_987
timestamp 1679585382
transform 1 0 95328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_994
timestamp 1679585382
transform 1 0 96000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1001
timestamp 1679585382
transform 1 0 96672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1008
timestamp 1679585382
transform 1 0 97344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1015
timestamp 1679585382
transform 1 0 98016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1022
timestamp 1679585382
transform 1 0 98688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679585382
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679585382
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679585382
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679585382
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679585382
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679585382
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679585382
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679585382
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679585382
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679585382
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679585382
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679585382
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679585382
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679585382
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679585382
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679585382
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679585382
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679585382
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679585382
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679585382
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679585382
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679585382
transform 1 0 14688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679585382
transform 1 0 15360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679585382
transform 1 0 16032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679585382
transform 1 0 16704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679585382
transform 1 0 17376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679585382
transform 1 0 18048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679585382
transform 1 0 18720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679585382
transform 1 0 19392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679585382
transform 1 0 20064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679585382
transform 1 0 20736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679585382
transform 1 0 21408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679585382
transform 1 0 22080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679585382
transform 1 0 22752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679585382
transform 1 0 23424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679585382
transform 1 0 24096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679585382
transform 1 0 24768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679585382
transform 1 0 25440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679585382
transform 1 0 26112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679585382
transform 1 0 26784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679585382
transform 1 0 27456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679585382
transform 1 0 28128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679585382
transform 1 0 28800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679585382
transform 1 0 29472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679585382
transform 1 0 30144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679585382
transform 1 0 30816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679585382
transform 1 0 31488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679585382
transform 1 0 32160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679585382
transform 1 0 32832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679585382
transform 1 0 33504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679585382
transform 1 0 34176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679585382
transform 1 0 34848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679585382
transform 1 0 35520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679585382
transform 1 0 36192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679585382
transform 1 0 36864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679585382
transform 1 0 37536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679585382
transform 1 0 38208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_399
timestamp 1679585382
transform 1 0 38880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_406
timestamp 1679585382
transform 1 0 39552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_413
timestamp 1679585382
transform 1 0 40224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_420
timestamp 1679585382
transform 1 0 40896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_427
timestamp 1679585382
transform 1 0 41568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_434
timestamp 1679585382
transform 1 0 42240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_441
timestamp 1679585382
transform 1 0 42912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_448
timestamp 1679585382
transform 1 0 43584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_455
timestamp 1679585382
transform 1 0 44256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_462
timestamp 1679585382
transform 1 0 44928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_469
timestamp 1679585382
transform 1 0 45600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_476
timestamp 1679585382
transform 1 0 46272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_483
timestamp 1679585382
transform 1 0 46944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_490
timestamp 1679585382
transform 1 0 47616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_497
timestamp 1679585382
transform 1 0 48288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_504
timestamp 1679585382
transform 1 0 48960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_511
timestamp 1679585382
transform 1 0 49632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_518
timestamp 1679585382
transform 1 0 50304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_525
timestamp 1679585382
transform 1 0 50976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_532
timestamp 1679585382
transform 1 0 51648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_539
timestamp 1679585382
transform 1 0 52320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_546
timestamp 1679585382
transform 1 0 52992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_553
timestamp 1679585382
transform 1 0 53664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_560
timestamp 1679585382
transform 1 0 54336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_567
timestamp 1679585382
transform 1 0 55008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_574
timestamp 1679585382
transform 1 0 55680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_581
timestamp 1679585382
transform 1 0 56352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_588
timestamp 1679585382
transform 1 0 57024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_595
timestamp 1679585382
transform 1 0 57696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_602
timestamp 1679585382
transform 1 0 58368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_609
timestamp 1679585382
transform 1 0 59040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_616
timestamp 1679585382
transform 1 0 59712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_623
timestamp 1679585382
transform 1 0 60384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_630
timestamp 1679585382
transform 1 0 61056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_637
timestamp 1679585382
transform 1 0 61728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_644
timestamp 1679585382
transform 1 0 62400 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_651
timestamp 1679585382
transform 1 0 63072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_658
timestamp 1679585382
transform 1 0 63744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_665
timestamp 1679585382
transform 1 0 64416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_672
timestamp 1679585382
transform 1 0 65088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_679
timestamp 1679585382
transform 1 0 65760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_686
timestamp 1679585382
transform 1 0 66432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_693
timestamp 1679585382
transform 1 0 67104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_700
timestamp 1679585382
transform 1 0 67776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_707
timestamp 1679585382
transform 1 0 68448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_714
timestamp 1679585382
transform 1 0 69120 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_721
timestamp 1679585382
transform 1 0 69792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_728
timestamp 1679585382
transform 1 0 70464 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_735
timestamp 1679585382
transform 1 0 71136 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_742
timestamp 1679585382
transform 1 0 71808 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_749
timestamp 1679585382
transform 1 0 72480 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_756
timestamp 1679585382
transform 1 0 73152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_763
timestamp 1679585382
transform 1 0 73824 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_770
timestamp 1679585382
transform 1 0 74496 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_777
timestamp 1679585382
transform 1 0 75168 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_784
timestamp 1679585382
transform 1 0 75840 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_791
timestamp 1679585382
transform 1 0 76512 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_798
timestamp 1679585382
transform 1 0 77184 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_805
timestamp 1679585382
transform 1 0 77856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_812
timestamp 1679585382
transform 1 0 78528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_819
timestamp 1679585382
transform 1 0 79200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_826
timestamp 1679585382
transform 1 0 79872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_833
timestamp 1679585382
transform 1 0 80544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_840
timestamp 1679585382
transform 1 0 81216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_847
timestamp 1679585382
transform 1 0 81888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_854
timestamp 1679585382
transform 1 0 82560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_861
timestamp 1679585382
transform 1 0 83232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_868
timestamp 1679585382
transform 1 0 83904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_875
timestamp 1679585382
transform 1 0 84576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_882
timestamp 1679585382
transform 1 0 85248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_889
timestamp 1679585382
transform 1 0 85920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_896
timestamp 1679585382
transform 1 0 86592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_903
timestamp 1679585382
transform 1 0 87264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_910
timestamp 1679585382
transform 1 0 87936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_917
timestamp 1679585382
transform 1 0 88608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_924
timestamp 1679585382
transform 1 0 89280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_931
timestamp 1679585382
transform 1 0 89952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_938
timestamp 1679585382
transform 1 0 90624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_945
timestamp 1679585382
transform 1 0 91296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_952
timestamp 1679585382
transform 1 0 91968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_959
timestamp 1679585382
transform 1 0 92640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_966
timestamp 1679585382
transform 1 0 93312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_973
timestamp 1679585382
transform 1 0 93984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_980
timestamp 1679585382
transform 1 0 94656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_987
timestamp 1679585382
transform 1 0 95328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_994
timestamp 1679585382
transform 1 0 96000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1001
timestamp 1679585382
transform 1 0 96672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1008
timestamp 1679585382
transform 1 0 97344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1015
timestamp 1679585382
transform 1 0 98016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1022
timestamp 1679585382
transform 1 0 98688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679585382
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679585382
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679585382
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679585382
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679585382
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679585382
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679585382
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679585382
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679585382
transform 1 0 5952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679585382
transform 1 0 6624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679585382
transform 1 0 7296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679585382
transform 1 0 7968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679585382
transform 1 0 8640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679585382
transform 1 0 9312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679585382
transform 1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679585382
transform 1 0 10656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679585382
transform 1 0 11328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679585382
transform 1 0 12000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679585382
transform 1 0 12672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679585382
transform 1 0 13344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679585382
transform 1 0 14016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679585382
transform 1 0 14688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679585382
transform 1 0 15360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679585382
transform 1 0 16032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679585382
transform 1 0 16704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679585382
transform 1 0 17376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679585382
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679585382
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679585382
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679585382
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679585382
transform 1 0 20736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679585382
transform 1 0 21408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679585382
transform 1 0 22080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679585382
transform 1 0 22752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679585382
transform 1 0 23424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679585382
transform 1 0 24096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679585382
transform 1 0 24768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679585382
transform 1 0 25440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679585382
transform 1 0 26112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679585382
transform 1 0 26784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679585382
transform 1 0 27456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679585382
transform 1 0 28128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679585382
transform 1 0 28800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679585382
transform 1 0 29472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679585382
transform 1 0 30144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679585382
transform 1 0 30816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679585382
transform 1 0 31488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679585382
transform 1 0 32160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679585382
transform 1 0 32832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679585382
transform 1 0 33504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679585382
transform 1 0 34176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679585382
transform 1 0 34848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679585382
transform 1 0 35520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679585382
transform 1 0 36192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679585382
transform 1 0 36864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679585382
transform 1 0 37536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679585382
transform 1 0 38208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679585382
transform 1 0 38880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679585382
transform 1 0 39552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_413
timestamp 1679585382
transform 1 0 40224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_420
timestamp 1679585382
transform 1 0 40896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_427
timestamp 1679585382
transform 1 0 41568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_434
timestamp 1679585382
transform 1 0 42240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_441
timestamp 1679585382
transform 1 0 42912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_448
timestamp 1679585382
transform 1 0 43584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_455
timestamp 1679585382
transform 1 0 44256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_462
timestamp 1679585382
transform 1 0 44928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_469
timestamp 1679585382
transform 1 0 45600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_476
timestamp 1679585382
transform 1 0 46272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_483
timestamp 1679585382
transform 1 0 46944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_490
timestamp 1679585382
transform 1 0 47616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_497
timestamp 1679585382
transform 1 0 48288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_504
timestamp 1679585382
transform 1 0 48960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_511
timestamp 1679585382
transform 1 0 49632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_518
timestamp 1679585382
transform 1 0 50304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_525
timestamp 1679585382
transform 1 0 50976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_532
timestamp 1679585382
transform 1 0 51648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_539
timestamp 1679585382
transform 1 0 52320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_546
timestamp 1679585382
transform 1 0 52992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_553
timestamp 1679585382
transform 1 0 53664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_560
timestamp 1679585382
transform 1 0 54336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_567
timestamp 1679585382
transform 1 0 55008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_574
timestamp 1679585382
transform 1 0 55680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_581
timestamp 1679585382
transform 1 0 56352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_588
timestamp 1679585382
transform 1 0 57024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_595
timestamp 1679585382
transform 1 0 57696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_602
timestamp 1679585382
transform 1 0 58368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_609
timestamp 1679585382
transform 1 0 59040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_616
timestamp 1679585382
transform 1 0 59712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_623
timestamp 1679585382
transform 1 0 60384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_630
timestamp 1679585382
transform 1 0 61056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_637
timestamp 1679585382
transform 1 0 61728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_644
timestamp 1679585382
transform 1 0 62400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_651
timestamp 1679585382
transform 1 0 63072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_658
timestamp 1679585382
transform 1 0 63744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_665
timestamp 1679585382
transform 1 0 64416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_672
timestamp 1679585382
transform 1 0 65088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_679
timestamp 1679585382
transform 1 0 65760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_686
timestamp 1679585382
transform 1 0 66432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_693
timestamp 1679585382
transform 1 0 67104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_700
timestamp 1679585382
transform 1 0 67776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_707
timestamp 1679585382
transform 1 0 68448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_714
timestamp 1679585382
transform 1 0 69120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_721
timestamp 1679585382
transform 1 0 69792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_728
timestamp 1679585382
transform 1 0 70464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_735
timestamp 1679585382
transform 1 0 71136 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_742
timestamp 1679585382
transform 1 0 71808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_749
timestamp 1679585382
transform 1 0 72480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_756
timestamp 1679585382
transform 1 0 73152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_763
timestamp 1679585382
transform 1 0 73824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_770
timestamp 1679585382
transform 1 0 74496 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_777
timestamp 1679585382
transform 1 0 75168 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_784
timestamp 1679585382
transform 1 0 75840 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_791
timestamp 1679585382
transform 1 0 76512 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_798
timestamp 1679585382
transform 1 0 77184 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_805
timestamp 1679585382
transform 1 0 77856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_812
timestamp 1679585382
transform 1 0 78528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_819
timestamp 1679585382
transform 1 0 79200 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_826
timestamp 1679585382
transform 1 0 79872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_833
timestamp 1679585382
transform 1 0 80544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_840
timestamp 1679585382
transform 1 0 81216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_847
timestamp 1679585382
transform 1 0 81888 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_854
timestamp 1679585382
transform 1 0 82560 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_861
timestamp 1679585382
transform 1 0 83232 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_868
timestamp 1679585382
transform 1 0 83904 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_875
timestamp 1679585382
transform 1 0 84576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_882
timestamp 1679585382
transform 1 0 85248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_889
timestamp 1679585382
transform 1 0 85920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_896
timestamp 1679585382
transform 1 0 86592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_903
timestamp 1679585382
transform 1 0 87264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_910
timestamp 1679585382
transform 1 0 87936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_917
timestamp 1679585382
transform 1 0 88608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_924
timestamp 1679585382
transform 1 0 89280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_931
timestamp 1679585382
transform 1 0 89952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_938
timestamp 1679585382
transform 1 0 90624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_945
timestamp 1679585382
transform 1 0 91296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_952
timestamp 1679585382
transform 1 0 91968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_959
timestamp 1679585382
transform 1 0 92640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_966
timestamp 1679585382
transform 1 0 93312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_973
timestamp 1679585382
transform 1 0 93984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_980
timestamp 1679585382
transform 1 0 94656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_987
timestamp 1679585382
transform 1 0 95328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_994
timestamp 1679585382
transform 1 0 96000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1001
timestamp 1679585382
transform 1 0 96672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1008
timestamp 1679585382
transform 1 0 97344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1015
timestamp 1679585382
transform 1 0 98016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1022
timestamp 1679585382
transform 1 0 98688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679585382
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679585382
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679585382
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679585382
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679585382
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679585382
transform 1 0 3936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679585382
transform 1 0 4608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679585382
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679585382
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679585382
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679585382
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679585382
transform 1 0 7968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679585382
transform 1 0 8640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679585382
transform 1 0 9312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679585382
transform 1 0 9984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679585382
transform 1 0 10656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679585382
transform 1 0 11328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679585382
transform 1 0 12000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679585382
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679585382
transform 1 0 13344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679585382
transform 1 0 14016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679585382
transform 1 0 14688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679585382
transform 1 0 15360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679585382
transform 1 0 16032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679585382
transform 1 0 16704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679585382
transform 1 0 17376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679585382
transform 1 0 18048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679585382
transform 1 0 18720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679585382
transform 1 0 19392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679585382
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679585382
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679585382
transform 1 0 21408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679585382
transform 1 0 22080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679585382
transform 1 0 22752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679585382
transform 1 0 23424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679585382
transform 1 0 24096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679585382
transform 1 0 24768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679585382
transform 1 0 25440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679585382
transform 1 0 26112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679585382
transform 1 0 26784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679585382
transform 1 0 27456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679585382
transform 1 0 28128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679585382
transform 1 0 28800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679585382
transform 1 0 29472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679585382
transform 1 0 30144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679585382
transform 1 0 30816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679585382
transform 1 0 31488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679585382
transform 1 0 32160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679585382
transform 1 0 32832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679585382
transform 1 0 33504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679585382
transform 1 0 34176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679585382
transform 1 0 34848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679585382
transform 1 0 35520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679585382
transform 1 0 36192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679585382
transform 1 0 36864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679585382
transform 1 0 37536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679585382
transform 1 0 38208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679585382
transform 1 0 38880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679585382
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679585382
transform 1 0 40224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_420
timestamp 1679585382
transform 1 0 40896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_427
timestamp 1679585382
transform 1 0 41568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_434
timestamp 1679585382
transform 1 0 42240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_441
timestamp 1679585382
transform 1 0 42912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_448
timestamp 1679585382
transform 1 0 43584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_455
timestamp 1679585382
transform 1 0 44256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_462
timestamp 1679585382
transform 1 0 44928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679585382
transform 1 0 45600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_476
timestamp 1679585382
transform 1 0 46272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_483
timestamp 1679585382
transform 1 0 46944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_490
timestamp 1679585382
transform 1 0 47616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_497
timestamp 1679585382
transform 1 0 48288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_504
timestamp 1679585382
transform 1 0 48960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_511
timestamp 1679585382
transform 1 0 49632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_518
timestamp 1679585382
transform 1 0 50304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_525
timestamp 1679585382
transform 1 0 50976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_532
timestamp 1679585382
transform 1 0 51648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_539
timestamp 1679585382
transform 1 0 52320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_546
timestamp 1679585382
transform 1 0 52992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679585382
transform 1 0 53664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_560
timestamp 1679585382
transform 1 0 54336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_567
timestamp 1679585382
transform 1 0 55008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_574
timestamp 1679585382
transform 1 0 55680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_581
timestamp 1679585382
transform 1 0 56352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_588
timestamp 1679585382
transform 1 0 57024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_595
timestamp 1679585382
transform 1 0 57696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_602
timestamp 1679585382
transform 1 0 58368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_609
timestamp 1679585382
transform 1 0 59040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_616
timestamp 1679585382
transform 1 0 59712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_623
timestamp 1679585382
transform 1 0 60384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_630
timestamp 1679585382
transform 1 0 61056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679585382
transform 1 0 61728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_644
timestamp 1679585382
transform 1 0 62400 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_651
timestamp 1679585382
transform 1 0 63072 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_658
timestamp 1679585382
transform 1 0 63744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_665
timestamp 1679585382
transform 1 0 64416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_672
timestamp 1679585382
transform 1 0 65088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_679
timestamp 1679585382
transform 1 0 65760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_686
timestamp 1679585382
transform 1 0 66432 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_693
timestamp 1679585382
transform 1 0 67104 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_700
timestamp 1679585382
transform 1 0 67776 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_707
timestamp 1679585382
transform 1 0 68448 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_714
timestamp 1679585382
transform 1 0 69120 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_721
timestamp 1679585382
transform 1 0 69792 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_728
timestamp 1679585382
transform 1 0 70464 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_735
timestamp 1679585382
transform 1 0 71136 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_742
timestamp 1679585382
transform 1 0 71808 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_749
timestamp 1679585382
transform 1 0 72480 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_756
timestamp 1679585382
transform 1 0 73152 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_763
timestamp 1679585382
transform 1 0 73824 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_770
timestamp 1679585382
transform 1 0 74496 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_777
timestamp 1679585382
transform 1 0 75168 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_784
timestamp 1679585382
transform 1 0 75840 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_791
timestamp 1679585382
transform 1 0 76512 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_798
timestamp 1679585382
transform 1 0 77184 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_805
timestamp 1679585382
transform 1 0 77856 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_812
timestamp 1679585382
transform 1 0 78528 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_819
timestamp 1679585382
transform 1 0 79200 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_826
timestamp 1679585382
transform 1 0 79872 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_833
timestamp 1679585382
transform 1 0 80544 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_840
timestamp 1679585382
transform 1 0 81216 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_847
timestamp 1679585382
transform 1 0 81888 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_854
timestamp 1679585382
transform 1 0 82560 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_861
timestamp 1679585382
transform 1 0 83232 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_868
timestamp 1679585382
transform 1 0 83904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_875
timestamp 1679585382
transform 1 0 84576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_882
timestamp 1679585382
transform 1 0 85248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_889
timestamp 1679585382
transform 1 0 85920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_896
timestamp 1679585382
transform 1 0 86592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_903
timestamp 1679585382
transform 1 0 87264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_910
timestamp 1679585382
transform 1 0 87936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_917
timestamp 1679585382
transform 1 0 88608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_924
timestamp 1679585382
transform 1 0 89280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_931
timestamp 1679585382
transform 1 0 89952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_938
timestamp 1679585382
transform 1 0 90624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_945
timestamp 1679585382
transform 1 0 91296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_952
timestamp 1679585382
transform 1 0 91968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_959
timestamp 1679585382
transform 1 0 92640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_966
timestamp 1679585382
transform 1 0 93312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_973
timestamp 1679585382
transform 1 0 93984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_980
timestamp 1679585382
transform 1 0 94656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_987
timestamp 1679585382
transform 1 0 95328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_994
timestamp 1679585382
transform 1 0 96000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1001
timestamp 1679585382
transform 1 0 96672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1008
timestamp 1679585382
transform 1 0 97344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1015
timestamp 1679585382
transform 1 0 98016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1022
timestamp 1679585382
transform 1 0 98688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679585382
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679585382
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679585382
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679585382
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679585382
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679585382
transform 1 0 3936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679585382
transform 1 0 4608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679585382
transform 1 0 5280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679585382
transform 1 0 5952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679585382
transform 1 0 6624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679585382
transform 1 0 7296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679585382
transform 1 0 7968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679585382
transform 1 0 8640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679585382
transform 1 0 9312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679585382
transform 1 0 9984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679585382
transform 1 0 10656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679585382
transform 1 0 11328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679585382
transform 1 0 12000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679585382
transform 1 0 12672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679585382
transform 1 0 13344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679585382
transform 1 0 14016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679585382
transform 1 0 14688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679585382
transform 1 0 15360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679585382
transform 1 0 16032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679585382
transform 1 0 16704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679585382
transform 1 0 17376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679585382
transform 1 0 18048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679585382
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679585382
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679585382
transform 1 0 20064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679585382
transform 1 0 20736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679585382
transform 1 0 21408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679585382
transform 1 0 22080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679585382
transform 1 0 22752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679585382
transform 1 0 23424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679585382
transform 1 0 24096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679585382
transform 1 0 24768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679585382
transform 1 0 25440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679585382
transform 1 0 26112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679585382
transform 1 0 26784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679585382
transform 1 0 27456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679585382
transform 1 0 28128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679585382
transform 1 0 28800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679585382
transform 1 0 29472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679585382
transform 1 0 30144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679585382
transform 1 0 30816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679585382
transform 1 0 31488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679585382
transform 1 0 32160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679585382
transform 1 0 32832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679585382
transform 1 0 33504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679585382
transform 1 0 34176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679585382
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679585382
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679585382
transform 1 0 36192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679585382
transform 1 0 36864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679585382
transform 1 0 37536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679585382
transform 1 0 38208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679585382
transform 1 0 38880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_406
timestamp 1679585382
transform 1 0 39552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_413
timestamp 1679585382
transform 1 0 40224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679585382
transform 1 0 40896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_427
timestamp 1679585382
transform 1 0 41568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679585382
transform 1 0 42240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_441
timestamp 1679585382
transform 1 0 42912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_448
timestamp 1679585382
transform 1 0 43584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_455
timestamp 1679585382
transform 1 0 44256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_462
timestamp 1679585382
transform 1 0 44928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_469
timestamp 1679585382
transform 1 0 45600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_476
timestamp 1679585382
transform 1 0 46272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679585382
transform 1 0 46944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679585382
transform 1 0 47616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_497
timestamp 1679585382
transform 1 0 48288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_504
timestamp 1679585382
transform 1 0 48960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_511
timestamp 1679585382
transform 1 0 49632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_518
timestamp 1679585382
transform 1 0 50304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_525
timestamp 1679585382
transform 1 0 50976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_532
timestamp 1679585382
transform 1 0 51648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_539
timestamp 1679585382
transform 1 0 52320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_546
timestamp 1679585382
transform 1 0 52992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_553
timestamp 1679585382
transform 1 0 53664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_560
timestamp 1679585382
transform 1 0 54336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_567
timestamp 1679585382
transform 1 0 55008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_574
timestamp 1679585382
transform 1 0 55680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_581
timestamp 1679585382
transform 1 0 56352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_588
timestamp 1679585382
transform 1 0 57024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_595
timestamp 1679585382
transform 1 0 57696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_602
timestamp 1679585382
transform 1 0 58368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_609
timestamp 1679585382
transform 1 0 59040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_616
timestamp 1679585382
transform 1 0 59712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_623
timestamp 1679585382
transform 1 0 60384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_630
timestamp 1679585382
transform 1 0 61056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_637
timestamp 1679585382
transform 1 0 61728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_644
timestamp 1679585382
transform 1 0 62400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_651
timestamp 1679585382
transform 1 0 63072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_658
timestamp 1679585382
transform 1 0 63744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_665
timestamp 1679585382
transform 1 0 64416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_672
timestamp 1679585382
transform 1 0 65088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_679
timestamp 1679585382
transform 1 0 65760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_686
timestamp 1679585382
transform 1 0 66432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_693
timestamp 1679585382
transform 1 0 67104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_700
timestamp 1679585382
transform 1 0 67776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_707
timestamp 1679585382
transform 1 0 68448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_714
timestamp 1679585382
transform 1 0 69120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_721
timestamp 1679585382
transform 1 0 69792 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_728
timestamp 1679585382
transform 1 0 70464 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_735
timestamp 1679585382
transform 1 0 71136 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_742
timestamp 1679585382
transform 1 0 71808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_749
timestamp 1679585382
transform 1 0 72480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_756
timestamp 1679585382
transform 1 0 73152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_763
timestamp 1679585382
transform 1 0 73824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_770
timestamp 1679585382
transform 1 0 74496 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_777
timestamp 1679585382
transform 1 0 75168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_784
timestamp 1679585382
transform 1 0 75840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_791
timestamp 1679585382
transform 1 0 76512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_798
timestamp 1679585382
transform 1 0 77184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_805
timestamp 1679585382
transform 1 0 77856 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_812
timestamp 1679585382
transform 1 0 78528 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_819
timestamp 1679585382
transform 1 0 79200 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_826
timestamp 1679585382
transform 1 0 79872 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_833
timestamp 1679585382
transform 1 0 80544 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_840
timestamp 1679585382
transform 1 0 81216 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_847
timestamp 1679585382
transform 1 0 81888 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_854
timestamp 1679585382
transform 1 0 82560 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_861
timestamp 1679585382
transform 1 0 83232 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_868
timestamp 1679585382
transform 1 0 83904 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_875
timestamp 1679585382
transform 1 0 84576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_882
timestamp 1679585382
transform 1 0 85248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_889
timestamp 1679585382
transform 1 0 85920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_896
timestamp 1679585382
transform 1 0 86592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_903
timestamp 1679585382
transform 1 0 87264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_910
timestamp 1679585382
transform 1 0 87936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_917
timestamp 1679585382
transform 1 0 88608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_924
timestamp 1679585382
transform 1 0 89280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_931
timestamp 1679585382
transform 1 0 89952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_938
timestamp 1679585382
transform 1 0 90624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_945
timestamp 1679585382
transform 1 0 91296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_952
timestamp 1679585382
transform 1 0 91968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_959
timestamp 1679585382
transform 1 0 92640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_966
timestamp 1679585382
transform 1 0 93312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_973
timestamp 1679585382
transform 1 0 93984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_980
timestamp 1679585382
transform 1 0 94656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_987
timestamp 1679585382
transform 1 0 95328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_994
timestamp 1679585382
transform 1 0 96000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1001
timestamp 1679585382
transform 1 0 96672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1008
timestamp 1679585382
transform 1 0 97344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1015
timestamp 1679585382
transform 1 0 98016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1022
timestamp 1679585382
transform 1 0 98688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679585382
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679585382
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679585382
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679585382
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679585382
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679585382
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679585382
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679585382
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679585382
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679585382
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679585382
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679585382
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679585382
transform 1 0 8640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679585382
transform 1 0 9312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679585382
transform 1 0 9984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679585382
transform 1 0 10656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679585382
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679585382
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679585382
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679585382
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679585382
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679585382
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679585382
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679585382
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679585382
transform 1 0 16704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679585382
transform 1 0 17376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679585382
transform 1 0 18048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679585382
transform 1 0 18720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679585382
transform 1 0 19392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679585382
transform 1 0 20064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679585382
transform 1 0 20736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679585382
transform 1 0 21408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679585382
transform 1 0 22080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679585382
transform 1 0 22752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679585382
transform 1 0 23424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679585382
transform 1 0 24096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679585382
transform 1 0 24768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679585382
transform 1 0 25440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679585382
transform 1 0 26112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679585382
transform 1 0 26784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679585382
transform 1 0 27456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679585382
transform 1 0 28128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679585382
transform 1 0 28800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679585382
transform 1 0 29472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679585382
transform 1 0 30144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679585382
transform 1 0 30816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679585382
transform 1 0 31488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679585382
transform 1 0 32160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679585382
transform 1 0 32832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679585382
transform 1 0 33504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679585382
transform 1 0 34176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679585382
transform 1 0 34848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679585382
transform 1 0 35520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679585382
transform 1 0 36192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679585382
transform 1 0 36864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679585382
transform 1 0 37536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679585382
transform 1 0 38208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679585382
transform 1 0 38880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679585382
transform 1 0 39552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_413
timestamp 1679585382
transform 1 0 40224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679585382
transform 1 0 40896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679585382
transform 1 0 41568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_434
timestamp 1679585382
transform 1 0 42240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_441
timestamp 1679585382
transform 1 0 42912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_448
timestamp 1679585382
transform 1 0 43584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_455
timestamp 1679585382
transform 1 0 44256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_462
timestamp 1679585382
transform 1 0 44928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_469
timestamp 1679585382
transform 1 0 45600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_476
timestamp 1679585382
transform 1 0 46272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_483
timestamp 1679585382
transform 1 0 46944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_490
timestamp 1679585382
transform 1 0 47616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_497
timestamp 1679585382
transform 1 0 48288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_504
timestamp 1679585382
transform 1 0 48960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_511
timestamp 1679585382
transform 1 0 49632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_518
timestamp 1679585382
transform 1 0 50304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_525
timestamp 1679585382
transform 1 0 50976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_532
timestamp 1679585382
transform 1 0 51648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_539
timestamp 1679585382
transform 1 0 52320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_546
timestamp 1679585382
transform 1 0 52992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_553
timestamp 1679585382
transform 1 0 53664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_560
timestamp 1679585382
transform 1 0 54336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_567
timestamp 1679585382
transform 1 0 55008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_574
timestamp 1679585382
transform 1 0 55680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_581
timestamp 1679585382
transform 1 0 56352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_588
timestamp 1679585382
transform 1 0 57024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_595
timestamp 1679585382
transform 1 0 57696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_602
timestamp 1679585382
transform 1 0 58368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_609
timestamp 1679585382
transform 1 0 59040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_616
timestamp 1679585382
transform 1 0 59712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_623
timestamp 1679585382
transform 1 0 60384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_630
timestamp 1679585382
transform 1 0 61056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_637
timestamp 1679585382
transform 1 0 61728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_644
timestamp 1679585382
transform 1 0 62400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_651
timestamp 1679585382
transform 1 0 63072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_658
timestamp 1679585382
transform 1 0 63744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_665
timestamp 1679585382
transform 1 0 64416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_672
timestamp 1679585382
transform 1 0 65088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_679
timestamp 1679585382
transform 1 0 65760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_686
timestamp 1679585382
transform 1 0 66432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_693
timestamp 1679585382
transform 1 0 67104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_700
timestamp 1679585382
transform 1 0 67776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_707
timestamp 1679585382
transform 1 0 68448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_714
timestamp 1679585382
transform 1 0 69120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_721
timestamp 1679585382
transform 1 0 69792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_728
timestamp 1679585382
transform 1 0 70464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_735
timestamp 1679585382
transform 1 0 71136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_742
timestamp 1679585382
transform 1 0 71808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_749
timestamp 1679585382
transform 1 0 72480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_756
timestamp 1679585382
transform 1 0 73152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_763
timestamp 1679585382
transform 1 0 73824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_770
timestamp 1679585382
transform 1 0 74496 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_777
timestamp 1679585382
transform 1 0 75168 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_784
timestamp 1679585382
transform 1 0 75840 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_791
timestamp 1679585382
transform 1 0 76512 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_798
timestamp 1679585382
transform 1 0 77184 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_805
timestamp 1679585382
transform 1 0 77856 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_812
timestamp 1679585382
transform 1 0 78528 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_819
timestamp 1679585382
transform 1 0 79200 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_826
timestamp 1679585382
transform 1 0 79872 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_833
timestamp 1679585382
transform 1 0 80544 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_840
timestamp 1679585382
transform 1 0 81216 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_847
timestamp 1679585382
transform 1 0 81888 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_854
timestamp 1679585382
transform 1 0 82560 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_861
timestamp 1679585382
transform 1 0 83232 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_868
timestamp 1679585382
transform 1 0 83904 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_875
timestamp 1679585382
transform 1 0 84576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_882
timestamp 1679585382
transform 1 0 85248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_889
timestamp 1679585382
transform 1 0 85920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_896
timestamp 1679585382
transform 1 0 86592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_903
timestamp 1679585382
transform 1 0 87264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_910
timestamp 1679585382
transform 1 0 87936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_917
timestamp 1679585382
transform 1 0 88608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_924
timestamp 1679585382
transform 1 0 89280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_931
timestamp 1679585382
transform 1 0 89952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_938
timestamp 1679585382
transform 1 0 90624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_945
timestamp 1679585382
transform 1 0 91296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_952
timestamp 1679585382
transform 1 0 91968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_959
timestamp 1679585382
transform 1 0 92640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_966
timestamp 1679585382
transform 1 0 93312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_973
timestamp 1679585382
transform 1 0 93984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_980
timestamp 1679585382
transform 1 0 94656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_987
timestamp 1679585382
transform 1 0 95328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_994
timestamp 1679585382
transform 1 0 96000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1001
timestamp 1679585382
transform 1 0 96672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1008
timestamp 1679585382
transform 1 0 97344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1015
timestamp 1679585382
transform 1 0 98016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1022
timestamp 1679585382
transform 1 0 98688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679585382
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679585382
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679585382
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679585382
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679585382
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679585382
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679585382
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679585382
transform 1 0 5280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679585382
transform 1 0 5952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679585382
transform 1 0 6624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679585382
transform 1 0 7296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679585382
transform 1 0 7968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679585382
transform 1 0 8640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679585382
transform 1 0 9312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679585382
transform 1 0 9984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679585382
transform 1 0 10656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679585382
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679585382
transform 1 0 12000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679585382
transform 1 0 12672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679585382
transform 1 0 13344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679585382
transform 1 0 14016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679585382
transform 1 0 14688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679585382
transform 1 0 15360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679585382
transform 1 0 16032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679585382
transform 1 0 16704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679585382
transform 1 0 17376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679585382
transform 1 0 18048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679585382
transform 1 0 18720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679585382
transform 1 0 19392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679585382
transform 1 0 20064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679585382
transform 1 0 20736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679585382
transform 1 0 21408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679585382
transform 1 0 22080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679585382
transform 1 0 22752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679585382
transform 1 0 23424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679585382
transform 1 0 24096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679585382
transform 1 0 24768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679585382
transform 1 0 25440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679585382
transform 1 0 26112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679585382
transform 1 0 26784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679585382
transform 1 0 27456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679585382
transform 1 0 28128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679585382
transform 1 0 28800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679585382
transform 1 0 29472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679585382
transform 1 0 30144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679585382
transform 1 0 30816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679585382
transform 1 0 31488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679585382
transform 1 0 32160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679585382
transform 1 0 32832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679585382
transform 1 0 33504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679585382
transform 1 0 34176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679585382
transform 1 0 34848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679585382
transform 1 0 35520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679585382
transform 1 0 36192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679585382
transform 1 0 36864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679585382
transform 1 0 37536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679585382
transform 1 0 38208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679585382
transform 1 0 38880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679585382
transform 1 0 39552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679585382
transform 1 0 40224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679585382
transform 1 0 40896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679585382
transform 1 0 41568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_434
timestamp 1679585382
transform 1 0 42240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_441
timestamp 1679585382
transform 1 0 42912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_448
timestamp 1679585382
transform 1 0 43584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_455
timestamp 1679585382
transform 1 0 44256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_462
timestamp 1679585382
transform 1 0 44928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_469
timestamp 1679585382
transform 1 0 45600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_476
timestamp 1679585382
transform 1 0 46272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_483
timestamp 1679585382
transform 1 0 46944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_490
timestamp 1679585382
transform 1 0 47616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_497
timestamp 1679585382
transform 1 0 48288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_504
timestamp 1679585382
transform 1 0 48960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_511
timestamp 1679585382
transform 1 0 49632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_518
timestamp 1679585382
transform 1 0 50304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_525
timestamp 1679585382
transform 1 0 50976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_532
timestamp 1679585382
transform 1 0 51648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_539
timestamp 1679585382
transform 1 0 52320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_546
timestamp 1679585382
transform 1 0 52992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_553
timestamp 1679585382
transform 1 0 53664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_560
timestamp 1679585382
transform 1 0 54336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_567
timestamp 1679585382
transform 1 0 55008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_574
timestamp 1679585382
transform 1 0 55680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_581
timestamp 1679585382
transform 1 0 56352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_588
timestamp 1679585382
transform 1 0 57024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_595
timestamp 1679585382
transform 1 0 57696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_602
timestamp 1679585382
transform 1 0 58368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_609
timestamp 1679585382
transform 1 0 59040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_616
timestamp 1679585382
transform 1 0 59712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_623
timestamp 1679585382
transform 1 0 60384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_630
timestamp 1679585382
transform 1 0 61056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_637
timestamp 1679585382
transform 1 0 61728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_644
timestamp 1679585382
transform 1 0 62400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_651
timestamp 1679585382
transform 1 0 63072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_658
timestamp 1679585382
transform 1 0 63744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_665
timestamp 1679585382
transform 1 0 64416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_672
timestamp 1679585382
transform 1 0 65088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_679
timestamp 1679585382
transform 1 0 65760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_686
timestamp 1679585382
transform 1 0 66432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_693
timestamp 1679585382
transform 1 0 67104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_700
timestamp 1679585382
transform 1 0 67776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_707
timestamp 1679585382
transform 1 0 68448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_714
timestamp 1679585382
transform 1 0 69120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_721
timestamp 1679585382
transform 1 0 69792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_728
timestamp 1679585382
transform 1 0 70464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_735
timestamp 1679585382
transform 1 0 71136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_742
timestamp 1679585382
transform 1 0 71808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_749
timestamp 1679585382
transform 1 0 72480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_756
timestamp 1679585382
transform 1 0 73152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_763
timestamp 1679585382
transform 1 0 73824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_770
timestamp 1679585382
transform 1 0 74496 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_777
timestamp 1679585382
transform 1 0 75168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_784
timestamp 1679585382
transform 1 0 75840 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_791
timestamp 1679585382
transform 1 0 76512 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_798
timestamp 1679585382
transform 1 0 77184 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_805
timestamp 1679585382
transform 1 0 77856 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_812
timestamp 1679585382
transform 1 0 78528 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_819
timestamp 1679585382
transform 1 0 79200 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_826
timestamp 1679585382
transform 1 0 79872 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_833
timestamp 1679585382
transform 1 0 80544 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_840
timestamp 1679585382
transform 1 0 81216 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_847
timestamp 1679585382
transform 1 0 81888 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_854
timestamp 1679585382
transform 1 0 82560 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_861
timestamp 1679585382
transform 1 0 83232 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_868
timestamp 1679585382
transform 1 0 83904 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_875
timestamp 1679585382
transform 1 0 84576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_882
timestamp 1679585382
transform 1 0 85248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_889
timestamp 1679585382
transform 1 0 85920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_896
timestamp 1679585382
transform 1 0 86592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_903
timestamp 1679585382
transform 1 0 87264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_910
timestamp 1679585382
transform 1 0 87936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_917
timestamp 1679585382
transform 1 0 88608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_924
timestamp 1679585382
transform 1 0 89280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_931
timestamp 1679585382
transform 1 0 89952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_938
timestamp 1679585382
transform 1 0 90624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_945
timestamp 1679585382
transform 1 0 91296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_952
timestamp 1679585382
transform 1 0 91968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_959
timestamp 1679585382
transform 1 0 92640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_966
timestamp 1679585382
transform 1 0 93312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_973
timestamp 1679585382
transform 1 0 93984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_980
timestamp 1679585382
transform 1 0 94656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_987
timestamp 1679585382
transform 1 0 95328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_994
timestamp 1679585382
transform 1 0 96000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1001
timestamp 1679585382
transform 1 0 96672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1008
timestamp 1679585382
transform 1 0 97344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1015
timestamp 1679585382
transform 1 0 98016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1022
timestamp 1679585382
transform 1 0 98688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679585382
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679585382
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679585382
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679585382
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679585382
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679585382
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679585382
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679585382
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679585382
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679585382
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679585382
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679585382
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679585382
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679585382
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679585382
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679585382
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679585382
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679585382
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679585382
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679585382
transform 1 0 13344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679585382
transform 1 0 14016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679585382
transform 1 0 14688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679585382
transform 1 0 15360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679585382
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679585382
transform 1 0 16704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679585382
transform 1 0 17376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679585382
transform 1 0 18048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679585382
transform 1 0 18720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679585382
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679585382
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679585382
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679585382
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679585382
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679585382
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679585382
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679585382
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679585382
transform 1 0 24768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679585382
transform 1 0 25440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679585382
transform 1 0 26112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679585382
transform 1 0 26784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679585382
transform 1 0 27456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679585382
transform 1 0 28128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679585382
transform 1 0 28800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679585382
transform 1 0 29472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679585382
transform 1 0 30144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679585382
transform 1 0 30816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679585382
transform 1 0 31488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679585382
transform 1 0 32160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679585382
transform 1 0 32832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679585382
transform 1 0 33504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679585382
transform 1 0 34176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679585382
transform 1 0 34848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679585382
transform 1 0 35520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679585382
transform 1 0 36192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679585382
transform 1 0 36864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679585382
transform 1 0 37536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679585382
transform 1 0 38208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679585382
transform 1 0 38880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679585382
transform 1 0 39552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679585382
transform 1 0 40224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679585382
transform 1 0 40896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679585382
transform 1 0 41568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679585382
transform 1 0 42240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679585382
transform 1 0 42912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679585382
transform 1 0 43584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679585382
transform 1 0 44256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679585382
transform 1 0 44928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679585382
transform 1 0 45600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_476
timestamp 1679585382
transform 1 0 46272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_483
timestamp 1679585382
transform 1 0 46944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679585382
transform 1 0 47616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679585382
transform 1 0 48288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_504
timestamp 1679585382
transform 1 0 48960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679585382
transform 1 0 49632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679585382
transform 1 0 50304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_525
timestamp 1679585382
transform 1 0 50976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_532
timestamp 1679585382
transform 1 0 51648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_539
timestamp 1679585382
transform 1 0 52320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_546
timestamp 1679585382
transform 1 0 52992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_553
timestamp 1679585382
transform 1 0 53664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_560
timestamp 1679585382
transform 1 0 54336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_567
timestamp 1679585382
transform 1 0 55008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_574
timestamp 1679585382
transform 1 0 55680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_581
timestamp 1679585382
transform 1 0 56352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_588
timestamp 1679585382
transform 1 0 57024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_595
timestamp 1679585382
transform 1 0 57696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_602
timestamp 1679585382
transform 1 0 58368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_609
timestamp 1679585382
transform 1 0 59040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_616
timestamp 1679585382
transform 1 0 59712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_623
timestamp 1679585382
transform 1 0 60384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_630
timestamp 1679585382
transform 1 0 61056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_637
timestamp 1679585382
transform 1 0 61728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_644
timestamp 1679585382
transform 1 0 62400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_651
timestamp 1679585382
transform 1 0 63072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_658
timestamp 1679585382
transform 1 0 63744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_665
timestamp 1679585382
transform 1 0 64416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_672
timestamp 1679585382
transform 1 0 65088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_679
timestamp 1679585382
transform 1 0 65760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_686
timestamp 1679585382
transform 1 0 66432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_693
timestamp 1679585382
transform 1 0 67104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_700
timestamp 1679585382
transform 1 0 67776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_707
timestamp 1679585382
transform 1 0 68448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_714
timestamp 1679585382
transform 1 0 69120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_721
timestamp 1679585382
transform 1 0 69792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_728
timestamp 1679585382
transform 1 0 70464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_735
timestamp 1679585382
transform 1 0 71136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_742
timestamp 1679585382
transform 1 0 71808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_749
timestamp 1679585382
transform 1 0 72480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_756
timestamp 1679585382
transform 1 0 73152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_763
timestamp 1679585382
transform 1 0 73824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_770
timestamp 1679585382
transform 1 0 74496 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_777
timestamp 1679585382
transform 1 0 75168 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_784
timestamp 1679585382
transform 1 0 75840 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_791
timestamp 1679585382
transform 1 0 76512 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_798
timestamp 1679585382
transform 1 0 77184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_805
timestamp 1679585382
transform 1 0 77856 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_812
timestamp 1679585382
transform 1 0 78528 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_819
timestamp 1679585382
transform 1 0 79200 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_826
timestamp 1679585382
transform 1 0 79872 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_833
timestamp 1679585382
transform 1 0 80544 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_840
timestamp 1679585382
transform 1 0 81216 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_847
timestamp 1679585382
transform 1 0 81888 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_854
timestamp 1679585382
transform 1 0 82560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_861
timestamp 1679585382
transform 1 0 83232 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_868
timestamp 1679585382
transform 1 0 83904 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_875
timestamp 1679585382
transform 1 0 84576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_882
timestamp 1679585382
transform 1 0 85248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_889
timestamp 1679585382
transform 1 0 85920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_896
timestamp 1679585382
transform 1 0 86592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_903
timestamp 1679585382
transform 1 0 87264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_910
timestamp 1679585382
transform 1 0 87936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_917
timestamp 1679585382
transform 1 0 88608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_924
timestamp 1679585382
transform 1 0 89280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_931
timestamp 1679585382
transform 1 0 89952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_938
timestamp 1679585382
transform 1 0 90624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_945
timestamp 1679585382
transform 1 0 91296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_952
timestamp 1679585382
transform 1 0 91968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_959
timestamp 1679585382
transform 1 0 92640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_966
timestamp 1679585382
transform 1 0 93312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_973
timestamp 1679585382
transform 1 0 93984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_980
timestamp 1679585382
transform 1 0 94656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_987
timestamp 1679585382
transform 1 0 95328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_994
timestamp 1679585382
transform 1 0 96000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1001
timestamp 1679585382
transform 1 0 96672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1008
timestamp 1679585382
transform 1 0 97344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1015
timestamp 1679585382
transform 1 0 98016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1022
timestamp 1679585382
transform 1 0 98688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679585382
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679585382
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679585382
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679585382
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679585382
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679585382
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679585382
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679585382
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679585382
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679585382
transform 1 0 6624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679585382
transform 1 0 7296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679585382
transform 1 0 7968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679585382
transform 1 0 8640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679585382
transform 1 0 9312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679585382
transform 1 0 9984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679585382
transform 1 0 10656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679585382
transform 1 0 11328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679585382
transform 1 0 12000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679585382
transform 1 0 12672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679585382
transform 1 0 13344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679585382
transform 1 0 14016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679585382
transform 1 0 14688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679585382
transform 1 0 15360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679585382
transform 1 0 16032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679585382
transform 1 0 16704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679585382
transform 1 0 17376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679585382
transform 1 0 18048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679585382
transform 1 0 18720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679585382
transform 1 0 19392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679585382
transform 1 0 20064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679585382
transform 1 0 20736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679585382
transform 1 0 21408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679585382
transform 1 0 22080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679585382
transform 1 0 22752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679585382
transform 1 0 23424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679585382
transform 1 0 24096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679585382
transform 1 0 24768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679585382
transform 1 0 25440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679585382
transform 1 0 26112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679585382
transform 1 0 26784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679585382
transform 1 0 27456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679585382
transform 1 0 28128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679585382
transform 1 0 28800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679585382
transform 1 0 29472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679585382
transform 1 0 30144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679585382
transform 1 0 30816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679585382
transform 1 0 31488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679585382
transform 1 0 32160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679585382
transform 1 0 32832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679585382
transform 1 0 33504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679585382
transform 1 0 34176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679585382
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679585382
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679585382
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679585382
transform 1 0 36864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679585382
transform 1 0 37536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679585382
transform 1 0 38208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679585382
transform 1 0 38880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679585382
transform 1 0 39552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679585382
transform 1 0 40224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679585382
transform 1 0 40896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679585382
transform 1 0 41568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679585382
transform 1 0 42240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679585382
transform 1 0 42912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679585382
transform 1 0 43584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679585382
transform 1 0 44256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679585382
transform 1 0 44928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_469
timestamp 1679585382
transform 1 0 45600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_476
timestamp 1679585382
transform 1 0 46272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_483
timestamp 1679585382
transform 1 0 46944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_490
timestamp 1679585382
transform 1 0 47616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_497
timestamp 1679585382
transform 1 0 48288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_504
timestamp 1679585382
transform 1 0 48960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679585382
transform 1 0 49632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_518
timestamp 1679585382
transform 1 0 50304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_525
timestamp 1679585382
transform 1 0 50976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_532
timestamp 1679585382
transform 1 0 51648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_539
timestamp 1679585382
transform 1 0 52320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_546
timestamp 1679585382
transform 1 0 52992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_553
timestamp 1679585382
transform 1 0 53664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_560
timestamp 1679585382
transform 1 0 54336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_567
timestamp 1679585382
transform 1 0 55008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_574
timestamp 1679585382
transform 1 0 55680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_581
timestamp 1679585382
transform 1 0 56352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_588
timestamp 1679585382
transform 1 0 57024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_595
timestamp 1679585382
transform 1 0 57696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_602
timestamp 1679585382
transform 1 0 58368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_609
timestamp 1679585382
transform 1 0 59040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_616
timestamp 1679585382
transform 1 0 59712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_623
timestamp 1679585382
transform 1 0 60384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_630
timestamp 1679585382
transform 1 0 61056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_637
timestamp 1679585382
transform 1 0 61728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_644
timestamp 1679585382
transform 1 0 62400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_651
timestamp 1679585382
transform 1 0 63072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_658
timestamp 1679585382
transform 1 0 63744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_665
timestamp 1679585382
transform 1 0 64416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_672
timestamp 1679585382
transform 1 0 65088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_679
timestamp 1679585382
transform 1 0 65760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_686
timestamp 1679585382
transform 1 0 66432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_693
timestamp 1679585382
transform 1 0 67104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_700
timestamp 1679585382
transform 1 0 67776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_707
timestamp 1679585382
transform 1 0 68448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_714
timestamp 1679585382
transform 1 0 69120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_721
timestamp 1679585382
transform 1 0 69792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_728
timestamp 1679585382
transform 1 0 70464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_735
timestamp 1679585382
transform 1 0 71136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_742
timestamp 1679585382
transform 1 0 71808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_749
timestamp 1679585382
transform 1 0 72480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_756
timestamp 1679585382
transform 1 0 73152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_763
timestamp 1679585382
transform 1 0 73824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_770
timestamp 1679585382
transform 1 0 74496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_777
timestamp 1679585382
transform 1 0 75168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_784
timestamp 1679585382
transform 1 0 75840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_791
timestamp 1679585382
transform 1 0 76512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_798
timestamp 1679585382
transform 1 0 77184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_805
timestamp 1679585382
transform 1 0 77856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_812
timestamp 1679585382
transform 1 0 78528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_819
timestamp 1679585382
transform 1 0 79200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_826
timestamp 1679585382
transform 1 0 79872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_833
timestamp 1679585382
transform 1 0 80544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_840
timestamp 1679585382
transform 1 0 81216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_847
timestamp 1679585382
transform 1 0 81888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_854
timestamp 1679585382
transform 1 0 82560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_861
timestamp 1679585382
transform 1 0 83232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_868
timestamp 1679585382
transform 1 0 83904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_875
timestamp 1679585382
transform 1 0 84576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_882
timestamp 1679585382
transform 1 0 85248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_889
timestamp 1679585382
transform 1 0 85920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_896
timestamp 1679585382
transform 1 0 86592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_903
timestamp 1679585382
transform 1 0 87264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_910
timestamp 1679585382
transform 1 0 87936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_917
timestamp 1679585382
transform 1 0 88608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_924
timestamp 1679585382
transform 1 0 89280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_931
timestamp 1679585382
transform 1 0 89952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_938
timestamp 1679585382
transform 1 0 90624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_945
timestamp 1679585382
transform 1 0 91296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_952
timestamp 1679585382
transform 1 0 91968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_959
timestamp 1679585382
transform 1 0 92640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_966
timestamp 1679585382
transform 1 0 93312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_973
timestamp 1679585382
transform 1 0 93984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_980
timestamp 1679585382
transform 1 0 94656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_987
timestamp 1679585382
transform 1 0 95328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_994
timestamp 1679585382
transform 1 0 96000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1001
timestamp 1679585382
transform 1 0 96672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1008
timestamp 1679585382
transform 1 0 97344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1015
timestamp 1679585382
transform 1 0 98016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1022
timestamp 1679585382
transform 1 0 98688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679585382
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679585382
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679585382
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679585382
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679585382
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679585382
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679585382
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679585382
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679585382
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679585382
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679585382
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679585382
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679585382
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679585382
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679585382
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679585382
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679585382
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679585382
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679585382
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679585382
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679585382
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679585382
transform 1 0 14688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679585382
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679585382
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679585382
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679585382
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679585382
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679585382
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679585382
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679585382
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679585382
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679585382
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679585382
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679585382
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679585382
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679585382
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679585382
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679585382
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679585382
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679585382
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679585382
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679585382
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679585382
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679585382
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679585382
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679585382
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679585382
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679585382
transform 1 0 32160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679585382
transform 1 0 32832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679585382
transform 1 0 33504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679585382
transform 1 0 34176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679585382
transform 1 0 34848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679585382
transform 1 0 35520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679585382
transform 1 0 36192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679585382
transform 1 0 36864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679585382
transform 1 0 37536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679585382
transform 1 0 38208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679585382
transform 1 0 38880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679585382
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679585382
transform 1 0 40224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679585382
transform 1 0 40896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679585382
transform 1 0 41568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679585382
transform 1 0 42240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679585382
transform 1 0 42912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679585382
transform 1 0 43584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679585382
transform 1 0 44256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679585382
transform 1 0 44928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679585382
transform 1 0 45600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679585382
transform 1 0 46272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679585382
transform 1 0 46944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679585382
transform 1 0 47616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_497
timestamp 1679585382
transform 1 0 48288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_504
timestamp 1679585382
transform 1 0 48960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_511
timestamp 1679585382
transform 1 0 49632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_518
timestamp 1679585382
transform 1 0 50304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_525
timestamp 1679585382
transform 1 0 50976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_532
timestamp 1679585382
transform 1 0 51648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_539
timestamp 1679585382
transform 1 0 52320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_546
timestamp 1679585382
transform 1 0 52992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_553
timestamp 1679585382
transform 1 0 53664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_560
timestamp 1679585382
transform 1 0 54336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_567
timestamp 1679585382
transform 1 0 55008 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_574
timestamp 1679585382
transform 1 0 55680 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_581
timestamp 1679585382
transform 1 0 56352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_588
timestamp 1679585382
transform 1 0 57024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_595
timestamp 1679585382
transform 1 0 57696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_602
timestamp 1679585382
transform 1 0 58368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_609
timestamp 1679585382
transform 1 0 59040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_616
timestamp 1679585382
transform 1 0 59712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679585382
transform 1 0 60384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_630
timestamp 1679585382
transform 1 0 61056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_637
timestamp 1679585382
transform 1 0 61728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_644
timestamp 1679585382
transform 1 0 62400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_651
timestamp 1679585382
transform 1 0 63072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_658
timestamp 1679585382
transform 1 0 63744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_665
timestamp 1679585382
transform 1 0 64416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_672
timestamp 1679585382
transform 1 0 65088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_679
timestamp 1679585382
transform 1 0 65760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_686
timestamp 1679585382
transform 1 0 66432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_693
timestamp 1679585382
transform 1 0 67104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_700
timestamp 1679585382
transform 1 0 67776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_707
timestamp 1679585382
transform 1 0 68448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_714
timestamp 1679585382
transform 1 0 69120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_721
timestamp 1679585382
transform 1 0 69792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_728
timestamp 1679585382
transform 1 0 70464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_735
timestamp 1679585382
transform 1 0 71136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_742
timestamp 1679585382
transform 1 0 71808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_749
timestamp 1679585382
transform 1 0 72480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_756
timestamp 1679585382
transform 1 0 73152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_763
timestamp 1679585382
transform 1 0 73824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_770
timestamp 1679585382
transform 1 0 74496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_777
timestamp 1679585382
transform 1 0 75168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_784
timestamp 1679585382
transform 1 0 75840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_791
timestamp 1679585382
transform 1 0 76512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_798
timestamp 1679585382
transform 1 0 77184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_805
timestamp 1679585382
transform 1 0 77856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_812
timestamp 1679585382
transform 1 0 78528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_819
timestamp 1679585382
transform 1 0 79200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_826
timestamp 1679585382
transform 1 0 79872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_833
timestamp 1679585382
transform 1 0 80544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_840
timestamp 1679585382
transform 1 0 81216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_847
timestamp 1679585382
transform 1 0 81888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_854
timestamp 1679585382
transform 1 0 82560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_861
timestamp 1679585382
transform 1 0 83232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_868
timestamp 1679585382
transform 1 0 83904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_875
timestamp 1679585382
transform 1 0 84576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_882
timestamp 1679585382
transform 1 0 85248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_889
timestamp 1679585382
transform 1 0 85920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_896
timestamp 1679585382
transform 1 0 86592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_903
timestamp 1679585382
transform 1 0 87264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_910
timestamp 1679585382
transform 1 0 87936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_917
timestamp 1679585382
transform 1 0 88608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_924
timestamp 1679585382
transform 1 0 89280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_931
timestamp 1679585382
transform 1 0 89952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_938
timestamp 1679585382
transform 1 0 90624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_945
timestamp 1679585382
transform 1 0 91296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_952
timestamp 1679585382
transform 1 0 91968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_959
timestamp 1679585382
transform 1 0 92640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_966
timestamp 1679585382
transform 1 0 93312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_973
timestamp 1679585382
transform 1 0 93984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_980
timestamp 1679585382
transform 1 0 94656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_987
timestamp 1679585382
transform 1 0 95328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_994
timestamp 1679585382
transform 1 0 96000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1001
timestamp 1679585382
transform 1 0 96672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1008
timestamp 1679585382
transform 1 0 97344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1015
timestamp 1679585382
transform 1 0 98016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1022
timestamp 1679585382
transform 1 0 98688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679585382
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679585382
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679585382
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679585382
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679585382
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679585382
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679585382
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679585382
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679585382
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679585382
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679585382
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679585382
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679585382
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679585382
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679585382
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679585382
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679585382
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679585382
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679585382
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679585382
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679585382
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679585382
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679585382
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679585382
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679585382
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679585382
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679585382
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679585382
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679585382
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679585382
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679585382
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679585382
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679585382
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679585382
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679585382
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679585382
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679585382
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679585382
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679585382
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679585382
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679585382
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679585382
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679585382
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679585382
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679585382
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679585382
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679585382
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679585382
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679585382
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679585382
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679585382
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679585382
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679585382
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679585382
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679585382
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679585382
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679585382
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679585382
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679585382
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679585382
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679585382
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679585382
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679585382
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679585382
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679585382
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679585382
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679585382
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679585382
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679585382
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679585382
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679585382
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679585382
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679585382
transform 1 0 48960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679585382
transform 1 0 49632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679585382
transform 1 0 50304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679585382
transform 1 0 50976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679585382
transform 1 0 51648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679585382
transform 1 0 52320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679585382
transform 1 0 52992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679585382
transform 1 0 53664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679585382
transform 1 0 54336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679585382
transform 1 0 55008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679585382
transform 1 0 55680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679585382
transform 1 0 56352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679585382
transform 1 0 57024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679585382
transform 1 0 57696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679585382
transform 1 0 58368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679585382
transform 1 0 59040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679585382
transform 1 0 59712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679585382
transform 1 0 60384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679585382
transform 1 0 61056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679585382
transform 1 0 61728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679585382
transform 1 0 62400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679585382
transform 1 0 63072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679585382
transform 1 0 63744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679585382
transform 1 0 64416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679585382
transform 1 0 65088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679585382
transform 1 0 65760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679585382
transform 1 0 66432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679585382
transform 1 0 67104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679585382
transform 1 0 67776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679585382
transform 1 0 68448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679585382
transform 1 0 69120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679585382
transform 1 0 69792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679585382
transform 1 0 70464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679585382
transform 1 0 71136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679585382
transform 1 0 71808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679585382
transform 1 0 72480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_756
timestamp 1679585382
transform 1 0 73152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_763
timestamp 1679585382
transform 1 0 73824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_770
timestamp 1679585382
transform 1 0 74496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_777
timestamp 1679585382
transform 1 0 75168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_784
timestamp 1679585382
transform 1 0 75840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_791
timestamp 1679585382
transform 1 0 76512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_798
timestamp 1679585382
transform 1 0 77184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_805
timestamp 1679585382
transform 1 0 77856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_812
timestamp 1679585382
transform 1 0 78528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_819
timestamp 1679585382
transform 1 0 79200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_826
timestamp 1679585382
transform 1 0 79872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_833
timestamp 1679585382
transform 1 0 80544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_840
timestamp 1679585382
transform 1 0 81216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_847
timestamp 1679585382
transform 1 0 81888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_854
timestamp 1679585382
transform 1 0 82560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_861
timestamp 1679585382
transform 1 0 83232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_868
timestamp 1679585382
transform 1 0 83904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_875
timestamp 1679585382
transform 1 0 84576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_882
timestamp 1679585382
transform 1 0 85248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_889
timestamp 1679585382
transform 1 0 85920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_896
timestamp 1679585382
transform 1 0 86592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_903
timestamp 1679585382
transform 1 0 87264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_910
timestamp 1679585382
transform 1 0 87936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_917
timestamp 1679585382
transform 1 0 88608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_924
timestamp 1679585382
transform 1 0 89280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_931
timestamp 1679585382
transform 1 0 89952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_938
timestamp 1679585382
transform 1 0 90624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_945
timestamp 1679585382
transform 1 0 91296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_952
timestamp 1679585382
transform 1 0 91968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_959
timestamp 1679585382
transform 1 0 92640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_966
timestamp 1679585382
transform 1 0 93312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_973
timestamp 1679585382
transform 1 0 93984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_980
timestamp 1679585382
transform 1 0 94656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_987
timestamp 1679585382
transform 1 0 95328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_994
timestamp 1679585382
transform 1 0 96000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1001
timestamp 1679585382
transform 1 0 96672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1008
timestamp 1679585382
transform 1 0 97344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1015
timestamp 1679585382
transform 1 0 98016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1022
timestamp 1679585382
transform 1 0 98688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679585382
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679585382
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679585382
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679585382
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679585382
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679585382
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679585382
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679585382
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679585382
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679585382
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679585382
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679585382
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679585382
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679585382
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679585382
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679585382
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679585382
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679585382
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679585382
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679585382
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679585382
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679585382
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679585382
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679585382
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679585382
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679585382
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679585382
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679585382
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679585382
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679585382
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679585382
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679585382
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679585382
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679585382
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679585382
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679585382
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679585382
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679585382
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679585382
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679585382
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679585382
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679585382
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679585382
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679585382
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679585382
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679585382
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679585382
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679585382
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679585382
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679585382
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679585382
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679585382
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679585382
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679585382
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679585382
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679585382
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679585382
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679585382
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679585382
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679585382
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679585382
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679585382
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679585382
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679585382
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679585382
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679585382
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679585382
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679585382
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679585382
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679585382
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679585382
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679585382
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679585382
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679585382
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679585382
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679585382
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679585382
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679585382
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679585382
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679585382
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679585382
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679585382
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679585382
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679585382
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679585382
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679585382
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679585382
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679585382
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679585382
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679585382
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679585382
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679585382
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679585382
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679585382
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679585382
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679585382
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679585382
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679585382
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679585382
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679585382
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679585382
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679585382
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679585382
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679585382
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679585382
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679585382
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679585382
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679585382
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679585382
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679585382
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679585382
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679585382
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679585382
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679585382
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679585382
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679585382
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679585382
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679585382
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679585382
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679585382
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679585382
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679585382
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679585382
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_861
timestamp 1679585382
transform 1 0 83232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_868
timestamp 1679585382
transform 1 0 83904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_875
timestamp 1679585382
transform 1 0 84576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_882
timestamp 1679585382
transform 1 0 85248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_889
timestamp 1679585382
transform 1 0 85920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_896
timestamp 1679585382
transform 1 0 86592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_903
timestamp 1679585382
transform 1 0 87264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_910
timestamp 1679585382
transform 1 0 87936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_917
timestamp 1679585382
transform 1 0 88608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_924
timestamp 1679585382
transform 1 0 89280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_931
timestamp 1679585382
transform 1 0 89952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_938
timestamp 1679585382
transform 1 0 90624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_945
timestamp 1679585382
transform 1 0 91296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_952
timestamp 1679585382
transform 1 0 91968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_959
timestamp 1679585382
transform 1 0 92640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_966
timestamp 1679585382
transform 1 0 93312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_973
timestamp 1679585382
transform 1 0 93984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_980
timestamp 1679585382
transform 1 0 94656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_987
timestamp 1679585382
transform 1 0 95328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_994
timestamp 1679585382
transform 1 0 96000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1001
timestamp 1679585382
transform 1 0 96672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1008
timestamp 1679585382
transform 1 0 97344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1015
timestamp 1679585382
transform 1 0 98016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1022
timestamp 1679585382
transform 1 0 98688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679585382
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679585382
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679585382
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679585382
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679585382
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679585382
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679585382
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679585382
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679585382
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679585382
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679585382
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679585382
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679585382
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679585382
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679585382
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679585382
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679585382
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679585382
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679585382
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679585382
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679585382
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679585382
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679585382
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679585382
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679585382
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679585382
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679585382
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679585382
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679585382
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679585382
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679585382
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679585382
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679585382
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679585382
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679585382
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679585382
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679585382
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679585382
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679585382
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679585382
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679585382
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679585382
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679585382
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679585382
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679585382
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679585382
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679585382
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679585382
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679585382
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679585382
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679585382
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679585382
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679585382
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679585382
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679585382
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679585382
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679585382
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679585382
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679585382
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679585382
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679585382
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679585382
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679585382
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679585382
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679585382
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679585382
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679585382
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679585382
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679585382
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679585382
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679585382
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679585382
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679585382
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679585382
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679585382
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679585382
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679585382
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679585382
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679585382
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679585382
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679585382
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679585382
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679585382
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679585382
transform 1 0 56352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679585382
transform 1 0 57024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679585382
transform 1 0 57696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679585382
transform 1 0 58368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679585382
transform 1 0 59040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679585382
transform 1 0 59712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679585382
transform 1 0 60384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679585382
transform 1 0 61056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679585382
transform 1 0 61728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679585382
transform 1 0 62400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679585382
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679585382
transform 1 0 63744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679585382
transform 1 0 64416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679585382
transform 1 0 65088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679585382
transform 1 0 65760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679585382
transform 1 0 66432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679585382
transform 1 0 67104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679585382
transform 1 0 67776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679585382
transform 1 0 68448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679585382
transform 1 0 69120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679585382
transform 1 0 69792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679585382
transform 1 0 70464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679585382
transform 1 0 71136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679585382
transform 1 0 71808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679585382
transform 1 0 72480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679585382
transform 1 0 73152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679585382
transform 1 0 73824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679585382
transform 1 0 74496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679585382
transform 1 0 75168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679585382
transform 1 0 75840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679585382
transform 1 0 76512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679585382
transform 1 0 77184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679585382
transform 1 0 77856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679585382
transform 1 0 78528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679585382
transform 1 0 79200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679585382
transform 1 0 79872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679585382
transform 1 0 80544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_840
timestamp 1679585382
transform 1 0 81216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_847
timestamp 1679585382
transform 1 0 81888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_854
timestamp 1679585382
transform 1 0 82560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_861
timestamp 1679585382
transform 1 0 83232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_868
timestamp 1679585382
transform 1 0 83904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_875
timestamp 1679585382
transform 1 0 84576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_882
timestamp 1679585382
transform 1 0 85248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_889
timestamp 1679585382
transform 1 0 85920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_896
timestamp 1679585382
transform 1 0 86592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_903
timestamp 1679585382
transform 1 0 87264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_910
timestamp 1679585382
transform 1 0 87936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_917
timestamp 1679585382
transform 1 0 88608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_924
timestamp 1679585382
transform 1 0 89280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_931
timestamp 1679585382
transform 1 0 89952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_938
timestamp 1679585382
transform 1 0 90624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_945
timestamp 1679585382
transform 1 0 91296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_952
timestamp 1679585382
transform 1 0 91968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_959
timestamp 1679585382
transform 1 0 92640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_966
timestamp 1679585382
transform 1 0 93312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_973
timestamp 1679585382
transform 1 0 93984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_980
timestamp 1679585382
transform 1 0 94656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_987
timestamp 1679585382
transform 1 0 95328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_994
timestamp 1679585382
transform 1 0 96000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1001
timestamp 1679585382
transform 1 0 96672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1008
timestamp 1679585382
transform 1 0 97344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1015
timestamp 1679585382
transform 1 0 98016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1022
timestamp 1679585382
transform 1 0 98688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679585382
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679585382
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679585382
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679585382
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679585382
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679585382
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679585382
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679585382
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679585382
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679585382
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679585382
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679585382
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679585382
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679585382
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679585382
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679585382
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679585382
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679585382
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679585382
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679585382
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679585382
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679585382
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679585382
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679585382
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679585382
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679585382
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679585382
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679585382
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679585382
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679585382
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_214
timestamp 1679585382
transform 1 0 21120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_221
timestamp 1679585382
transform 1 0 21792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_228
timestamp 1679585382
transform 1 0 22464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_235
timestamp 1679585382
transform 1 0 23136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_242
timestamp 1679585382
transform 1 0 23808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_249
timestamp 1679585382
transform 1 0 24480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_256
timestamp 1679585382
transform 1 0 25152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_263
timestamp 1679585382
transform 1 0 25824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_270
timestamp 1679585382
transform 1 0 26496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_277
timestamp 1679585382
transform 1 0 27168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_284
timestamp 1679585382
transform 1 0 27840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_291
timestamp 1679585382
transform 1 0 28512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_298
timestamp 1679585382
transform 1 0 29184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_305
timestamp 1679585382
transform 1 0 29856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_312
timestamp 1679585382
transform 1 0 30528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_319
timestamp 1679585382
transform 1 0 31200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_326
timestamp 1679585382
transform 1 0 31872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_333
timestamp 1679585382
transform 1 0 32544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_340
timestamp 1679585382
transform 1 0 33216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_347
timestamp 1679585382
transform 1 0 33888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_354
timestamp 1679585382
transform 1 0 34560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_361
timestamp 1679585382
transform 1 0 35232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_368
timestamp 1679585382
transform 1 0 35904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_375
timestamp 1679585382
transform 1 0 36576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_382
timestamp 1679585382
transform 1 0 37248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_389
timestamp 1679585382
transform 1 0 37920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_396
timestamp 1679585382
transform 1 0 38592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679585382
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679585382
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_417
timestamp 1679585382
transform 1 0 40608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_424
timestamp 1679585382
transform 1 0 41280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_431
timestamp 1679585382
transform 1 0 41952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_438
timestamp 1679585382
transform 1 0 42624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_445
timestamp 1679585382
transform 1 0 43296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_452
timestamp 1679585382
transform 1 0 43968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_459
timestamp 1679585382
transform 1 0 44640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_466
timestamp 1679585382
transform 1 0 45312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_473
timestamp 1679585382
transform 1 0 45984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_480
timestamp 1679585382
transform 1 0 46656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_487
timestamp 1679585382
transform 1 0 47328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_494
timestamp 1679585382
transform 1 0 48000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_501
timestamp 1679585382
transform 1 0 48672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_508
timestamp 1679585382
transform 1 0 49344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_515
timestamp 1679585382
transform 1 0 50016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_522
timestamp 1679585382
transform 1 0 50688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_529
timestamp 1679585382
transform 1 0 51360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_536
timestamp 1679585382
transform 1 0 52032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_543
timestamp 1679585382
transform 1 0 52704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_550
timestamp 1679585382
transform 1 0 53376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_557
timestamp 1679585382
transform 1 0 54048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_564
timestamp 1679585382
transform 1 0 54720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_571
timestamp 1679585382
transform 1 0 55392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_578
timestamp 1679585382
transform 1 0 56064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_585
timestamp 1679585382
transform 1 0 56736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_592
timestamp 1679585382
transform 1 0 57408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_599
timestamp 1679585382
transform 1 0 58080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_606
timestamp 1679585382
transform 1 0 58752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_613
timestamp 1679585382
transform 1 0 59424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_620
timestamp 1679585382
transform 1 0 60096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_627
timestamp 1679585382
transform 1 0 60768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_634
timestamp 1679585382
transform 1 0 61440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_641
timestamp 1679585382
transform 1 0 62112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_648
timestamp 1679585382
transform 1 0 62784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_655
timestamp 1679585382
transform 1 0 63456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_662
timestamp 1679585382
transform 1 0 64128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_669
timestamp 1679585382
transform 1 0 64800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_676
timestamp 1679585382
transform 1 0 65472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_683
timestamp 1679585382
transform 1 0 66144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_690
timestamp 1679585382
transform 1 0 66816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_697
timestamp 1679585382
transform 1 0 67488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_704
timestamp 1679585382
transform 1 0 68160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_711
timestamp 1679585382
transform 1 0 68832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_718
timestamp 1679585382
transform 1 0 69504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_725
timestamp 1679585382
transform 1 0 70176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_732
timestamp 1679585382
transform 1 0 70848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_739
timestamp 1679585382
transform 1 0 71520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_746
timestamp 1679585382
transform 1 0 72192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_753
timestamp 1679585382
transform 1 0 72864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_760
timestamp 1679585382
transform 1 0 73536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_767
timestamp 1679585382
transform 1 0 74208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_774
timestamp 1679585382
transform 1 0 74880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_781
timestamp 1679585382
transform 1 0 75552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_788
timestamp 1679585382
transform 1 0 76224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_795
timestamp 1679585382
transform 1 0 76896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_802
timestamp 1679585382
transform 1 0 77568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_809
timestamp 1679585382
transform 1 0 78240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_816
timestamp 1679585382
transform 1 0 78912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_823
timestamp 1679585382
transform 1 0 79584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_830
timestamp 1679585382
transform 1 0 80256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_837
timestamp 1679585382
transform 1 0 80928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_844
timestamp 1679585382
transform 1 0 81600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_851
timestamp 1679585382
transform 1 0 82272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_858
timestamp 1679585382
transform 1 0 82944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_865
timestamp 1679585382
transform 1 0 83616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_872
timestamp 1679585382
transform 1 0 84288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_879
timestamp 1679585382
transform 1 0 84960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_886
timestamp 1679585382
transform 1 0 85632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_893
timestamp 1679585382
transform 1 0 86304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_900
timestamp 1679585382
transform 1 0 86976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_907
timestamp 1679585382
transform 1 0 87648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_914
timestamp 1679585382
transform 1 0 88320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_921
timestamp 1679585382
transform 1 0 88992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_928
timestamp 1679585382
transform 1 0 89664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_935
timestamp 1679585382
transform 1 0 90336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_942
timestamp 1679585382
transform 1 0 91008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_949
timestamp 1679585382
transform 1 0 91680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_956
timestamp 1679585382
transform 1 0 92352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_963
timestamp 1679585382
transform 1 0 93024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_970
timestamp 1679585382
transform 1 0 93696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_977
timestamp 1679585382
transform 1 0 94368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_984
timestamp 1679585382
transform 1 0 95040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_991
timestamp 1679585382
transform 1 0 95712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_998
timestamp 1679585382
transform 1 0 96384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1005
timestamp 1679585382
transform 1 0 97056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1012
timestamp 1679585382
transform 1 0 97728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1019
timestamp 1679585382
transform 1 0 98400 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_1026
timestamp 1677583704
transform 1 0 99072 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_1028
timestamp 1677583258
transform 1 0 99264 0 -1 38556
box -48 -56 144 834
use sg13g2_tiehi  heichips25_template_27
timestamp 1680007851
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_28
timestamp 1680007851
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_29
timestamp 1680007851
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_30
timestamp 1680007851
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_31
timestamp 1680007851
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_32
timestamp 1680007851
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_33
timestamp 1680007851
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template
timestamp 1680007851
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1677675658
transform -1 0 3744 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1677675658
transform 1 0 3360 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1677675658
transform -1 0 10272 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1677675658
transform -1 0 8928 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1677675658
transform -1 0 14208 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1677675658
transform -1 0 10944 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1677675658
transform 1 0 12000 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1677675658
transform -1 0 5952 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1677675658
transform -1 0 5088 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1677675658
transform -1 0 4896 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1677675658
transform -1 0 12192 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1677675658
transform 1 0 10368 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1677675658
transform -1 0 14304 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1677675658
transform -1 0 6336 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1677675658
transform -1 0 11424 0 1 3780
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1676385511
transform 1 0 576 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676385511
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676385511
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676385511
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676385511
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676385511
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676385511
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676385511
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676385511
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676385511
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676385511
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676385511
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676385511
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676385511
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676385511
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676385511
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676385511
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676385511
transform -1 0 960 0 1 8316
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via1 49968 38556 49968 38556 0 VGND
rlabel metal1 49968 37800 49968 37800 0 VPWR
rlabel metal3 12240 14196 12240 14196 0 _00_
rlabel metal3 10944 11172 10944 11172 0 _01_
rlabel metal3 8640 16464 8640 16464 0 _02_
rlabel metal2 3408 21000 3408 21000 0 _03_
rlabel metal2 4512 12264 4512 12264 0 _04_
rlabel metal2 9216 3738 9216 3738 0 _05_
rlabel metal2 4800 4410 4800 4410 0 _06_
rlabel metal2 10464 8064 10464 8064 0 _07_
rlabel metal3 8688 7980 8688 7980 0 _08_
rlabel metal2 4224 9828 4224 9828 0 _09_
rlabel metal2 5280 6048 5280 6048 0 _10_
rlabel via1 9293 7980 9293 7980 0 _11_
rlabel metal2 10368 13062 10368 13062 0 _12_
rlabel metal3 10800 13188 10800 13188 0 _13_
rlabel metal2 10848 11760 10848 11760 0 _14_
rlabel metal2 8544 11802 8544 11802 0 _15_
rlabel metal3 8688 16044 8688 16044 0 _16_
rlabel metal3 3072 20748 3072 20748 0 _17_
rlabel metal2 3456 11760 3456 11760 0 _18_
rlabel metal2 9264 4116 9264 4116 0 _19_
rlabel metal3 4512 5124 4512 5124 0 _20_
rlabel metal3 5280 7392 5280 7392 0 _21_
rlabel metal2 4656 4956 4656 4956 0 _22_
rlabel metal2 9888 12726 9888 12726 0 clk
rlabel metal2 11328 10710 11328 10710 0 clknet_0_clk
rlabel metal2 10464 3024 10464 3024 0 clknet_1_0__leaf_clk
rlabel metal2 8928 19656 8928 19656 0 clknet_1_1__leaf_clk
rlabel metal3 4416 13356 4416 13356 0 net
rlabel metal2 2784 20832 2784 20832 0 net1
rlabel metal2 864 15330 864 15330 0 net10
rlabel metal2 864 2730 864 2730 0 net11
rlabel metal2 912 3360 912 3360 0 net12
rlabel metal2 864 4242 864 4242 0 net13
rlabel metal2 864 4830 864 4830 0 net14
rlabel metal2 864 5964 864 5964 0 net15
rlabel metal2 816 7224 816 7224 0 net16
rlabel metal2 912 7896 912 7896 0 net17
rlabel metal3 1776 8736 1776 8736 0 net18
rlabel metal2 4080 3276 4080 3276 0 net19
rlabel metal3 1728 20748 1728 20748 0 net2
rlabel metal2 5376 21252 5376 21252 0 net20
rlabel metal2 12096 7170 12096 7170 0 net21
rlabel metal2 8064 17502 8064 17502 0 net22
rlabel metal2 9696 3108 9696 3108 0 net23
rlabel metal2 14544 10332 14544 10332 0 net24
rlabel metal2 13584 15372 13584 15372 0 net25
rlabel metal3 366 15708 366 15708 0 net26
rlabel metal3 366 16548 366 16548 0 net27
rlabel metal3 366 17388 366 17388 0 net28
rlabel metal3 366 18228 366 18228 0 net29
rlabel metal2 2832 2688 2832 2688 0 net3
rlabel metal3 366 19068 366 19068 0 net30
rlabel metal3 366 19908 366 19908 0 net31
rlabel metal3 366 20748 366 20748 0 net32
rlabel metal3 366 21588 366 21588 0 net33
rlabel metal2 2976 12348 2976 12348 0 net34
rlabel metal2 4224 11676 4224 11676 0 net35
rlabel metal2 9216 16506 9216 16506 0 net36
rlabel metal2 8064 17892 8064 17892 0 net37
rlabel metal3 11712 11676 11712 11676 0 net38
rlabel metal2 9888 10920 9888 10920 0 net39
rlabel metal3 1824 10248 1824 10248 0 net4
rlabel metal2 14064 11088 14064 11088 0 net40
rlabel metal2 5616 7140 5616 7140 0 net41
rlabel metal2 4320 5040 4320 5040 0 net42
rlabel metal2 3648 3276 3648 3276 0 net43
rlabel metal2 7104 8274 7104 8274 0 net44
rlabel metal3 11424 7728 11424 7728 0 net45
rlabel metal3 12384 14028 12384 14028 0 net46
rlabel metal3 4560 20748 4560 20748 0 net47
rlabel metal3 10080 4116 10080 4116 0 net48
rlabel metal2 3936 4662 3936 4662 0 net5
rlabel metal3 1968 4872 1968 4872 0 net6
rlabel metal3 2496 6384 2496 6384 0 net7
rlabel metal2 2496 11004 2496 11004 0 net8
rlabel metal2 2880 8820 2880 8820 0 net9
rlabel metal3 366 37548 366 37548 0 rst_n
rlabel metal3 318 22428 318 22428 0 ui_in[0]
rlabel metal3 366 8988 366 8988 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 366 10668 366 10668 0 uio_out[2]
rlabel metal3 366 11508 366 11508 0 uio_out[3]
rlabel metal3 366 12348 366 12348 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 366 14028 366 14028 0 uio_out[6]
rlabel metal3 366 14868 366 14868 0 uio_out[7]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 366 3948 366 3948 0 uo_out[2]
rlabel metal3 366 4788 366 4788 0 uo_out[3]
rlabel metal3 366 5628 366 5628 0 uo_out[4]
rlabel metal2 672 6720 672 6720 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
