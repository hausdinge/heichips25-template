VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc
  CLASS BLOCK ;
  FOREIGN adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 80.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 15.380 0.000 17.580 80.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.380 0.000 62.580 80.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 16.280 80.000 18.480 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 46.280 80.000 48.480 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 21.580 0.000 23.780 80.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.580 0.000 68.780 80.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 22.480 80.000 24.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 52.480 80.000 54.680 ;
    END
  END VSS
  PIN analog_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.020 0.400 38.420 ;
    END
  END analog_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 39.700 80.000 40.100 ;
    END
  END clk
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 37.180 80.000 37.580 ;
    END
  END data_out[0]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 41.560 0.000 41.960 0.400 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 38.860 80.000 39.260 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 38.020 80.000 38.420 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 39.640 0.000 40.040 0.400 ;
    END
  END data_out[7]
  PIN ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 40.540 80.000 40.940 ;
    END
  END ready
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.860 0.400 39.260 ;
    END
  END start
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 76.800 75.750 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 76.800 75.820 ;
      LAYER Metal2 ;
        RECT 3.255 0.610 79.305 75.745 ;
        RECT 3.255 0.400 38.470 0.610 ;
        RECT 39.290 0.400 39.430 0.610 ;
        RECT 40.250 0.400 40.390 0.610 ;
        RECT 41.210 0.400 41.350 0.610 ;
        RECT 42.170 0.400 42.310 0.610 ;
        RECT 43.130 0.400 79.305 0.610 ;
      LAYER Metal3 ;
        RECT 0.400 41.150 79.600 75.700 ;
        RECT 0.400 40.330 79.390 41.150 ;
        RECT 0.400 40.310 79.600 40.330 ;
        RECT 0.400 39.490 79.390 40.310 ;
        RECT 0.400 39.470 79.600 39.490 ;
        RECT 0.610 38.650 79.390 39.470 ;
        RECT 0.400 38.630 79.600 38.650 ;
        RECT 0.610 37.810 79.390 38.630 ;
        RECT 0.400 37.790 79.600 37.810 ;
        RECT 0.400 36.970 79.390 37.790 ;
        RECT 0.400 3.680 79.600 36.970 ;
  END
END adc
END LIBRARY

