* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_28_907 VPWR VGND sg13g2_decap_8
XFILLER_39_266 VPWR VGND sg13g2_decap_8
XFILLER_36_973 VPWR VGND sg13g2_decap_8
XFILLER_22_100 VPWR VGND sg13g2_decap_8
XFILLER_35_483 VPWR VGND sg13g2_decap_8
XFILLER_23_634 VPWR VGND sg13g2_decap_8
XFILLER_10_317 VPWR VGND sg13g2_decap_8
XFILLER_22_177 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_45_203 VPWR VGND sg13g2_decap_8
XFILLER_27_940 VPWR VGND sg13g2_decap_8
XFILLER_42_910 VPWR VGND sg13g2_decap_8
XFILLER_26_74 VPWR VGND sg13g2_decap_8
XFILLER_41_420 VPWR VGND sg13g2_decap_8
XFILLER_26_494 VPWR VGND sg13g2_decap_8
XFILLER_42_987 VPWR VGND sg13g2_decap_8
XFILLER_14_667 VPWR VGND sg13g2_decap_8
XFILLER_41_497 VPWR VGND sg13g2_decap_8
XFILLER_13_188 VPWR VGND sg13g2_decap_8
XFILLER_42_84 VPWR VGND sg13g2_decap_8
XFILLER_10_884 VPWR VGND sg13g2_decap_8
XFILLER_6_866 VPWR VGND sg13g2_decap_8
XFILLER_5_332 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_49_564 VPWR VGND sg13g2_decap_8
X_83_ net8 net16 VPWR VGND sg13g2_buf_1
XFILLER_36_203 VPWR VGND sg13g2_decap_8
XFILLER_18_962 VPWR VGND sg13g2_decap_8
XFILLER_45_770 VPWR VGND sg13g2_decap_8
XFILLER_17_472 VPWR VGND sg13g2_decap_8
XFILLER_33_910 VPWR VGND sg13g2_decap_8
XFILLER_44_280 VPWR VGND sg13g2_decap_8
XFILLER_32_420 VPWR VGND sg13g2_decap_8
XFILLER_33_987 VPWR VGND sg13g2_decap_8
XFILLER_20_637 VPWR VGND sg13g2_decap_8
XFILLER_32_497 VPWR VGND sg13g2_decap_8
XFILLER_9_671 VPWR VGND sg13g2_decap_8
XFILLER_8_170 VPWR VGND sg13g2_decap_8
XFILLER_28_704 VPWR VGND sg13g2_decap_8
XFILLER_43_707 VPWR VGND sg13g2_decap_8
XFILLER_27_247 VPWR VGND sg13g2_decap_8
XFILLER_42_217 VPWR VGND sg13g2_decap_8
XFILLER_24_921 VPWR VGND sg13g2_decap_8
XFILLER_36_770 VPWR VGND sg13g2_decap_8
XFILLER_23_431 VPWR VGND sg13g2_decap_8
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_24_998 VPWR VGND sg13g2_decap_8
XFILLER_10_114 VPWR VGND sg13g2_decap_8
XFILLER_11_637 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_3_858 VPWR VGND sg13g2_decap_8
XFILLER_2_357 VPWR VGND sg13g2_decap_8
XFILLER_19_748 VPWR VGND sg13g2_decap_8
XFILLER_46_567 VPWR VGND sg13g2_decap_8
XFILLER_34_707 VPWR VGND sg13g2_decap_8
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_18_269 VPWR VGND sg13g2_decap_8
XFILLER_33_217 VPWR VGND sg13g2_decap_8
XFILLER_15_932 VPWR VGND sg13g2_decap_8
XFILLER_18_1004 VPWR VGND sg13g2_decap_8
XFILLER_26_291 VPWR VGND sg13g2_decap_8
XFILLER_14_464 VPWR VGND sg13g2_decap_8
XFILLER_30_924 VPWR VGND sg13g2_decap_8
XFILLER_42_784 VPWR VGND sg13g2_decap_8
XFILLER_41_294 VPWR VGND sg13g2_decap_8
XFILLER_10_681 VPWR VGND sg13g2_decap_8
XFILLER_6_663 VPWR VGND sg13g2_decap_8
XFILLER_25_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_37_567 VPWR VGND sg13g2_decap_8
XFILLER_25_718 VPWR VGND sg13g2_decap_8
XFILLER_24_228 VPWR VGND sg13g2_decap_8
XFILLER_21_913 VPWR VGND sg13g2_decap_8
XFILLER_33_784 VPWR VGND sg13g2_decap_8
XFILLER_20_434 VPWR VGND sg13g2_decap_8
XFILLER_32_294 VPWR VGND sg13g2_decap_8
XFILLER_28_501 VPWR VGND sg13g2_decap_8
XFILLER_43_504 VPWR VGND sg13g2_decap_8
XFILLER_28_578 VPWR VGND sg13g2_decap_8
XFILLER_15_239 VPWR VGND sg13g2_decap_8
XFILLER_24_795 VPWR VGND sg13g2_decap_8
XFILLER_11_434 VPWR VGND sg13g2_decap_8
XFILLER_12_968 VPWR VGND sg13g2_decap_8
XFILLER_23_53 VPWR VGND sg13g2_decap_8
XFILLER_48_1008 VPWR VGND sg13g2_decap_8
XFILLER_3_655 VPWR VGND sg13g2_decap_8
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_545 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_34_504 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_42_581 VPWR VGND sg13g2_decap_8
XFILLER_14_261 VPWR VGND sg13g2_decap_8
XFILLER_30_721 VPWR VGND sg13g2_decap_8
XFILLER_9_99 VPWR VGND sg13g2_fill_2
XFILLER_30_798 VPWR VGND sg13g2_decap_8
XFILLER_31_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_950 VPWR VGND sg13g2_decap_8
XFILLER_6_460 VPWR VGND sg13g2_decap_8
XFILLER_38_854 VPWR VGND sg13g2_decap_8
X_49_ VGND VPWR net5 _10_ _20_ net41 sg13g2_a21oi_1
XFILLER_25_515 VPWR VGND sg13g2_decap_8
XFILLER_37_364 VPWR VGND sg13g2_decap_8
XFILLER_40_518 VPWR VGND sg13g2_decap_8
XFILLER_21_710 VPWR VGND sg13g2_decap_8
XFILLER_33_581 VPWR VGND sg13g2_decap_8
XFILLER_20_231 VPWR VGND sg13g2_decap_8
XFILLER_21_787 VPWR VGND sg13g2_decap_8
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_29_865 VPWR VGND sg13g2_decap_8
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_28_375 VPWR VGND sg13g2_decap_8
XFILLER_44_868 VPWR VGND sg13g2_decap_8
XFILLER_16_559 VPWR VGND sg13g2_decap_8
XFILLER_31_518 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_34_63 VPWR VGND sg13g2_decap_8
XFILLER_11_231 VPWR VGND sg13g2_decap_8
XFILLER_12_765 VPWR VGND sg13g2_decap_8
XFILLER_24_592 VPWR VGND sg13g2_decap_8
XFILLER_8_758 VPWR VGND sg13g2_decap_8
XFILLER_7_257 VPWR VGND sg13g2_decap_8
XFILLER_4_953 VPWR VGND sg13g2_decap_8
XFILLER_3_452 VPWR VGND sg13g2_decap_8
XFILLER_47_651 VPWR VGND sg13g2_decap_8
XFILLER_19_342 VPWR VGND sg13g2_decap_8
XFILLER_46_161 VPWR VGND sg13g2_decap_8
XFILLER_34_301 VPWR VGND sg13g2_decap_8
XFILLER_35_868 VPWR VGND sg13g2_decap_8
XFILLER_34_378 VPWR VGND sg13g2_decap_8
XFILLER_30_595 VPWR VGND sg13g2_decap_8
XFILLER_26_802 VPWR VGND sg13g2_decap_8
XFILLER_38_651 VPWR VGND sg13g2_decap_8
XFILLER_25_312 VPWR VGND sg13g2_decap_8
XFILLER_37_161 VPWR VGND sg13g2_decap_8
XFILLER_41_805 VPWR VGND sg13g2_decap_8
XFILLER_26_879 VPWR VGND sg13g2_decap_8
XFILLER_25_389 VPWR VGND sg13g2_decap_8
XFILLER_40_315 VPWR VGND sg13g2_decap_8
XFILLER_21_584 VPWR VGND sg13g2_decap_8
XFILLER_5_717 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_1_945 VPWR VGND sg13g2_decap_8
XFILLER_20_98 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_49_949 VPWR VGND sg13g2_decap_8
Xhold41 net6 VPWR VGND net41 sg13g2_dlygate4sd3_1
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_21_1011 VPWR VGND sg13g2_decap_8
XFILLER_29_74 VPWR VGND sg13g2_decap_8
XFILLER_29_662 VPWR VGND sg13g2_decap_8
XFILLER_17_857 VPWR VGND sg13g2_decap_8
XFILLER_28_172 VPWR VGND sg13g2_decap_8
XFILLER_44_665 VPWR VGND sg13g2_decap_8
XFILLER_16_356 VPWR VGND sg13g2_decap_8
XFILLER_32_805 VPWR VGND sg13g2_decap_8
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_43_175 VPWR VGND sg13g2_decap_8
XFILLER_31_315 VPWR VGND sg13g2_decap_8
XFILLER_12_562 VPWR VGND sg13g2_decap_8
XFILLER_40_882 VPWR VGND sg13g2_decap_8
XFILLER_8_555 VPWR VGND sg13g2_decap_8
XFILLER_6_89 VPWR VGND sg13g2_decap_8
XFILLER_4_750 VPWR VGND sg13g2_decap_8
XFILLER_6_1027 VPWR VGND sg13g2_fill_2
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_39_448 VPWR VGND sg13g2_decap_8
XFILLER_26_109 VPWR VGND sg13g2_decap_8
XFILLER_35_665 VPWR VGND sg13g2_decap_8
XFILLER_23_816 VPWR VGND sg13g2_decap_8
XFILLER_34_175 VPWR VGND sg13g2_decap_8
XFILLER_22_359 VPWR VGND sg13g2_decap_8
XFILLER_31_882 VPWR VGND sg13g2_decap_8
XFILLER_30_392 VPWR VGND sg13g2_decap_8
XFILLER_44_1022 VPWR VGND sg13g2_decap_8
Xheichips25_template_32 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_41_602 VPWR VGND sg13g2_decap_8
XFILLER_14_849 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_26_676 VPWR VGND sg13g2_decap_8
XFILLER_25_186 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_41_679 VPWR VGND sg13g2_decap_8
XFILLER_21_381 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_5_514 VPWR VGND sg13g2_decap_8
XFILLER_31_42 VPWR VGND sg13g2_decap_8
Xoutput7 net7 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_742 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_49_746 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_45_952 VPWR VGND sg13g2_decap_8
XFILLER_17_654 VPWR VGND sg13g2_decap_8
XFILLER_44_462 VPWR VGND sg13g2_decap_8
XFILLER_16_153 VPWR VGND sg13g2_decap_8
XFILLER_32_602 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_decap_8
XFILLER_13_860 VPWR VGND sg13g2_decap_8
XFILLER_20_819 VPWR VGND sg13g2_decap_8
XFILLER_32_679 VPWR VGND sg13g2_decap_8
XFILLER_9_853 VPWR VGND sg13g2_decap_8
XFILLER_31_189 VPWR VGND sg13g2_decap_8
XFILLER_8_352 VPWR VGND sg13g2_decap_8
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_245 VPWR VGND sg13g2_decap_8
XFILLER_27_429 VPWR VGND sg13g2_decap_8
XFILLER_36_952 VPWR VGND sg13g2_decap_8
XFILLER_23_613 VPWR VGND sg13g2_decap_8
XFILLER_35_462 VPWR VGND sg13g2_decap_8
XFILLER_11_819 VPWR VGND sg13g2_decap_8
XFILLER_22_156 VPWR VGND sg13g2_decap_8
XFILLER_2_539 VPWR VGND sg13g2_decap_8
XFILLER_46_749 VPWR VGND sg13g2_decap_8
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_26_473 VPWR VGND sg13g2_decap_8
XFILLER_27_996 VPWR VGND sg13g2_decap_8
XFILLER_42_966 VPWR VGND sg13g2_decap_8
XFILLER_14_646 VPWR VGND sg13g2_decap_8
XFILLER_41_476 VPWR VGND sg13g2_decap_8
XFILLER_13_134 VPWR VGND sg13g2_decap_4
XFILLER_13_167 VPWR VGND sg13g2_decap_8
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_10_863 VPWR VGND sg13g2_decap_8
XFILLER_6_845 VPWR VGND sg13g2_decap_8
XFILLER_5_311 VPWR VGND sg13g2_decap_8
XFILLER_5_388 VPWR VGND sg13g2_decap_8
XFILLER_3_68 VPWR VGND sg13g2_decap_8
XFILLER_49_543 VPWR VGND sg13g2_decap_8
X_82_ net7 net15 VPWR VGND sg13g2_buf_1
XFILLER_3_1019 VPWR VGND sg13g2_decap_8
XFILLER_37_749 VPWR VGND sg13g2_decap_8
XFILLER_18_941 VPWR VGND sg13g2_decap_8
XFILLER_36_259 VPWR VGND sg13g2_decap_8
XFILLER_17_451 VPWR VGND sg13g2_decap_8
XFILLER_20_616 VPWR VGND sg13g2_decap_8
XFILLER_33_966 VPWR VGND sg13g2_decap_8
XFILLER_32_476 VPWR VGND sg13g2_decap_8
XFILLER_9_650 VPWR VGND sg13g2_decap_8
XFILLER_27_226 VPWR VGND sg13g2_decap_8
XFILLER_24_900 VPWR VGND sg13g2_decap_8
XFILLER_23_410 VPWR VGND sg13g2_decap_8
XFILLER_24_977 VPWR VGND sg13g2_decap_8
XFILLER_11_616 VPWR VGND sg13g2_decap_8
XFILLER_23_487 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_12_88 VPWR VGND sg13g2_decap_8
XFILLER_3_837 VPWR VGND sg13g2_decap_8
XFILLER_2_336 VPWR VGND sg13g2_decap_8
XFILLER_19_727 VPWR VGND sg13g2_decap_8
XFILLER_46_546 VPWR VGND sg13g2_decap_8
XFILLER_18_248 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_15_911 VPWR VGND sg13g2_decap_8
XFILLER_26_270 VPWR VGND sg13g2_decap_8
XFILLER_27_793 VPWR VGND sg13g2_decap_8
XFILLER_42_763 VPWR VGND sg13g2_decap_8
XFILLER_14_443 VPWR VGND sg13g2_decap_8
XFILLER_15_988 VPWR VGND sg13g2_decap_8
XFILLER_30_903 VPWR VGND sg13g2_decap_8
XFILLER_41_273 VPWR VGND sg13g2_decap_8
XFILLER_10_660 VPWR VGND sg13g2_decap_8
XFILLER_6_642 VPWR VGND sg13g2_decap_8
XFILLER_5_185 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
XFILLER_37_546 VPWR VGND sg13g2_decap_8
XFILLER_24_207 VPWR VGND sg13g2_decap_8
XFILLER_33_763 VPWR VGND sg13g2_decap_8
XFILLER_20_413 VPWR VGND sg13g2_decap_8
XFILLER_32_273 VPWR VGND sg13g2_decap_8
XFILLER_21_969 VPWR VGND sg13g2_decap_8
XFILLER_28_557 VPWR VGND sg13g2_decap_8
XFILLER_15_218 VPWR VGND sg13g2_decap_8
XFILLER_11_413 VPWR VGND sg13g2_decap_8
XFILLER_12_947 VPWR VGND sg13g2_decap_8
XFILLER_24_774 VPWR VGND sg13g2_decap_8
XFILLER_23_32 VPWR VGND sg13g2_decap_8
XFILLER_23_284 VPWR VGND sg13g2_decap_8
XFILLER_7_439 VPWR VGND sg13g2_decap_8
XFILLER_20_980 VPWR VGND sg13g2_decap_8
XFILLER_3_634 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_decap_8
XFILLER_47_833 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_19_524 VPWR VGND sg13g2_decap_8
XFILLER_46_343 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_27_590 VPWR VGND sg13g2_decap_8
XFILLER_14_240 VPWR VGND sg13g2_decap_8
XFILLER_42_560 VPWR VGND sg13g2_decap_8
XFILLER_15_785 VPWR VGND sg13g2_decap_8
XFILLER_30_700 VPWR VGND sg13g2_decap_8
XFILLER_9_67 VPWR VGND sg13g2_decap_8
XFILLER_30_777 VPWR VGND sg13g2_decap_8
XFILLER_11_980 VPWR VGND sg13g2_decap_8
XFILLER_9_1014 VPWR VGND sg13g2_decap_8
XFILLER_38_833 VPWR VGND sg13g2_decap_8
X_48_ VGND VPWR net48 _10_ _05_ _19_ sg13g2_a21oi_1
XFILLER_37_343 VPWR VGND sg13g2_decap_8
XFILLER_33_560 VPWR VGND sg13g2_decap_8
XFILLER_20_210 VPWR VGND sg13g2_decap_8
XFILLER_21_766 VPWR VGND sg13g2_decap_8
XFILLER_20_287 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_29_844 VPWR VGND sg13g2_decap_8
XFILLER_28_354 VPWR VGND sg13g2_decap_8
XFILLER_44_847 VPWR VGND sg13g2_decap_8
XFILLER_16_538 VPWR VGND sg13g2_decap_8
XFILLER_43_357 VPWR VGND sg13g2_decap_8
XFILLER_24_571 VPWR VGND sg13g2_decap_8
XFILLER_34_42 VPWR VGND sg13g2_decap_8
XFILLER_11_210 VPWR VGND sg13g2_decap_8
XFILLER_12_744 VPWR VGND sg13g2_decap_8
XFILLER_8_737 VPWR VGND sg13g2_decap_8
XFILLER_7_236 VPWR VGND sg13g2_decap_8
XFILLER_11_287 VPWR VGND sg13g2_decap_8
XFILLER_4_932 VPWR VGND sg13g2_decap_8
XFILLER_3_431 VPWR VGND sg13g2_decap_8
XFILLER_47_630 VPWR VGND sg13g2_decap_8
XFILLER_19_321 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_19_398 VPWR VGND sg13g2_decap_8
XFILLER_35_847 VPWR VGND sg13g2_decap_8
XFILLER_34_357 VPWR VGND sg13g2_decap_8
XFILLER_15_582 VPWR VGND sg13g2_decap_8
XFILLER_30_574 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_38_630 VPWR VGND sg13g2_decap_8
XFILLER_37_140 VPWR VGND sg13g2_decap_8
XFILLER_26_858 VPWR VGND sg13g2_decap_8
XFILLER_38_1008 VPWR VGND sg13g2_decap_8
XFILLER_25_368 VPWR VGND sg13g2_decap_8
XFILLER_21_563 VPWR VGND sg13g2_decap_8
XFILLER_4_239 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_1_924 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_49_928 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_29_53 VPWR VGND sg13g2_decap_8
Xhold42 _20_ VPWR VGND net42 sg13g2_dlygate4sd3_1
XFILLER_29_641 VPWR VGND sg13g2_decap_8
XFILLER_17_836 VPWR VGND sg13g2_decap_8
XFILLER_28_151 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_8
XFILLER_44_644 VPWR VGND sg13g2_decap_8
XFILLER_16_335 VPWR VGND sg13g2_decap_8
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_12_541 VPWR VGND sg13g2_decap_8
XFILLER_40_861 VPWR VGND sg13g2_decap_8
XFILLER_8_534 VPWR VGND sg13g2_decap_8
XFILLER_6_68 VPWR VGND sg13g2_decap_8
XFILLER_6_1006 VPWR VGND sg13g2_decap_8
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_39_427 VPWR VGND sg13g2_decap_8
XFILLER_48_994 VPWR VGND sg13g2_decap_8
XFILLER_19_195 VPWR VGND sg13g2_decap_8
XFILLER_35_644 VPWR VGND sg13g2_decap_8
XFILLER_34_154 VPWR VGND sg13g2_decap_8
XFILLER_22_338 VPWR VGND sg13g2_decap_8
XFILLER_31_861 VPWR VGND sg13g2_decap_8
XFILLER_30_371 VPWR VGND sg13g2_decap_8
XFILLER_44_1001 VPWR VGND sg13g2_decap_8
Xheichips25_template_33 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_39_994 VPWR VGND sg13g2_decap_8
XFILLER_26_655 VPWR VGND sg13g2_decap_8
XFILLER_14_828 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_25_165 VPWR VGND sg13g2_decap_8
XFILLER_41_658 VPWR VGND sg13g2_decap_8
XFILLER_13_349 VPWR VGND sg13g2_decap_8
XFILLER_15_88 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
XFILLER_21_360 VPWR VGND sg13g2_decap_8
XFILLER_31_21 VPWR VGND sg13g2_decap_8
XFILLER_31_98 VPWR VGND sg13g2_decap_8
Xoutput8 net8 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_721 VPWR VGND sg13g2_decap_8
XFILLER_49_725 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_45_931 VPWR VGND sg13g2_decap_8
XFILLER_44_441 VPWR VGND sg13g2_decap_8
XFILLER_16_132 VPWR VGND sg13g2_decap_8
XFILLER_17_633 VPWR VGND sg13g2_decap_8
XFILLER_32_658 VPWR VGND sg13g2_decap_8
XFILLER_31_168 VPWR VGND sg13g2_decap_8
XFILLER_9_832 VPWR VGND sg13g2_decap_8
XFILLER_8_331 VPWR VGND sg13g2_decap_8
XFILLER_39_224 VPWR VGND sg13g2_decap_8
XFILLER_27_408 VPWR VGND sg13g2_decap_8
XFILLER_48_791 VPWR VGND sg13g2_decap_8
XFILLER_36_931 VPWR VGND sg13g2_decap_8
XFILLER_35_441 VPWR VGND sg13g2_decap_8
XFILLER_22_135 VPWR VGND sg13g2_decap_8
XFILLER_23_669 VPWR VGND sg13g2_decap_8
XFILLER_11_1022 VPWR VGND sg13g2_decap_8
XFILLER_2_518 VPWR VGND sg13g2_decap_8
XFILLER_19_909 VPWR VGND sg13g2_decap_8
XFILLER_46_728 VPWR VGND sg13g2_decap_8
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_39_791 VPWR VGND sg13g2_decap_8
XFILLER_26_452 VPWR VGND sg13g2_decap_8
XFILLER_27_975 VPWR VGND sg13g2_decap_8
XFILLER_42_945 VPWR VGND sg13g2_decap_8
XFILLER_13_113 VPWR VGND sg13g2_decap_8
XFILLER_14_625 VPWR VGND sg13g2_decap_8
XFILLER_41_455 VPWR VGND sg13g2_decap_8
XFILLER_42_42 VPWR VGND sg13g2_decap_8
XFILLER_9_139 VPWR VGND sg13g2_decap_8
XFILLER_10_842 VPWR VGND sg13g2_decap_8
XFILLER_6_824 VPWR VGND sg13g2_decap_8
XFILLER_5_367 VPWR VGND sg13g2_decap_8
XFILLER_3_47 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_8
X_81_ net6 net14 VPWR VGND sg13g2_buf_1
XFILLER_49_599 VPWR VGND sg13g2_decap_8
XFILLER_18_920 VPWR VGND sg13g2_decap_8
XFILLER_37_728 VPWR VGND sg13g2_decap_8
XFILLER_17_430 VPWR VGND sg13g2_decap_8
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_18_997 VPWR VGND sg13g2_decap_8
XFILLER_33_945 VPWR VGND sg13g2_decap_8
XFILLER_32_455 VPWR VGND sg13g2_decap_8
XFILLER_34_1022 VPWR VGND sg13g2_decap_8
XFILLER_41_1015 VPWR VGND sg13g2_decap_8
XFILLER_27_205 VPWR VGND sg13g2_decap_8
XFILLER_28_739 VPWR VGND sg13g2_decap_8
XFILLER_24_956 VPWR VGND sg13g2_decap_8
XFILLER_23_466 VPWR VGND sg13g2_decap_8
XFILLER_10_149 VPWR VGND sg13g2_decap_8
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_2_315 VPWR VGND sg13g2_decap_8
XFILLER_19_706 VPWR VGND sg13g2_decap_8
XFILLER_46_525 VPWR VGND sg13g2_decap_8
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_18_227 VPWR VGND sg13g2_decap_8
XFILLER_27_772 VPWR VGND sg13g2_decap_8
XFILLER_14_422 VPWR VGND sg13g2_decap_8
XFILLER_42_742 VPWR VGND sg13g2_decap_8
XFILLER_15_967 VPWR VGND sg13g2_decap_8
XFILLER_14_499 VPWR VGND sg13g2_decap_8
XFILLER_41_252 VPWR VGND sg13g2_decap_8
XFILLER_30_959 VPWR VGND sg13g2_decap_8
XFILLER_6_621 VPWR VGND sg13g2_decap_8
XFILLER_5_164 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_6_698 VPWR VGND sg13g2_decap_8
XFILLER_2_882 VPWR VGND sg13g2_decap_8
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_37_525 VPWR VGND sg13g2_decap_8
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_18_794 VPWR VGND sg13g2_decap_8
XFILLER_33_742 VPWR VGND sg13g2_decap_8
XFILLER_21_948 VPWR VGND sg13g2_decap_8
XFILLER_32_252 VPWR VGND sg13g2_decap_8
XFILLER_20_469 VPWR VGND sg13g2_decap_8
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_28_536 VPWR VGND sg13g2_decap_8
XFILLER_43_539 VPWR VGND sg13g2_decap_8
XFILLER_24_753 VPWR VGND sg13g2_decap_8
XFILLER_12_926 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_23_263 VPWR VGND sg13g2_decap_8
XFILLER_8_919 VPWR VGND sg13g2_decap_8
XFILLER_7_418 VPWR VGND sg13g2_decap_8
XFILLER_11_469 VPWR VGND sg13g2_decap_8
XFILLER_23_88 VPWR VGND sg13g2_decap_8
XFILLER_3_613 VPWR VGND sg13g2_decap_8
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_47_812 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_19_503 VPWR VGND sg13g2_decap_8
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_47_889 VPWR VGND sg13g2_decap_8
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_34_539 VPWR VGND sg13g2_decap_8
XFILLER_15_764 VPWR VGND sg13g2_decap_8
XFILLER_9_46 VPWR VGND sg13g2_decap_8
XFILLER_14_296 VPWR VGND sg13g2_decap_8
XFILLER_30_756 VPWR VGND sg13g2_decap_8
XFILLER_7_985 VPWR VGND sg13g2_decap_8
XFILLER_6_495 VPWR VGND sg13g2_decap_8
XFILLER_38_812 VPWR VGND sg13g2_decap_8
XFILLER_49_193 VPWR VGND sg13g2_decap_8
XFILLER_37_322 VPWR VGND sg13g2_decap_8
X_47_ net1 VPWR _19_ VGND net48 _10_ sg13g2_o21ai_1
XFILLER_38_889 VPWR VGND sg13g2_decap_8
XFILLER_37_399 VPWR VGND sg13g2_decap_8
XFILLER_18_591 VPWR VGND sg13g2_decap_8
XFILLER_21_745 VPWR VGND sg13g2_decap_8
XFILLER_20_266 VPWR VGND sg13g2_decap_8
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_48_609 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_29_823 VPWR VGND sg13g2_decap_8
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_28_333 VPWR VGND sg13g2_decap_8
XFILLER_44_826 VPWR VGND sg13g2_decap_8
XFILLER_16_517 VPWR VGND sg13g2_decap_8
XFILLER_18_88 VPWR VGND sg13g2_decap_8
XFILLER_43_336 VPWR VGND sg13g2_decap_8
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_24_550 VPWR VGND sg13g2_decap_8
XFILLER_12_723 VPWR VGND sg13g2_decap_8
XFILLER_15_1009 VPWR VGND sg13g2_decap_8
XFILLER_34_98 VPWR VGND sg13g2_decap_8
XFILLER_8_716 VPWR VGND sg13g2_decap_8
XFILLER_11_266 VPWR VGND sg13g2_decap_8
XFILLER_7_215 VPWR VGND sg13g2_decap_8
XFILLER_4_911 VPWR VGND sg13g2_decap_8
XFILLER_3_410 VPWR VGND sg13g2_decap_8
XFILLER_4_988 VPWR VGND sg13g2_decap_8
XFILLER_3_487 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_39_609 VPWR VGND sg13g2_decap_8
XFILLER_38_119 VPWR VGND sg13g2_decap_8
XFILLER_19_300 VPWR VGND sg13g2_decap_8
XFILLER_47_686 VPWR VGND sg13g2_decap_8
XFILLER_19_377 VPWR VGND sg13g2_decap_8
XFILLER_35_826 VPWR VGND sg13g2_decap_8
XFILLER_46_196 VPWR VGND sg13g2_decap_8
XFILLER_34_336 VPWR VGND sg13g2_decap_8
XFILLER_15_561 VPWR VGND sg13g2_decap_8
XFILLER_30_553 VPWR VGND sg13g2_decap_8
XFILLER_7_782 VPWR VGND sg13g2_decap_8
XFILLER_6_292 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_26_837 VPWR VGND sg13g2_decap_8
XFILLER_38_686 VPWR VGND sg13g2_decap_8
XFILLER_25_347 VPWR VGND sg13g2_decap_8
XFILLER_37_196 VPWR VGND sg13g2_decap_8
XFILLER_21_542 VPWR VGND sg13g2_decap_8
XFILLER_4_218 VPWR VGND sg13g2_decap_8
XFILLER_1_903 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_49_907 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_29_32 VPWR VGND sg13g2_decap_8
Xhold43 _06_ VPWR VGND net43 sg13g2_dlygate4sd3_1
XFILLER_29_620 VPWR VGND sg13g2_decap_8
XFILLER_28_130 VPWR VGND sg13g2_decap_8
XFILLER_44_623 VPWR VGND sg13g2_decap_8
XFILLER_16_314 VPWR VGND sg13g2_decap_8
XFILLER_17_815 VPWR VGND sg13g2_decap_8
XFILLER_29_697 VPWR VGND sg13g2_decap_8
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_43_133 VPWR VGND sg13g2_decap_8
XFILLER_12_520 VPWR VGND sg13g2_decap_8
XFILLER_8_513 VPWR VGND sg13g2_decap_8
XFILLER_40_840 VPWR VGND sg13g2_decap_8
XFILLER_12_597 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
XFILLER_6_47 VPWR VGND sg13g2_decap_8
XFILLER_6_36 VPWR VGND sg13g2_fill_2
XFILLER_4_785 VPWR VGND sg13g2_decap_8
XFILLER_3_284 VPWR VGND sg13g2_decap_8
XFILLER_39_406 VPWR VGND sg13g2_decap_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
XFILLER_48_973 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
XFILLER_19_174 VPWR VGND sg13g2_decap_8
XFILLER_35_623 VPWR VGND sg13g2_decap_8
XFILLER_34_133 VPWR VGND sg13g2_decap_8
XFILLER_16_881 VPWR VGND sg13g2_decap_8
XFILLER_22_317 VPWR VGND sg13g2_decap_8
XFILLER_31_840 VPWR VGND sg13g2_decap_8
XFILLER_30_350 VPWR VGND sg13g2_decap_8
XFILLER_39_973 VPWR VGND sg13g2_decap_8
XFILLER_38_483 VPWR VGND sg13g2_decap_8
XFILLER_26_634 VPWR VGND sg13g2_decap_8
XFILLER_14_807 VPWR VGND sg13g2_decap_8
XFILLER_25_144 VPWR VGND sg13g2_decap_8
XFILLER_41_637 VPWR VGND sg13g2_decap_8
XFILLER_13_328 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_22_884 VPWR VGND sg13g2_decap_8
XFILLER_31_77 VPWR VGND sg13g2_decap_8
XFILLER_5_549 VPWR VGND sg13g2_decap_8
XFILLER_1_700 VPWR VGND sg13g2_decap_8
Xoutput11 net11 uo_out[0] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_49_704 VPWR VGND sg13g2_decap_8
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_45_910 VPWR VGND sg13g2_decap_8
XFILLER_17_612 VPWR VGND sg13g2_decap_8
XFILLER_44_420 VPWR VGND sg13g2_decap_8
XFILLER_16_111 VPWR VGND sg13g2_decap_8
XFILLER_29_494 VPWR VGND sg13g2_decap_8
XFILLER_45_987 VPWR VGND sg13g2_decap_8
XFILLER_17_689 VPWR VGND sg13g2_decap_8
XFILLER_44_497 VPWR VGND sg13g2_decap_8
XFILLER_16_188 VPWR VGND sg13g2_decap_8
XFILLER_32_637 VPWR VGND sg13g2_decap_8
XFILLER_9_811 VPWR VGND sg13g2_decap_8
XFILLER_31_147 VPWR VGND sg13g2_decap_8
XFILLER_8_310 VPWR VGND sg13g2_decap_8
XFILLER_13_895 VPWR VGND sg13g2_decap_8
XFILLER_9_888 VPWR VGND sg13g2_decap_8
XFILLER_12_394 VPWR VGND sg13g2_decap_8
XFILLER_8_387 VPWR VGND sg13g2_decap_8
XFILLER_4_582 VPWR VGND sg13g2_decap_8
XFILLER_28_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_203 VPWR VGND sg13g2_decap_8
XFILLER_48_770 VPWR VGND sg13g2_decap_8
XFILLER_36_910 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_decap_8
XFILLER_35_420 VPWR VGND sg13g2_decap_8
XFILLER_36_987 VPWR VGND sg13g2_decap_8
XFILLER_22_114 VPWR VGND sg13g2_decap_8
XFILLER_23_648 VPWR VGND sg13g2_decap_8
XFILLER_35_497 VPWR VGND sg13g2_decap_8
XFILLER_11_1001 VPWR VGND sg13g2_decap_8
XFILLER_46_707 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_18_409 VPWR VGND sg13g2_decap_8
XFILLER_39_770 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_26_431 VPWR VGND sg13g2_decap_8
XFILLER_27_954 VPWR VGND sg13g2_decap_8
XFILLER_38_280 VPWR VGND sg13g2_decap_8
XFILLER_14_604 VPWR VGND sg13g2_decap_8
XFILLER_42_924 VPWR VGND sg13g2_decap_8
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_41_434 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_10_821 VPWR VGND sg13g2_decap_8
XFILLER_6_803 VPWR VGND sg13g2_decap_8
XFILLER_22_681 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_5_346 VPWR VGND sg13g2_decap_8
XFILLER_10_898 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
X_80_ net5 net13 VPWR VGND sg13g2_buf_1
XFILLER_37_707 VPWR VGND sg13g2_decap_8
XFILLER_49_578 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_29_291 VPWR VGND sg13g2_decap_8
XFILLER_18_976 VPWR VGND sg13g2_decap_8
XFILLER_45_784 VPWR VGND sg13g2_decap_8
XFILLER_17_486 VPWR VGND sg13g2_decap_8
XFILLER_33_924 VPWR VGND sg13g2_decap_8
XFILLER_44_294 VPWR VGND sg13g2_decap_8
XFILLER_32_434 VPWR VGND sg13g2_decap_8
XFILLER_34_1001 VPWR VGND sg13g2_decap_8
XFILLER_13_692 VPWR VGND sg13g2_decap_8
XFILLER_9_685 VPWR VGND sg13g2_decap_8
XFILLER_12_191 VPWR VGND sg13g2_decap_8
XFILLER_8_184 VPWR VGND sg13g2_decap_8
XFILLER_28_718 VPWR VGND sg13g2_decap_8
XFILLER_24_935 VPWR VGND sg13g2_decap_8
XFILLER_36_784 VPWR VGND sg13g2_decap_8
XFILLER_23_445 VPWR VGND sg13g2_decap_8
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_10_128 VPWR VGND sg13g2_decap_8
XFILLER_12_46 VPWR VGND sg13g2_decap_8
XFILLER_46_504 VPWR VGND sg13g2_decap_8
XFILLER_18_206 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_27_751 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_42_721 VPWR VGND sg13g2_decap_8
XFILLER_14_401 VPWR VGND sg13g2_decap_8
XFILLER_15_946 VPWR VGND sg13g2_decap_8
XFILLER_18_1018 VPWR VGND sg13g2_decap_8
XFILLER_41_231 VPWR VGND sg13g2_decap_8
XFILLER_42_798 VPWR VGND sg13g2_decap_8
XFILLER_14_478 VPWR VGND sg13g2_decap_8
XFILLER_30_938 VPWR VGND sg13g2_decap_8
XFILLER_6_600 VPWR VGND sg13g2_decap_8
XFILLER_10_695 VPWR VGND sg13g2_decap_8
XFILLER_6_677 VPWR VGND sg13g2_decap_8
XFILLER_5_143 VPWR VGND sg13g2_decap_8
XFILLER_2_861 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_37_504 VPWR VGND sg13g2_decap_8
XFILLER_45_581 VPWR VGND sg13g2_decap_8
XFILLER_18_773 VPWR VGND sg13g2_decap_8
XFILLER_33_721 VPWR VGND sg13g2_decap_8
XFILLER_17_283 VPWR VGND sg13g2_decap_8
XFILLER_32_231 VPWR VGND sg13g2_decap_8
XFILLER_21_927 VPWR VGND sg13g2_decap_8
XFILLER_33_798 VPWR VGND sg13g2_decap_8
XFILLER_20_448 VPWR VGND sg13g2_decap_8
XFILLER_9_482 VPWR VGND sg13g2_decap_8
XFILLER_28_515 VPWR VGND sg13g2_decap_8
XFILLER_43_518 VPWR VGND sg13g2_decap_8
XFILLER_36_581 VPWR VGND sg13g2_decap_8
XFILLER_12_905 VPWR VGND sg13g2_decap_8
XFILLER_24_732 VPWR VGND sg13g2_decap_8
XFILLER_23_242 VPWR VGND sg13g2_decap_8
XFILLER_11_448 VPWR VGND sg13g2_decap_8
XFILLER_23_67 VPWR VGND sg13g2_decap_8
XFILLER_3_669 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_19_559 VPWR VGND sg13g2_decap_8
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_34_518 VPWR VGND sg13g2_decap_8
XFILLER_15_743 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_decap_8
XFILLER_42_595 VPWR VGND sg13g2_decap_8
XFILLER_14_275 VPWR VGND sg13g2_decap_8
XFILLER_30_735 VPWR VGND sg13g2_decap_8
XFILLER_31_1015 VPWR VGND sg13g2_decap_8
XFILLER_10_492 VPWR VGND sg13g2_decap_8
XFILLER_7_964 VPWR VGND sg13g2_decap_8
XFILLER_6_474 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_37_301 VPWR VGND sg13g2_decap_8
X_46_ _09_ _10_ net35 _04_ VPWR VGND sg13g2_nor3_1
XFILLER_38_868 VPWR VGND sg13g2_decap_8
XFILLER_18_570 VPWR VGND sg13g2_decap_8
XFILLER_25_529 VPWR VGND sg13g2_decap_8
XFILLER_37_378 VPWR VGND sg13g2_decap_8
XFILLER_21_724 VPWR VGND sg13g2_decap_8
XFILLER_33_595 VPWR VGND sg13g2_decap_8
XFILLER_20_245 VPWR VGND sg13g2_decap_8
XFILLER_47_1022 VPWR VGND sg13g2_decap_8
XFILLER_29_802 VPWR VGND sg13g2_decap_8
XFILLER_28_312 VPWR VGND sg13g2_decap_8
XFILLER_44_805 VPWR VGND sg13g2_decap_8
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_29_879 VPWR VGND sg13g2_decap_8
XFILLER_43_315 VPWR VGND sg13g2_decap_8
XFILLER_28_389 VPWR VGND sg13g2_decap_8
XFILLER_12_702 VPWR VGND sg13g2_decap_8
XFILLER_34_77 VPWR VGND sg13g2_decap_8
XFILLER_11_245 VPWR VGND sg13g2_decap_8
XFILLER_12_779 VPWR VGND sg13g2_decap_8
XFILLER_4_967 VPWR VGND sg13g2_decap_8
XFILLER_3_466 VPWR VGND sg13g2_decap_8
XFILLER_47_665 VPWR VGND sg13g2_decap_8
XFILLER_19_356 VPWR VGND sg13g2_decap_8
XFILLER_35_805 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_34_315 VPWR VGND sg13g2_decap_8
XFILLER_15_540 VPWR VGND sg13g2_decap_8
XFILLER_43_882 VPWR VGND sg13g2_decap_8
XFILLER_42_392 VPWR VGND sg13g2_decap_8
XFILLER_30_532 VPWR VGND sg13g2_decap_8
XFILLER_7_761 VPWR VGND sg13g2_decap_8
XFILLER_6_271 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_29_109 VPWR VGND sg13g2_decap_8
XFILLER_38_665 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_26_816 VPWR VGND sg13g2_decap_8
XFILLER_37_175 VPWR VGND sg13g2_decap_8
XFILLER_25_326 VPWR VGND sg13g2_decap_8
XFILLER_41_819 VPWR VGND sg13g2_decap_8
XFILLER_21_521 VPWR VGND sg13g2_decap_8
XFILLER_34_882 VPWR VGND sg13g2_decap_8
XFILLER_40_329 VPWR VGND sg13g2_decap_8
XFILLER_33_392 VPWR VGND sg13g2_decap_8
XFILLER_14_1010 VPWR VGND sg13g2_decap_8
XFILLER_21_598 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_1_959 VPWR VGND sg13g2_decap_8
XFILLER_29_11 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
Xhold44 net7 VPWR VGND net44 sg13g2_dlygate4sd3_1
XFILLER_21_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_88 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_44_602 VPWR VGND sg13g2_decap_8
XFILLER_29_676 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_28_186 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_44_679 VPWR VGND sg13g2_decap_8
XFILLER_32_819 VPWR VGND sg13g2_decap_8
XFILLER_43_189 VPWR VGND sg13g2_decap_8
XFILLER_25_893 VPWR VGND sg13g2_decap_8
XFILLER_31_329 VPWR VGND sg13g2_decap_8
XFILLER_12_576 VPWR VGND sg13g2_decap_8
XFILLER_40_896 VPWR VGND sg13g2_decap_8
XFILLER_8_569 VPWR VGND sg13g2_decap_8
XFILLER_4_764 VPWR VGND sg13g2_decap_8
XFILLER_3_263 VPWR VGND sg13g2_decap_8
XFILLER_48_952 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_19_153 VPWR VGND sg13g2_decap_8
XFILLER_35_602 VPWR VGND sg13g2_decap_8
XFILLER_34_112 VPWR VGND sg13g2_decap_8
XFILLER_16_860 VPWR VGND sg13g2_decap_8
XFILLER_35_679 VPWR VGND sg13g2_decap_8
XFILLER_34_189 VPWR VGND sg13g2_decap_8
XFILLER_31_896 VPWR VGND sg13g2_decap_8
XFILLER_39_952 VPWR VGND sg13g2_decap_8
XFILLER_26_613 VPWR VGND sg13g2_decap_8
XFILLER_38_462 VPWR VGND sg13g2_decap_8
XFILLER_25_123 VPWR VGND sg13g2_decap_8
XFILLER_41_616 VPWR VGND sg13g2_decap_8
XFILLER_13_307 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_22_863 VPWR VGND sg13g2_decap_8
XFILLER_21_395 VPWR VGND sg13g2_decap_8
XFILLER_5_528 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_decap_8
Xoutput12 net12 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_756 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_29_473 VPWR VGND sg13g2_decap_8
XFILLER_45_966 VPWR VGND sg13g2_decap_8
XFILLER_17_668 VPWR VGND sg13g2_decap_8
XFILLER_44_476 VPWR VGND sg13g2_decap_8
XFILLER_16_167 VPWR VGND sg13g2_decap_8
XFILLER_32_616 VPWR VGND sg13g2_decap_8
XFILLER_25_690 VPWR VGND sg13g2_decap_8
XFILLER_31_126 VPWR VGND sg13g2_decap_8
XFILLER_13_874 VPWR VGND sg13g2_decap_8
XFILLER_9_867 VPWR VGND sg13g2_decap_8
XFILLER_12_373 VPWR VGND sg13g2_decap_8
XFILLER_40_693 VPWR VGND sg13g2_decap_8
XFILLER_8_366 VPWR VGND sg13g2_decap_8
XFILLER_4_561 VPWR VGND sg13g2_decap_8
XFILLER_39_259 VPWR VGND sg13g2_decap_8
XFILLER_36_966 VPWR VGND sg13g2_decap_8
XFILLER_23_627 VPWR VGND sg13g2_decap_8
XFILLER_35_476 VPWR VGND sg13g2_decap_8
XFILLER_31_693 VPWR VGND sg13g2_decap_8
XFILLER_26_410 VPWR VGND sg13g2_decap_8
XFILLER_27_933 VPWR VGND sg13g2_decap_8
XFILLER_42_903 VPWR VGND sg13g2_decap_8
XFILLER_41_413 VPWR VGND sg13g2_decap_8
XFILLER_26_67 VPWR VGND sg13g2_decap_8
XFILLER_26_487 VPWR VGND sg13g2_decap_8
XFILLER_10_800 VPWR VGND sg13g2_decap_8
XFILLER_22_660 VPWR VGND sg13g2_decap_8
XFILLER_42_77 VPWR VGND sg13g2_decap_8
XFILLER_10_877 VPWR VGND sg13g2_decap_8
XFILLER_21_192 VPWR VGND sg13g2_decap_8
XFILLER_6_859 VPWR VGND sg13g2_decap_8
XFILLER_5_325 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_18_955 VPWR VGND sg13g2_decap_8
XFILLER_29_270 VPWR VGND sg13g2_decap_8
XFILLER_45_763 VPWR VGND sg13g2_decap_8
XFILLER_33_903 VPWR VGND sg13g2_decap_8
XFILLER_44_273 VPWR VGND sg13g2_decap_8
XFILLER_17_465 VPWR VGND sg13g2_decap_8
XFILLER_32_413 VPWR VGND sg13g2_decap_8
XFILLER_41_980 VPWR VGND sg13g2_decap_8
XFILLER_13_671 VPWR VGND sg13g2_decap_8
XFILLER_12_170 VPWR VGND sg13g2_decap_8
XFILLER_40_490 VPWR VGND sg13g2_decap_8
XFILLER_8_163 VPWR VGND sg13g2_decap_8
XFILLER_9_664 VPWR VGND sg13g2_decap_8
XFILLER_5_892 VPWR VGND sg13g2_decap_8
XFILLER_36_763 VPWR VGND sg13g2_decap_8
XFILLER_24_914 VPWR VGND sg13g2_decap_8
XFILLER_35_273 VPWR VGND sg13g2_decap_8
XFILLER_23_424 VPWR VGND sg13g2_decap_8
XFILLER_10_107 VPWR VGND sg13g2_decap_8
XFILLER_32_980 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_decap_8
XFILLER_31_490 VPWR VGND sg13g2_decap_8
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
XFILLER_27_730 VPWR VGND sg13g2_decap_8
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_42_700 VPWR VGND sg13g2_decap_8
XFILLER_15_925 VPWR VGND sg13g2_decap_8
XFILLER_26_284 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_decap_8
XFILLER_42_777 VPWR VGND sg13g2_decap_8
XFILLER_14_457 VPWR VGND sg13g2_decap_8
XFILLER_30_917 VPWR VGND sg13g2_decap_8
XFILLER_23_991 VPWR VGND sg13g2_decap_8
XFILLER_41_287 VPWR VGND sg13g2_decap_8
XFILLER_5_122 VPWR VGND sg13g2_decap_8
XFILLER_10_674 VPWR VGND sg13g2_decap_8
XFILLER_6_656 VPWR VGND sg13g2_decap_8
XFILLER_5_199 VPWR VGND sg13g2_decap_8
XFILLER_2_840 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_18_752 VPWR VGND sg13g2_decap_8
XFILLER_45_560 VPWR VGND sg13g2_decap_8
XFILLER_17_262 VPWR VGND sg13g2_decap_8
XFILLER_33_700 VPWR VGND sg13g2_decap_8
XFILLER_32_210 VPWR VGND sg13g2_decap_8
XFILLER_21_906 VPWR VGND sg13g2_decap_8
XFILLER_33_777 VPWR VGND sg13g2_decap_8
XFILLER_20_427 VPWR VGND sg13g2_decap_8
XFILLER_32_287 VPWR VGND sg13g2_decap_8
XFILLER_9_461 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_8
XFILLER_24_711 VPWR VGND sg13g2_decap_8
XFILLER_36_560 VPWR VGND sg13g2_decap_8
XFILLER_23_221 VPWR VGND sg13g2_decap_8
XFILLER_24_788 VPWR VGND sg13g2_decap_8
XFILLER_11_427 VPWR VGND sg13g2_decap_8
XFILLER_23_46 VPWR VGND sg13g2_decap_8
XFILLER_23_298 VPWR VGND sg13g2_decap_8
XFILLER_20_994 VPWR VGND sg13g2_decap_8
XFILLER_3_648 VPWR VGND sg13g2_decap_8
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_24_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_19_538 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_15_722 VPWR VGND sg13g2_decap_8
XFILLER_42_574 VPWR VGND sg13g2_decap_8
XFILLER_14_254 VPWR VGND sg13g2_decap_8
XFILLER_30_714 VPWR VGND sg13g2_decap_8
XFILLER_15_799 VPWR VGND sg13g2_decap_8
XFILLER_10_471 VPWR VGND sg13g2_decap_8
XFILLER_7_943 VPWR VGND sg13g2_decap_8
XFILLER_11_994 VPWR VGND sg13g2_decap_8
XFILLER_6_453 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_4 VPWR VGND sg13g2_decap_8
XFILLER_49_151 VPWR VGND sg13g2_decap_8
XFILLER_38_847 VPWR VGND sg13g2_decap_8
X_45_ VGND VPWR net2 net3 _18_ net34 sg13g2_a21oi_1
XFILLER_37_357 VPWR VGND sg13g2_decap_8
XFILLER_25_508 VPWR VGND sg13g2_decap_8
XFILLER_21_703 VPWR VGND sg13g2_decap_8
XFILLER_20_224 VPWR VGND sg13g2_decap_8
XFILLER_33_574 VPWR VGND sg13g2_decap_8
XFILLER_47_1001 VPWR VGND sg13g2_decap_8
XFILLER_18_46 VPWR VGND sg13g2_decap_8
XFILLER_29_858 VPWR VGND sg13g2_decap_8
XFILLER_28_368 VPWR VGND sg13g2_decap_8
XFILLER_24_585 VPWR VGND sg13g2_decap_8
XFILLER_34_56 VPWR VGND sg13g2_decap_8
XFILLER_11_224 VPWR VGND sg13g2_decap_8
XFILLER_12_758 VPWR VGND sg13g2_decap_8
XFILLER_20_791 VPWR VGND sg13g2_decap_8
XFILLER_4_946 VPWR VGND sg13g2_decap_8
XFILLER_3_445 VPWR VGND sg13g2_decap_8
XFILLER_47_644 VPWR VGND sg13g2_decap_8
XFILLER_19_335 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_43_861 VPWR VGND sg13g2_decap_8
XFILLER_42_371 VPWR VGND sg13g2_decap_8
XFILLER_15_596 VPWR VGND sg13g2_decap_8
XFILLER_30_511 VPWR VGND sg13g2_decap_8
XFILLER_30_588 VPWR VGND sg13g2_decap_8
XFILLER_7_740 VPWR VGND sg13g2_decap_8
XFILLER_11_791 VPWR VGND sg13g2_decap_8
XFILLER_6_250 VPWR VGND sg13g2_decap_8
XFILLER_38_644 VPWR VGND sg13g2_decap_8
XFILLER_25_305 VPWR VGND sg13g2_decap_8
XFILLER_37_154 VPWR VGND sg13g2_decap_8
XFILLER_34_861 VPWR VGND sg13g2_decap_8
XFILLER_40_308 VPWR VGND sg13g2_decap_8
XFILLER_21_500 VPWR VGND sg13g2_decap_8
XFILLER_33_371 VPWR VGND sg13g2_decap_8
XFILLER_21_577 VPWR VGND sg13g2_decap_8
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_1_938 VPWR VGND sg13g2_decap_8
XFILLER_0_448 VPWR VGND sg13g2_decap_8
Xhold45 _07_ VPWR VGND net45 sg13g2_dlygate4sd3_1
Xhold34 net4 VPWR VGND net34 sg13g2_dlygate4sd3_1
XFILLER_29_67 VPWR VGND sg13g2_decap_8
XFILLER_21_1004 VPWR VGND sg13g2_decap_8
XFILLER_29_655 VPWR VGND sg13g2_decap_8
XFILLER_28_165 VPWR VGND sg13g2_decap_8
XFILLER_44_658 VPWR VGND sg13g2_decap_8
XFILLER_16_349 VPWR VGND sg13g2_decap_8
XFILLER_45_77 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_8
XFILLER_31_308 VPWR VGND sg13g2_decap_8
XFILLER_25_872 VPWR VGND sg13g2_decap_8
XFILLER_12_555 VPWR VGND sg13g2_decap_8
XFILLER_24_382 VPWR VGND sg13g2_decap_8
XFILLER_40_875 VPWR VGND sg13g2_decap_8
XFILLER_8_548 VPWR VGND sg13g2_decap_8
XFILLER_4_743 VPWR VGND sg13g2_decap_8
XFILLER_3_242 VPWR VGND sg13g2_decap_8
XFILLER_48_931 VPWR VGND sg13g2_decap_8
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_19_132 VPWR VGND sg13g2_fill_2
XFILLER_23_809 VPWR VGND sg13g2_decap_8
XFILLER_35_658 VPWR VGND sg13g2_decap_8
XFILLER_34_168 VPWR VGND sg13g2_decap_8
XFILLER_37_1022 VPWR VGND sg13g2_decap_8
XFILLER_15_393 VPWR VGND sg13g2_decap_8
XFILLER_31_875 VPWR VGND sg13g2_decap_8
XFILLER_30_385 VPWR VGND sg13g2_decap_8
XFILLER_44_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_931 VPWR VGND sg13g2_decap_8
XFILLER_38_441 VPWR VGND sg13g2_decap_8
XFILLER_25_102 VPWR VGND sg13g2_decap_8
XFILLER_26_669 VPWR VGND sg13g2_decap_8
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_25_179 VPWR VGND sg13g2_decap_8
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_22_842 VPWR VGND sg13g2_decap_8
XFILLER_21_374 VPWR VGND sg13g2_decap_8
XFILLER_31_35 VPWR VGND sg13g2_decap_8
XFILLER_5_507 VPWR VGND sg13g2_decap_8
Xoutput13 net13 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_735 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_49_739 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_29_452 VPWR VGND sg13g2_decap_8
XFILLER_45_945 VPWR VGND sg13g2_decap_8
XFILLER_17_647 VPWR VGND sg13g2_decap_8
XFILLER_44_455 VPWR VGND sg13g2_decap_8
XFILLER_16_146 VPWR VGND sg13g2_decap_8
XFILLER_31_105 VPWR VGND sg13g2_decap_8
XFILLER_13_853 VPWR VGND sg13g2_decap_8
XFILLER_12_352 VPWR VGND sg13g2_decap_8
XFILLER_40_672 VPWR VGND sg13g2_decap_8
XFILLER_8_345 VPWR VGND sg13g2_decap_8
XFILLER_9_846 VPWR VGND sg13g2_decap_8
XFILLER_4_540 VPWR VGND sg13g2_decap_8
XFILLER_39_238 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_36_945 VPWR VGND sg13g2_decap_8
XFILLER_23_606 VPWR VGND sg13g2_decap_8
XFILLER_35_455 VPWR VGND sg13g2_decap_8
XFILLER_22_149 VPWR VGND sg13g2_decap_8
XFILLER_15_190 VPWR VGND sg13g2_decap_8
XFILLER_31_672 VPWR VGND sg13g2_decap_8
XFILLER_30_182 VPWR VGND sg13g2_decap_8
XFILLER_27_912 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_fill_1
XFILLER_27_989 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_decap_8
XFILLER_26_466 VPWR VGND sg13g2_decap_8
XFILLER_42_959 VPWR VGND sg13g2_decap_8
XFILLER_13_127 VPWR VGND sg13g2_decap_8
XFILLER_13_138 VPWR VGND sg13g2_fill_2
XFILLER_41_469 VPWR VGND sg13g2_decap_8
XFILLER_42_56 VPWR VGND sg13g2_decap_8
XFILLER_21_171 VPWR VGND sg13g2_decap_8
XFILLER_5_304 VPWR VGND sg13g2_decap_8
XFILLER_10_856 VPWR VGND sg13g2_decap_8
XFILLER_6_838 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_27_1010 VPWR VGND sg13g2_decap_8
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_18_934 VPWR VGND sg13g2_decap_8
XFILLER_45_742 VPWR VGND sg13g2_decap_8
XFILLER_17_444 VPWR VGND sg13g2_decap_8
XFILLER_44_252 VPWR VGND sg13g2_decap_8
XFILLER_33_959 VPWR VGND sg13g2_decap_8
XFILLER_13_650 VPWR VGND sg13g2_decap_8
XFILLER_20_609 VPWR VGND sg13g2_decap_8
XFILLER_32_469 VPWR VGND sg13g2_decap_8
XFILLER_9_643 VPWR VGND sg13g2_decap_8
XFILLER_8_142 VPWR VGND sg13g2_decap_8
XFILLER_5_871 VPWR VGND sg13g2_decap_8
XFILLER_27_219 VPWR VGND sg13g2_decap_8
XFILLER_36_742 VPWR VGND sg13g2_decap_8
XFILLER_23_403 VPWR VGND sg13g2_decap_8
XFILLER_35_252 VPWR VGND sg13g2_decap_8
XFILLER_11_609 VPWR VGND sg13g2_decap_8
XFILLER_2_329 VPWR VGND sg13g2_decap_8
XFILLER_46_539 VPWR VGND sg13g2_decap_8
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_15_904 VPWR VGND sg13g2_decap_8
XFILLER_26_263 VPWR VGND sg13g2_decap_8
XFILLER_27_786 VPWR VGND sg13g2_decap_8
XFILLER_42_756 VPWR VGND sg13g2_decap_8
XFILLER_14_436 VPWR VGND sg13g2_decap_8
XFILLER_23_970 VPWR VGND sg13g2_decap_8
XFILLER_41_266 VPWR VGND sg13g2_decap_8
XFILLER_10_653 VPWR VGND sg13g2_decap_8
XFILLER_6_635 VPWR VGND sg13g2_decap_8
XFILLER_5_101 VPWR VGND sg13g2_decap_8
XFILLER_5_178 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_2_896 VPWR VGND sg13g2_decap_8
X_61_ net21 VGND VPWR net45 net7 clknet_1_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_37_539 VPWR VGND sg13g2_decap_8
XFILLER_18_731 VPWR VGND sg13g2_decap_8
XFILLER_17_241 VPWR VGND sg13g2_decap_8
XFILLER_33_756 VPWR VGND sg13g2_decap_8
XFILLER_20_406 VPWR VGND sg13g2_decap_8
XFILLER_32_266 VPWR VGND sg13g2_decap_8
XFILLER_9_440 VPWR VGND sg13g2_decap_8
XFILLER_23_200 VPWR VGND sg13g2_decap_8
XFILLER_11_406 VPWR VGND sg13g2_decap_8
XFILLER_24_767 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_8
XFILLER_23_277 VPWR VGND sg13g2_decap_8
XFILLER_20_973 VPWR VGND sg13g2_decap_8
XFILLER_3_627 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_47_826 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_19_517 VPWR VGND sg13g2_decap_8
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_15_701 VPWR VGND sg13g2_decap_8
XFILLER_27_583 VPWR VGND sg13g2_decap_8
XFILLER_42_553 VPWR VGND sg13g2_decap_8
XFILLER_14_233 VPWR VGND sg13g2_decap_8
XFILLER_15_778 VPWR VGND sg13g2_decap_8
XFILLER_10_450 VPWR VGND sg13g2_decap_8
XFILLER_7_922 VPWR VGND sg13g2_decap_8
XFILLER_11_973 VPWR VGND sg13g2_decap_8
XFILLER_6_432 VPWR VGND sg13g2_decap_8
XFILLER_7_999 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_9_1007 VPWR VGND sg13g2_decap_8
XFILLER_2_693 VPWR VGND sg13g2_decap_8
XFILLER_49_130 VPWR VGND sg13g2_decap_8
XFILLER_38_826 VPWR VGND sg13g2_decap_8
X_44_ VGND VPWR net2 net47 _03_ _17_ sg13g2_a21oi_1
XFILLER_37_336 VPWR VGND sg13g2_decap_8
XFILLER_33_553 VPWR VGND sg13g2_decap_8
XFILLER_20_203 VPWR VGND sg13g2_decap_8
XFILLER_21_759 VPWR VGND sg13g2_decap_8
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_29_837 VPWR VGND sg13g2_decap_8
XFILLER_28_347 VPWR VGND sg13g2_decap_8
XFILLER_24_564 VPWR VGND sg13g2_decap_8
XFILLER_34_35 VPWR VGND sg13g2_decap_8
XFILLER_11_203 VPWR VGND sg13g2_decap_8
XFILLER_12_737 VPWR VGND sg13g2_decap_8
XFILLER_7_229 VPWR VGND sg13g2_decap_8
XFILLER_20_770 VPWR VGND sg13g2_decap_8
XFILLER_4_925 VPWR VGND sg13g2_decap_8
XFILLER_3_424 VPWR VGND sg13g2_decap_8
XFILLER_47_623 VPWR VGND sg13g2_decap_8
XFILLER_19_314 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_27_380 VPWR VGND sg13g2_decap_8
XFILLER_43_840 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_decap_8
XFILLER_15_575 VPWR VGND sg13g2_decap_8
XFILLER_11_770 VPWR VGND sg13g2_decap_8
XFILLER_30_567 VPWR VGND sg13g2_decap_8
XFILLER_7_796 VPWR VGND sg13g2_decap_8
XFILLER_3_991 VPWR VGND sg13g2_decap_8
XFILLER_2_490 VPWR VGND sg13g2_decap_8
XFILLER_38_623 VPWR VGND sg13g2_decap_8
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_19_881 VPWR VGND sg13g2_decap_8
XFILLER_34_840 VPWR VGND sg13g2_decap_8
XFILLER_33_350 VPWR VGND sg13g2_decap_8
XFILLER_21_556 VPWR VGND sg13g2_decap_8
XFILLER_1_917 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
Xhold35 _18_ VPWR VGND net35 sg13g2_dlygate4sd3_1
Xhold46 net8 VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_29_46 VPWR VGND sg13g2_decap_8
XFILLER_29_634 VPWR VGND sg13g2_decap_8
XFILLER_17_829 VPWR VGND sg13g2_decap_8
XFILLER_28_144 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
XFILLER_44_637 VPWR VGND sg13g2_decap_8
XFILLER_16_328 VPWR VGND sg13g2_decap_8
XFILLER_43_147 VPWR VGND sg13g2_decap_8
XFILLER_25_851 VPWR VGND sg13g2_decap_8
XFILLER_24_361 VPWR VGND sg13g2_decap_8
XFILLER_12_534 VPWR VGND sg13g2_decap_8
XFILLER_40_854 VPWR VGND sg13g2_decap_8
XFILLER_8_527 VPWR VGND sg13g2_decap_8
XFILLER_4_722 VPWR VGND sg13g2_decap_8
XFILLER_3_221 VPWR VGND sg13g2_decap_8
XFILLER_4_799 VPWR VGND sg13g2_decap_8
XFILLER_3_298 VPWR VGND sg13g2_decap_8
XFILLER_48_910 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_19_111 VPWR VGND sg13g2_decap_8
XFILLER_48_987 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_19_188 VPWR VGND sg13g2_decap_8
XFILLER_35_637 VPWR VGND sg13g2_decap_8
XFILLER_34_147 VPWR VGND sg13g2_decap_8
XFILLER_37_1001 VPWR VGND sg13g2_decap_8
XFILLER_15_372 VPWR VGND sg13g2_decap_8
XFILLER_16_895 VPWR VGND sg13g2_decap_8
XFILLER_31_854 VPWR VGND sg13g2_decap_8
XFILLER_30_364 VPWR VGND sg13g2_decap_8
XFILLER_7_593 VPWR VGND sg13g2_decap_8
XFILLER_32_0 VPWR VGND sg13g2_decap_8
XFILLER_39_910 VPWR VGND sg13g2_decap_8
XFILLER_38_420 VPWR VGND sg13g2_decap_8
XFILLER_39_987 VPWR VGND sg13g2_decap_8
XFILLER_26_648 VPWR VGND sg13g2_decap_8
XFILLER_38_497 VPWR VGND sg13g2_decap_8
XFILLER_25_158 VPWR VGND sg13g2_decap_8
XFILLER_22_821 VPWR VGND sg13g2_decap_8
XFILLER_21_353 VPWR VGND sg13g2_decap_8
XFILLER_22_898 VPWR VGND sg13g2_decap_8
XFILLER_31_14 VPWR VGND sg13g2_decap_8
Xoutput14 net14 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_714 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_49_718 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_29_431 VPWR VGND sg13g2_decap_8
XFILLER_45_924 VPWR VGND sg13g2_decap_8
XFILLER_17_626 VPWR VGND sg13g2_decap_8
XFILLER_44_434 VPWR VGND sg13g2_decap_8
XFILLER_16_125 VPWR VGND sg13g2_decap_8
XFILLER_13_832 VPWR VGND sg13g2_decap_8
XFILLER_9_825 VPWR VGND sg13g2_decap_8
XFILLER_12_331 VPWR VGND sg13g2_decap_8
XFILLER_40_651 VPWR VGND sg13g2_decap_8
XFILLER_8_324 VPWR VGND sg13g2_decap_8
XFILLER_21_91 VPWR VGND sg13g2_fill_1
XFILLER_4_596 VPWR VGND sg13g2_decap_8
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_39_217 VPWR VGND sg13g2_decap_8
XFILLER_48_784 VPWR VGND sg13g2_decap_8
XFILLER_36_924 VPWR VGND sg13g2_decap_8
XFILLER_47_294 VPWR VGND sg13g2_decap_8
XFILLER_35_434 VPWR VGND sg13g2_decap_8
XFILLER_16_692 VPWR VGND sg13g2_decap_8
XFILLER_22_128 VPWR VGND sg13g2_decap_8
XFILLER_31_651 VPWR VGND sg13g2_decap_8
XFILLER_30_161 VPWR VGND sg13g2_decap_8
XFILLER_8_891 VPWR VGND sg13g2_decap_8
XFILLER_7_82 VPWR VGND sg13g2_decap_8
XFILLER_11_1015 VPWR VGND sg13g2_decap_8
XFILLER_7_390 VPWR VGND sg13g2_decap_8
XFILLER_39_784 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_fill_2
XFILLER_26_445 VPWR VGND sg13g2_decap_8
XFILLER_27_968 VPWR VGND sg13g2_decap_8
XFILLER_38_294 VPWR VGND sg13g2_decap_8
XFILLER_42_938 VPWR VGND sg13g2_decap_8
XFILLER_13_106 VPWR VGND sg13g2_decap_8
XFILLER_14_618 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_decap_8
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_10_835 VPWR VGND sg13g2_decap_8
XFILLER_21_150 VPWR VGND sg13g2_decap_8
XFILLER_22_695 VPWR VGND sg13g2_decap_8
XFILLER_6_817 VPWR VGND sg13g2_decap_8
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
XFILLER_45_721 VPWR VGND sg13g2_decap_8
XFILLER_18_913 VPWR VGND sg13g2_decap_8
XFILLER_44_231 VPWR VGND sg13g2_decap_8
XFILLER_17_423 VPWR VGND sg13g2_decap_8
XFILLER_45_798 VPWR VGND sg13g2_decap_8
XFILLER_33_938 VPWR VGND sg13g2_decap_8
XFILLER_32_448 VPWR VGND sg13g2_decap_8
XFILLER_34_1015 VPWR VGND sg13g2_decap_8
XFILLER_9_622 VPWR VGND sg13g2_decap_8
XFILLER_9_699 VPWR VGND sg13g2_decap_8
XFILLER_8_198 VPWR VGND sg13g2_decap_8
XFILLER_5_850 VPWR VGND sg13g2_decap_8
XFILLER_4_393 VPWR VGND sg13g2_decap_8
XFILLER_41_1008 VPWR VGND sg13g2_decap_8
XFILLER_48_581 VPWR VGND sg13g2_decap_8
XFILLER_36_721 VPWR VGND sg13g2_decap_8
XFILLER_35_231 VPWR VGND sg13g2_decap_8
XFILLER_36_798 VPWR VGND sg13g2_decap_8
XFILLER_17_990 VPWR VGND sg13g2_decap_8
XFILLER_24_949 VPWR VGND sg13g2_decap_8
XFILLER_23_459 VPWR VGND sg13g2_decap_8
XFILLER_3_809 VPWR VGND sg13g2_decap_8
XFILLER_2_308 VPWR VGND sg13g2_decap_8
XFILLER_46_518 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_39_581 VPWR VGND sg13g2_decap_8
XFILLER_26_242 VPWR VGND sg13g2_decap_8
XFILLER_27_765 VPWR VGND sg13g2_decap_8
XFILLER_42_735 VPWR VGND sg13g2_decap_8
XFILLER_14_415 VPWR VGND sg13g2_decap_8
XFILLER_41_245 VPWR VGND sg13g2_decap_8
XFILLER_10_632 VPWR VGND sg13g2_decap_8
XFILLER_22_492 VPWR VGND sg13g2_decap_8
XFILLER_6_614 VPWR VGND sg13g2_decap_8
XFILLER_5_157 VPWR VGND sg13g2_decap_8
XFILLER_2_875 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
X_60_ net19 VGND VPWR net43 net6 clknet_1_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_18_710 VPWR VGND sg13g2_decap_8
XFILLER_37_518 VPWR VGND sg13g2_decap_8
XFILLER_17_220 VPWR VGND sg13g2_decap_8
XFILLER_18_787 VPWR VGND sg13g2_decap_8
XFILLER_45_595 VPWR VGND sg13g2_decap_8
XFILLER_17_297 VPWR VGND sg13g2_decap_8
XFILLER_33_735 VPWR VGND sg13g2_decap_8
XFILLER_32_245 VPWR VGND sg13g2_decap_8
XFILLER_14_982 VPWR VGND sg13g2_decap_8
XFILLER_9_496 VPWR VGND sg13g2_decap_8
XFILLER_4_190 VPWR VGND sg13g2_decap_8
XFILLER_28_529 VPWR VGND sg13g2_decap_8
XFILLER_24_746 VPWR VGND sg13g2_decap_8
XFILLER_36_595 VPWR VGND sg13g2_decap_8
XFILLER_12_919 VPWR VGND sg13g2_decap_8
XFILLER_23_256 VPWR VGND sg13g2_decap_8
XFILLER_20_952 VPWR VGND sg13g2_decap_8
XFILLER_3_606 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_27_562 VPWR VGND sg13g2_decap_8
XFILLER_14_212 VPWR VGND sg13g2_decap_8
XFILLER_42_532 VPWR VGND sg13g2_decap_8
XFILLER_15_757 VPWR VGND sg13g2_decap_8
XFILLER_9_39 VPWR VGND sg13g2_decap_8
XFILLER_14_289 VPWR VGND sg13g2_decap_8
XFILLER_7_901 VPWR VGND sg13g2_decap_8
XFILLER_11_952 VPWR VGND sg13g2_decap_8
XFILLER_30_749 VPWR VGND sg13g2_decap_8
XFILLER_6_411 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_7_978 VPWR VGND sg13g2_decap_8
XFILLER_6_488 VPWR VGND sg13g2_decap_8
XFILLER_2_672 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_38_805 VPWR VGND sg13g2_decap_8
X_43_ net1 VPWR _17_ VGND net2 net47 sg13g2_o21ai_1
XFILLER_37_315 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_decap_8
XFILLER_46_882 VPWR VGND sg13g2_decap_8
XFILLER_18_584 VPWR VGND sg13g2_decap_8
XFILLER_45_392 VPWR VGND sg13g2_decap_8
XFILLER_33_532 VPWR VGND sg13g2_decap_8
XFILLER_21_738 VPWR VGND sg13g2_decap_8
XFILLER_20_259 VPWR VGND sg13g2_decap_8
XFILLER_9_293 VPWR VGND sg13g2_decap_8
XFILLER_0_609 VPWR VGND sg13g2_decap_8
XFILLER_29_816 VPWR VGND sg13g2_decap_8
XFILLER_28_326 VPWR VGND sg13g2_decap_8
XFILLER_44_819 VPWR VGND sg13g2_decap_8
XFILLER_43_329 VPWR VGND sg13g2_decap_8
XFILLER_37_882 VPWR VGND sg13g2_decap_8
XFILLER_24_543 VPWR VGND sg13g2_decap_8
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_36_392 VPWR VGND sg13g2_decap_8
XFILLER_12_716 VPWR VGND sg13g2_decap_8
XFILLER_8_709 VPWR VGND sg13g2_decap_8
XFILLER_7_208 VPWR VGND sg13g2_decap_8
XFILLER_11_259 VPWR VGND sg13g2_decap_8
XFILLER_4_904 VPWR VGND sg13g2_decap_8
XFILLER_3_403 VPWR VGND sg13g2_decap_8
XFILLER_47_602 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_47_679 VPWR VGND sg13g2_decap_8
XFILLER_35_819 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_28_893 VPWR VGND sg13g2_decap_8
XFILLER_34_329 VPWR VGND sg13g2_decap_8
XFILLER_15_554 VPWR VGND sg13g2_decap_8
XFILLER_43_896 VPWR VGND sg13g2_decap_8
XFILLER_30_546 VPWR VGND sg13g2_decap_8
XFILLER_7_775 VPWR VGND sg13g2_decap_8
XFILLER_6_285 VPWR VGND sg13g2_decap_8
XFILLER_3_970 VPWR VGND sg13g2_decap_8
XFILLER_38_602 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_19_860 VPWR VGND sg13g2_decap_8
XFILLER_38_679 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_37_189 VPWR VGND sg13g2_decap_8
XFILLER_18_381 VPWR VGND sg13g2_decap_8
XFILLER_34_896 VPWR VGND sg13g2_decap_8
XFILLER_21_535 VPWR VGND sg13g2_decap_8
XFILLER_14_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_29_25 VPWR VGND sg13g2_decap_8
Xhold36 net10 VPWR VGND net36 sg13g2_dlygate4sd3_1
Xhold47 net3 VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_29_613 VPWR VGND sg13g2_decap_8
XFILLER_28_123 VPWR VGND sg13g2_decap_8
XFILLER_17_808 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_44_616 VPWR VGND sg13g2_decap_8
XFILLER_16_307 VPWR VGND sg13g2_decap_8
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_25_830 VPWR VGND sg13g2_decap_8
XFILLER_24_340 VPWR VGND sg13g2_decap_8
XFILLER_12_513 VPWR VGND sg13g2_decap_8
XFILLER_40_833 VPWR VGND sg13g2_decap_8
XFILLER_8_506 VPWR VGND sg13g2_decap_8
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_4_701 VPWR VGND sg13g2_decap_8
XFILLER_3_200 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_4
XFILLER_4_778 VPWR VGND sg13g2_decap_8
XFILLER_3_277 VPWR VGND sg13g2_decap_8
XFILLER_10_93 VPWR VGND sg13g2_decap_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
XFILLER_48_966 VPWR VGND sg13g2_decap_8
XFILLER_19_134 VPWR VGND sg13g2_fill_1
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_19_167 VPWR VGND sg13g2_decap_8
XFILLER_35_616 VPWR VGND sg13g2_decap_8
XFILLER_28_690 VPWR VGND sg13g2_decap_8
XFILLER_34_126 VPWR VGND sg13g2_decap_8
XFILLER_15_351 VPWR VGND sg13g2_decap_8
XFILLER_16_874 VPWR VGND sg13g2_decap_8
XFILLER_43_693 VPWR VGND sg13g2_decap_8
XFILLER_31_833 VPWR VGND sg13g2_decap_8
XFILLER_30_343 VPWR VGND sg13g2_decap_8
XFILLER_7_572 VPWR VGND sg13g2_decap_8
Xheichips25_template_27 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_39_966 VPWR VGND sg13g2_decap_8
XFILLER_26_627 VPWR VGND sg13g2_decap_8
XFILLER_38_476 VPWR VGND sg13g2_decap_8
XFILLER_25_137 VPWR VGND sg13g2_decap_8
XFILLER_22_800 VPWR VGND sg13g2_decap_8
XFILLER_34_693 VPWR VGND sg13g2_decap_8
XFILLER_21_332 VPWR VGND sg13g2_decap_8
XFILLER_22_877 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_5_1011 VPWR VGND sg13g2_decap_8
XFILLER_29_410 VPWR VGND sg13g2_decap_8
XFILLER_45_903 VPWR VGND sg13g2_decap_8
XFILLER_44_413 VPWR VGND sg13g2_decap_8
XFILLER_16_104 VPWR VGND sg13g2_decap_8
XFILLER_17_605 VPWR VGND sg13g2_decap_8
XFILLER_29_487 VPWR VGND sg13g2_decap_8
XFILLER_13_811 VPWR VGND sg13g2_decap_8
XFILLER_12_310 VPWR VGND sg13g2_decap_8
XFILLER_40_630 VPWR VGND sg13g2_decap_8
XFILLER_8_303 VPWR VGND sg13g2_decap_8
XFILLER_9_804 VPWR VGND sg13g2_decap_8
XFILLER_12_387 VPWR VGND sg13g2_decap_8
XFILLER_13_888 VPWR VGND sg13g2_decap_8
XFILLER_4_575 VPWR VGND sg13g2_decap_8
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_48_763 VPWR VGND sg13g2_decap_8
XFILLER_36_903 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_35_413 VPWR VGND sg13g2_decap_8
XFILLER_22_107 VPWR VGND sg13g2_decap_8
XFILLER_44_980 VPWR VGND sg13g2_decap_8
XFILLER_16_671 VPWR VGND sg13g2_decap_8
XFILLER_43_490 VPWR VGND sg13g2_decap_8
XFILLER_31_630 VPWR VGND sg13g2_decap_8
XFILLER_30_140 VPWR VGND sg13g2_decap_8
XFILLER_8_870 VPWR VGND sg13g2_decap_8
XFILLER_7_61 VPWR VGND sg13g2_decap_8
XFILLER_39_763 VPWR VGND sg13g2_decap_8
XFILLER_38_273 VPWR VGND sg13g2_decap_8
XFILLER_26_424 VPWR VGND sg13g2_decap_8
XFILLER_27_947 VPWR VGND sg13g2_decap_8
XFILLER_42_917 VPWR VGND sg13g2_decap_8
XFILLER_41_427 VPWR VGND sg13g2_decap_8
XFILLER_35_980 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_34_490 VPWR VGND sg13g2_decap_8
XFILLER_10_814 VPWR VGND sg13g2_decap_8
XFILLER_22_674 VPWR VGND sg13g2_decap_8
XFILLER_5_339 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_45_700 VPWR VGND sg13g2_decap_8
XFILLER_17_402 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_decap_8
XFILLER_18_969 VPWR VGND sg13g2_decap_8
XFILLER_29_284 VPWR VGND sg13g2_decap_8
XFILLER_45_777 VPWR VGND sg13g2_decap_8
XFILLER_17_479 VPWR VGND sg13g2_decap_8
XFILLER_33_917 VPWR VGND sg13g2_decap_8
XFILLER_44_287 VPWR VGND sg13g2_decap_8
XFILLER_26_991 VPWR VGND sg13g2_decap_8
XFILLER_32_427 VPWR VGND sg13g2_decap_8
XFILLER_9_601 VPWR VGND sg13g2_decap_8
XFILLER_41_994 VPWR VGND sg13g2_decap_8
XFILLER_13_685 VPWR VGND sg13g2_decap_8
XFILLER_9_678 VPWR VGND sg13g2_decap_8
XFILLER_12_184 VPWR VGND sg13g2_decap_8
XFILLER_8_177 VPWR VGND sg13g2_decap_8
XFILLER_32_91 VPWR VGND sg13g2_decap_8
XFILLER_4_372 VPWR VGND sg13g2_decap_8
XFILLER_48_560 VPWR VGND sg13g2_decap_8
XFILLER_36_700 VPWR VGND sg13g2_decap_8
XFILLER_35_210 VPWR VGND sg13g2_decap_8
XFILLER_24_928 VPWR VGND sg13g2_decap_8
XFILLER_36_777 VPWR VGND sg13g2_decap_8
XFILLER_23_438 VPWR VGND sg13g2_decap_8
XFILLER_35_287 VPWR VGND sg13g2_decap_8
XFILLER_32_994 VPWR VGND sg13g2_decap_8
XFILLER_12_39 VPWR VGND sg13g2_decap_8
XFILLER_37_14 VPWR VGND sg13g2_decap_8
XFILLER_39_560 VPWR VGND sg13g2_decap_8
XFILLER_26_221 VPWR VGND sg13g2_decap_8
XFILLER_27_744 VPWR VGND sg13g2_decap_8
XFILLER_42_714 VPWR VGND sg13g2_decap_8
XFILLER_15_939 VPWR VGND sg13g2_decap_8
XFILLER_26_298 VPWR VGND sg13g2_decap_8
XFILLER_41_224 VPWR VGND sg13g2_decap_8
XFILLER_10_611 VPWR VGND sg13g2_decap_8
XFILLER_22_471 VPWR VGND sg13g2_decap_8
XFILLER_5_136 VPWR VGND sg13g2_decap_8
XFILLER_10_688 VPWR VGND sg13g2_decap_8
XFILLER_2_854 VPWR VGND sg13g2_decap_8
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_18_766 VPWR VGND sg13g2_decap_8
XFILLER_45_574 VPWR VGND sg13g2_decap_8
XFILLER_17_276 VPWR VGND sg13g2_decap_8
XFILLER_33_714 VPWR VGND sg13g2_decap_8
XFILLER_32_224 VPWR VGND sg13g2_decap_8
XFILLER_14_961 VPWR VGND sg13g2_decap_8
XFILLER_41_791 VPWR VGND sg13g2_decap_8
XFILLER_13_482 VPWR VGND sg13g2_decap_8
XFILLER_9_475 VPWR VGND sg13g2_decap_8
XFILLER_4_95 VPWR VGND sg13g2_decap_8
XFILLER_4_84 VPWR VGND sg13g2_decap_4
XFILLER_28_508 VPWR VGND sg13g2_decap_8
XFILLER_24_725 VPWR VGND sg13g2_decap_8
XFILLER_36_574 VPWR VGND sg13g2_decap_8
XFILLER_23_235 VPWR VGND sg13g2_decap_8
XFILLER_17_1011 VPWR VGND sg13g2_decap_8
XFILLER_20_931 VPWR VGND sg13g2_decap_8
XFILLER_32_791 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_24_1026 VPWR VGND sg13g2_fill_2
XFILLER_27_541 VPWR VGND sg13g2_decap_8
XFILLER_42_511 VPWR VGND sg13g2_decap_8
XFILLER_15_736 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_fill_2
XFILLER_42_588 VPWR VGND sg13g2_decap_8
XFILLER_14_268 VPWR VGND sg13g2_decap_8
XFILLER_30_728 VPWR VGND sg13g2_decap_8
XFILLER_11_931 VPWR VGND sg13g2_decap_8
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_31_1008 VPWR VGND sg13g2_decap_8
XFILLER_10_485 VPWR VGND sg13g2_decap_8
XFILLER_7_957 VPWR VGND sg13g2_decap_8
XFILLER_6_467 VPWR VGND sg13g2_decap_8
XFILLER_2_651 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_49_165 VPWR VGND sg13g2_decap_8
X_42_ VGND VPWR net36 _15_ _02_ _16_ sg13g2_a21oi_1
XFILLER_46_861 VPWR VGND sg13g2_decap_8
XFILLER_45_371 VPWR VGND sg13g2_decap_8
XFILLER_18_563 VPWR VGND sg13g2_decap_8
XFILLER_33_511 VPWR VGND sg13g2_decap_8
XFILLER_21_717 VPWR VGND sg13g2_decap_8
XFILLER_33_588 VPWR VGND sg13g2_decap_8
XFILLER_20_238 VPWR VGND sg13g2_decap_8
XFILLER_9_272 VPWR VGND sg13g2_decap_8
XFILLER_47_1015 VPWR VGND sg13g2_decap_8
XFILLER_28_305 VPWR VGND sg13g2_decap_8
XFILLER_43_308 VPWR VGND sg13g2_decap_8
XFILLER_37_861 VPWR VGND sg13g2_decap_8
XFILLER_36_371 VPWR VGND sg13g2_decap_8
XFILLER_24_522 VPWR VGND sg13g2_decap_8
XFILLER_11_238 VPWR VGND sg13g2_decap_8
XFILLER_24_599 VPWR VGND sg13g2_decap_8
XFILLER_3_459 VPWR VGND sg13g2_decap_8
XFILLER_47_658 VPWR VGND sg13g2_decap_8
XFILLER_19_349 VPWR VGND sg13g2_decap_8
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_28_872 VPWR VGND sg13g2_decap_8
XFILLER_34_308 VPWR VGND sg13g2_decap_8
XFILLER_15_533 VPWR VGND sg13g2_decap_8
XFILLER_43_875 VPWR VGND sg13g2_decap_8
XFILLER_42_385 VPWR VGND sg13g2_decap_8
XFILLER_30_525 VPWR VGND sg13g2_decap_8
XFILLER_24_81 VPWR VGND sg13g2_decap_8
XFILLER_10_282 VPWR VGND sg13g2_decap_8
XFILLER_7_754 VPWR VGND sg13g2_decap_8
XFILLER_6_264 VPWR VGND sg13g2_decap_8
XFILLER_40_91 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_26_809 VPWR VGND sg13g2_decap_8
XFILLER_38_658 VPWR VGND sg13g2_decap_8
XFILLER_18_360 VPWR VGND sg13g2_decap_8
XFILLER_25_319 VPWR VGND sg13g2_decap_8
XFILLER_37_168 VPWR VGND sg13g2_decap_8
XFILLER_34_875 VPWR VGND sg13g2_decap_8
XFILLER_21_514 VPWR VGND sg13g2_decap_8
XFILLER_33_385 VPWR VGND sg13g2_decap_8
XFILLER_14_1003 VPWR VGND sg13g2_decap_8
XFILLER_20_39 VPWR VGND sg13g2_decap_8
Xhold37 _02_ VPWR VGND net37 sg13g2_dlygate4sd3_1
Xhold48 net5 VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_21_1018 VPWR VGND sg13g2_decap_8
XFILLER_28_102 VPWR VGND sg13g2_decap_8
XFILLER_29_669 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_28_179 VPWR VGND sg13g2_decap_8
XFILLER_25_886 VPWR VGND sg13g2_decap_8
XFILLER_40_812 VPWR VGND sg13g2_decap_8
XFILLER_24_396 VPWR VGND sg13g2_decap_8
XFILLER_12_569 VPWR VGND sg13g2_decap_8
XFILLER_40_889 VPWR VGND sg13g2_decap_8
XFILLER_4_757 VPWR VGND sg13g2_decap_8
XFILLER_10_72 VPWR VGND sg13g2_decap_8
XFILLER_3_256 VPWR VGND sg13g2_decap_8
XFILLER_0_952 VPWR VGND sg13g2_decap_8
XFILLER_48_945 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_4
XFILLER_19_146 VPWR VGND sg13g2_decap_8
XFILLER_34_105 VPWR VGND sg13g2_decap_8
XFILLER_16_853 VPWR VGND sg13g2_decap_8
XFILLER_43_672 VPWR VGND sg13g2_decap_8
XFILLER_15_330 VPWR VGND sg13g2_decap_8
XFILLER_31_812 VPWR VGND sg13g2_decap_8
XFILLER_42_182 VPWR VGND sg13g2_decap_8
XFILLER_30_322 VPWR VGND sg13g2_decap_8
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_31_889 VPWR VGND sg13g2_decap_8
XFILLER_7_551 VPWR VGND sg13g2_decap_8
XFILLER_30_399 VPWR VGND sg13g2_decap_8
Xheichips25_template_28 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_39_945 VPWR VGND sg13g2_decap_8
XFILLER_38_455 VPWR VGND sg13g2_decap_8
XFILLER_26_606 VPWR VGND sg13g2_decap_8
XFILLER_25_116 VPWR VGND sg13g2_decap_8
XFILLER_41_609 VPWR VGND sg13g2_decap_8
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_21_311 VPWR VGND sg13g2_decap_8
XFILLER_34_672 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
XFILLER_22_856 VPWR VGND sg13g2_decap_8
XFILLER_33_182 VPWR VGND sg13g2_decap_8
XFILLER_21_388 VPWR VGND sg13g2_decap_8
XFILLER_31_49 VPWR VGND sg13g2_decap_8
Xoutput16 net16 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_749 VPWR VGND sg13g2_decap_8
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_29_466 VPWR VGND sg13g2_decap_8
XFILLER_45_959 VPWR VGND sg13g2_decap_8
XFILLER_44_469 VPWR VGND sg13g2_decap_8
XFILLER_32_609 VPWR VGND sg13g2_decap_8
XFILLER_25_683 VPWR VGND sg13g2_decap_8
XFILLER_31_119 VPWR VGND sg13g2_decap_8
XFILLER_13_867 VPWR VGND sg13g2_decap_8
XFILLER_24_193 VPWR VGND sg13g2_decap_8
XFILLER_12_366 VPWR VGND sg13g2_decap_8
XFILLER_40_686 VPWR VGND sg13g2_decap_8
XFILLER_8_359 VPWR VGND sg13g2_decap_8
XFILLER_21_60 VPWR VGND sg13g2_decap_8
XFILLER_4_554 VPWR VGND sg13g2_decap_8
XFILLER_48_742 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_36_959 VPWR VGND sg13g2_decap_8
XFILLER_16_650 VPWR VGND sg13g2_decap_8
XFILLER_35_469 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clknet_0_clk clk VPWR VGND sg13g2_buf_16
XFILLER_31_686 VPWR VGND sg13g2_decap_8
XFILLER_30_196 VPWR VGND sg13g2_decap_8
XFILLER_39_742 VPWR VGND sg13g2_decap_8
XFILLER_26_403 VPWR VGND sg13g2_decap_8
XFILLER_27_926 VPWR VGND sg13g2_decap_8
XFILLER_38_252 VPWR VGND sg13g2_decap_8
XFILLER_41_406 VPWR VGND sg13g2_decap_8
XFILLER_22_653 VPWR VGND sg13g2_decap_8
XFILLER_21_185 VPWR VGND sg13g2_decap_8
XFILLER_5_318 VPWR VGND sg13g2_decap_8
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_27_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_263 VPWR VGND sg13g2_decap_8
XFILLER_18_948 VPWR VGND sg13g2_decap_8
XFILLER_45_756 VPWR VGND sg13g2_decap_8
XFILLER_17_458 VPWR VGND sg13g2_decap_8
XFILLER_32_406 VPWR VGND sg13g2_decap_8
XFILLER_44_266 VPWR VGND sg13g2_decap_8
XFILLER_26_970 VPWR VGND sg13g2_decap_8
XFILLER_16_93 VPWR VGND sg13g2_decap_4
XFILLER_25_480 VPWR VGND sg13g2_decap_8
XFILLER_41_973 VPWR VGND sg13g2_decap_8
XFILLER_12_130 VPWR VGND sg13g2_decap_8
XFILLER_12_163 VPWR VGND sg13g2_decap_8
XFILLER_13_664 VPWR VGND sg13g2_decap_8
XFILLER_9_657 VPWR VGND sg13g2_decap_8
XFILLER_40_483 VPWR VGND sg13g2_decap_8
XFILLER_8_156 VPWR VGND sg13g2_decap_8
XFILLER_32_70 VPWR VGND sg13g2_decap_8
XFILLER_4_351 VPWR VGND sg13g2_decap_8
XFILLER_5_885 VPWR VGND sg13g2_decap_8
XFILLER_24_907 VPWR VGND sg13g2_decap_8
XFILLER_36_756 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_decap_8
XFILLER_35_266 VPWR VGND sg13g2_decap_8
XFILLER_32_973 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
XFILLER_31_483 VPWR VGND sg13g2_decap_8
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_26_200 VPWR VGND sg13g2_decap_8
XFILLER_27_723 VPWR VGND sg13g2_decap_8
XFILLER_15_918 VPWR VGND sg13g2_decap_8
XFILLER_26_277 VPWR VGND sg13g2_decap_8
XFILLER_41_203 VPWR VGND sg13g2_decap_8
XFILLER_22_450 VPWR VGND sg13g2_decap_8
XFILLER_23_984 VPWR VGND sg13g2_decap_8
XFILLER_10_667 VPWR VGND sg13g2_decap_8
XFILLER_6_649 VPWR VGND sg13g2_decap_8
XFILLER_5_115 VPWR VGND sg13g2_decap_8
XFILLER_2_833 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_18_745 VPWR VGND sg13g2_decap_8
XFILLER_45_553 VPWR VGND sg13g2_decap_8
XFILLER_17_255 VPWR VGND sg13g2_decap_8
XFILLER_32_203 VPWR VGND sg13g2_decap_8
XFILLER_14_940 VPWR VGND sg13g2_decap_8
XFILLER_41_770 VPWR VGND sg13g2_decap_8
XFILLER_13_461 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
XFILLER_40_280 VPWR VGND sg13g2_decap_8
XFILLER_9_454 VPWR VGND sg13g2_decap_8
XFILLER_5_682 VPWR VGND sg13g2_decap_8
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_24_704 VPWR VGND sg13g2_decap_8
XFILLER_36_553 VPWR VGND sg13g2_decap_8
XFILLER_23_214 VPWR VGND sg13g2_decap_8
XFILLER_20_910 VPWR VGND sg13g2_decap_8
XFILLER_32_770 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_decap_8
XFILLER_31_280 VPWR VGND sg13g2_decap_8
XFILLER_20_987 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1005 VPWR VGND sg13g2_decap_8
XFILLER_27_520 VPWR VGND sg13g2_decap_8
XFILLER_15_715 VPWR VGND sg13g2_decap_8
XFILLER_14_247 VPWR VGND sg13g2_decap_8
XFILLER_27_597 VPWR VGND sg13g2_decap_8
XFILLER_42_567 VPWR VGND sg13g2_decap_8
XFILLER_11_910 VPWR VGND sg13g2_decap_8
XFILLER_30_707 VPWR VGND sg13g2_decap_8
XFILLER_23_781 VPWR VGND sg13g2_decap_8
XFILLER_10_464 VPWR VGND sg13g2_decap_8
XFILLER_7_936 VPWR VGND sg13g2_decap_8
XFILLER_11_987 VPWR VGND sg13g2_decap_8
XFILLER_6_446 VPWR VGND sg13g2_decap_8
XFILLER_2_630 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_49_144 VPWR VGND sg13g2_decap_8
X_41_ net1 VPWR _16_ VGND net36 _15_ sg13g2_o21ai_1
XFILLER_46_840 VPWR VGND sg13g2_decap_8
XFILLER_18_542 VPWR VGND sg13g2_decap_8
XFILLER_38_91 VPWR VGND sg13g2_decap_8
XFILLER_45_350 VPWR VGND sg13g2_decap_8
XFILLER_33_567 VPWR VGND sg13g2_decap_8
XFILLER_20_217 VPWR VGND sg13g2_decap_8
XFILLER_9_251 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_decap_8
XFILLER_37_840 VPWR VGND sg13g2_decap_8
XFILLER_24_501 VPWR VGND sg13g2_decap_8
XFILLER_36_350 VPWR VGND sg13g2_decap_8
XFILLER_24_578 VPWR VGND sg13g2_decap_8
XFILLER_34_49 VPWR VGND sg13g2_decap_8
XFILLER_11_217 VPWR VGND sg13g2_decap_8
XFILLER_20_784 VPWR VGND sg13g2_decap_8
XFILLER_4_939 VPWR VGND sg13g2_decap_8
XFILLER_3_438 VPWR VGND sg13g2_decap_8
XFILLER_8_1010 VPWR VGND sg13g2_decap_8
XFILLER_47_637 VPWR VGND sg13g2_decap_8
XFILLER_19_328 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_28_851 VPWR VGND sg13g2_decap_8
XFILLER_15_512 VPWR VGND sg13g2_decap_8
XFILLER_43_854 VPWR VGND sg13g2_decap_8
XFILLER_27_394 VPWR VGND sg13g2_decap_8
XFILLER_42_364 VPWR VGND sg13g2_decap_8
XFILLER_30_504 VPWR VGND sg13g2_decap_8
XFILLER_15_589 VPWR VGND sg13g2_decap_8
XFILLER_24_60 VPWR VGND sg13g2_decap_8
XFILLER_10_261 VPWR VGND sg13g2_decap_8
XFILLER_7_733 VPWR VGND sg13g2_decap_8
XFILLER_11_784 VPWR VGND sg13g2_decap_8
XFILLER_6_243 VPWR VGND sg13g2_decap_8
XFILLER_40_70 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_38_637 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_8
XFILLER_19_895 VPWR VGND sg13g2_decap_8
XFILLER_34_854 VPWR VGND sg13g2_decap_8
XFILLER_33_364 VPWR VGND sg13g2_decap_8
XFILLER_20_18 VPWR VGND sg13g2_decap_8
Xhold38 net9 VPWR VGND net38 sg13g2_dlygate4sd3_1
XFILLER_29_648 VPWR VGND sg13g2_decap_8
XFILLER_28_158 VPWR VGND sg13g2_decap_8
XFILLER_25_865 VPWR VGND sg13g2_decap_8
XFILLER_24_375 VPWR VGND sg13g2_decap_8
XFILLER_12_548 VPWR VGND sg13g2_decap_8
XFILLER_40_868 VPWR VGND sg13g2_decap_8
XFILLER_20_581 VPWR VGND sg13g2_decap_8
XFILLER_4_736 VPWR VGND sg13g2_decap_8
XFILLER_3_235 VPWR VGND sg13g2_decap_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
XFILLER_48_924 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_60 VPWR VGND sg13g2_decap_8
XFILLER_19_125 VPWR VGND sg13g2_decap_8
XFILLER_16_832 VPWR VGND sg13g2_decap_8
XFILLER_43_651 VPWR VGND sg13g2_decap_8
XFILLER_27_191 VPWR VGND sg13g2_decap_8
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_37_1015 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_15_386 VPWR VGND sg13g2_decap_8
XFILLER_30_301 VPWR VGND sg13g2_decap_8
XFILLER_31_868 VPWR VGND sg13g2_decap_8
XFILLER_30_378 VPWR VGND sg13g2_decap_8
XFILLER_7_530 VPWR VGND sg13g2_decap_8
XFILLER_11_581 VPWR VGND sg13g2_decap_8
XFILLER_44_1008 VPWR VGND sg13g2_decap_8
XFILLER_39_924 VPWR VGND sg13g2_decap_8
Xheichips25_template_29 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_38_434 VPWR VGND sg13g2_decap_8
XFILLER_19_692 VPWR VGND sg13g2_decap_8
XFILLER_15_18 VPWR VGND sg13g2_decap_8
XFILLER_34_651 VPWR VGND sg13g2_decap_8
XFILLER_22_835 VPWR VGND sg13g2_decap_8
XFILLER_33_161 VPWR VGND sg13g2_decap_8
XFILLER_21_367 VPWR VGND sg13g2_decap_8
XFILLER_31_28 VPWR VGND sg13g2_decap_8
Xoutput17 net17 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_728 VPWR VGND sg13g2_decap_8
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_29_445 VPWR VGND sg13g2_decap_8
XFILLER_45_938 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_decap_8
XFILLER_16_139 VPWR VGND sg13g2_decap_8
XFILLER_25_662 VPWR VGND sg13g2_decap_8
XFILLER_24_172 VPWR VGND sg13g2_decap_8
XFILLER_12_345 VPWR VGND sg13g2_decap_8
XFILLER_13_846 VPWR VGND sg13g2_decap_8
XFILLER_9_839 VPWR VGND sg13g2_decap_8
XFILLER_40_665 VPWR VGND sg13g2_decap_8
XFILLER_8_338 VPWR VGND sg13g2_decap_8
XFILLER_4_533 VPWR VGND sg13g2_decap_8
XFILLER_48_721 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_36_938 VPWR VGND sg13g2_decap_8
XFILLER_48_798 VPWR VGND sg13g2_decap_8
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_35_448 VPWR VGND sg13g2_decap_8
XFILLER_15_183 VPWR VGND sg13g2_decap_8
XFILLER_31_665 VPWR VGND sg13g2_decap_8
XFILLER_30_175 VPWR VGND sg13g2_decap_8
XFILLER_7_96 VPWR VGND sg13g2_decap_8
XFILLER_30_0 VPWR VGND sg13g2_decap_8
XFILLER_39_721 VPWR VGND sg13g2_decap_8
XFILLER_27_905 VPWR VGND sg13g2_decap_8
XFILLER_38_231 VPWR VGND sg13g2_decap_8
XFILLER_26_39 VPWR VGND sg13g2_decap_8
XFILLER_39_798 VPWR VGND sg13g2_decap_8
XFILLER_26_459 VPWR VGND sg13g2_decap_8
XFILLER_22_632 VPWR VGND sg13g2_decap_8
XFILLER_42_49 VPWR VGND sg13g2_decap_8
XFILLER_10_849 VPWR VGND sg13g2_decap_8
XFILLER_21_164 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_27_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_529 VPWR VGND sg13g2_decap_8
XFILLER_18_927 VPWR VGND sg13g2_decap_8
XFILLER_29_242 VPWR VGND sg13g2_decap_8
XFILLER_45_735 VPWR VGND sg13g2_decap_8
XFILLER_17_437 VPWR VGND sg13g2_decap_8
XFILLER_44_245 VPWR VGND sg13g2_decap_8
XFILLER_41_952 VPWR VGND sg13g2_decap_8
XFILLER_13_643 VPWR VGND sg13g2_decap_8
XFILLER_16_72 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_40_462 VPWR VGND sg13g2_decap_8
XFILLER_9_636 VPWR VGND sg13g2_decap_8
XFILLER_8_113 VPWR VGND sg13g2_fill_2
XFILLER_5_864 VPWR VGND sg13g2_decap_8
XFILLER_4_330 VPWR VGND sg13g2_decap_8
XFILLER_48_595 VPWR VGND sg13g2_decap_8
XFILLER_36_735 VPWR VGND sg13g2_decap_8
XFILLER_35_245 VPWR VGND sg13g2_decap_8
XFILLER_32_952 VPWR VGND sg13g2_decap_8
XFILLER_31_462 VPWR VGND sg13g2_decap_8
XFILLER_27_702 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_decap_8
XFILLER_39_595 VPWR VGND sg13g2_decap_8
XFILLER_27_779 VPWR VGND sg13g2_decap_8
XFILLER_14_429 VPWR VGND sg13g2_decap_8
XFILLER_26_256 VPWR VGND sg13g2_decap_8
XFILLER_42_749 VPWR VGND sg13g2_decap_8
XFILLER_23_963 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_decap_8
XFILLER_10_646 VPWR VGND sg13g2_decap_8
XFILLER_6_628 VPWR VGND sg13g2_decap_8
XFILLER_2_812 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_2_889 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_40_1022 VPWR VGND sg13g2_decap_8
XFILLER_18_724 VPWR VGND sg13g2_decap_8
XFILLER_45_532 VPWR VGND sg13g2_decap_8
XFILLER_17_234 VPWR VGND sg13g2_decap_8
XFILLER_27_93 VPWR VGND sg13g2_decap_8
XFILLER_33_749 VPWR VGND sg13g2_decap_8
XFILLER_13_440 VPWR VGND sg13g2_decap_8
XFILLER_32_259 VPWR VGND sg13g2_decap_8
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_9_433 VPWR VGND sg13g2_decap_8
XFILLER_14_996 VPWR VGND sg13g2_decap_8
XFILLER_5_661 VPWR VGND sg13g2_decap_8
XFILLER_4_20 VPWR VGND sg13g2_fill_1
XFILLER_49_893 VPWR VGND sg13g2_decap_8
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_36_532 VPWR VGND sg13g2_decap_8
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_20_966 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_39_392 VPWR VGND sg13g2_decap_8
XFILLER_27_576 VPWR VGND sg13g2_decap_8
XFILLER_42_546 VPWR VGND sg13g2_decap_8
XFILLER_14_226 VPWR VGND sg13g2_decap_8
XFILLER_23_760 VPWR VGND sg13g2_decap_8
XFILLER_10_443 VPWR VGND sg13g2_decap_8
XFILLER_7_915 VPWR VGND sg13g2_decap_8
XFILLER_11_966 VPWR VGND sg13g2_decap_8
XFILLER_6_425 VPWR VGND sg13g2_decap_8
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_2_686 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
X_40_ _09_ net39 _15_ _01_ VPWR VGND sg13g2_nor3_1
XFILLER_38_819 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
XFILLER_37_329 VPWR VGND sg13g2_decap_8
XFILLER_18_521 VPWR VGND sg13g2_decap_8
XFILLER_46_896 VPWR VGND sg13g2_decap_8
XFILLER_18_598 VPWR VGND sg13g2_decap_8
XFILLER_33_546 VPWR VGND sg13g2_decap_8
XFILLER_14_793 VPWR VGND sg13g2_decap_8
XFILLER_9_230 VPWR VGND sg13g2_decap_8
XFILLER_6_992 VPWR VGND sg13g2_decap_8
XFILLER_18_18 VPWR VGND sg13g2_decap_8
XFILLER_49_690 VPWR VGND sg13g2_decap_8
XFILLER_34_28 VPWR VGND sg13g2_decap_8
XFILLER_37_896 VPWR VGND sg13g2_decap_8
XFILLER_24_557 VPWR VGND sg13g2_decap_8
XFILLER_20_763 VPWR VGND sg13g2_decap_8
XFILLER_4_918 VPWR VGND sg13g2_decap_8
XFILLER_3_417 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_47_616 VPWR VGND sg13g2_decap_8
XFILLER_19_307 VPWR VGND sg13g2_decap_8
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_28_830 VPWR VGND sg13g2_decap_8
XFILLER_43_833 VPWR VGND sg13g2_decap_8
XFILLER_27_373 VPWR VGND sg13g2_decap_8
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_15_568 VPWR VGND sg13g2_decap_8
XFILLER_10_240 VPWR VGND sg13g2_decap_8
XFILLER_7_712 VPWR VGND sg13g2_decap_8
XFILLER_11_763 VPWR VGND sg13g2_decap_8
XFILLER_6_222 VPWR VGND sg13g2_decap_8
XFILLER_7_789 VPWR VGND sg13g2_decap_8
XFILLER_6_299 VPWR VGND sg13g2_decap_8
XFILLER_3_984 VPWR VGND sg13g2_decap_8
XFILLER_2_483 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_38_616 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_19_874 VPWR VGND sg13g2_decap_8
XFILLER_46_693 VPWR VGND sg13g2_decap_8
XFILLER_18_395 VPWR VGND sg13g2_decap_8
XFILLER_34_833 VPWR VGND sg13g2_decap_8
XFILLER_33_343 VPWR VGND sg13g2_decap_8
XFILLER_14_590 VPWR VGND sg13g2_decap_8
XFILLER_21_549 VPWR VGND sg13g2_decap_8
XFILLER_29_39 VPWR VGND sg13g2_decap_8
Xhold39 _14_ VPWR VGND net39 sg13g2_dlygate4sd3_1
XFILLER_29_627 VPWR VGND sg13g2_decap_8
XFILLER_28_137 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_8
XFILLER_25_844 VPWR VGND sg13g2_decap_8
XFILLER_37_693 VPWR VGND sg13g2_decap_8
XFILLER_24_354 VPWR VGND sg13g2_decap_8
XFILLER_12_527 VPWR VGND sg13g2_decap_8
XFILLER_40_847 VPWR VGND sg13g2_decap_8
XFILLER_20_560 VPWR VGND sg13g2_decap_8
XFILLER_4_715 VPWR VGND sg13g2_decap_8
XFILLER_3_214 VPWR VGND sg13g2_decap_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_48_903 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_16_811 VPWR VGND sg13g2_decap_8
XFILLER_27_170 VPWR VGND sg13g2_decap_8
XFILLER_43_630 VPWR VGND sg13g2_decap_8
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_15_365 VPWR VGND sg13g2_decap_8
XFILLER_16_888 VPWR VGND sg13g2_decap_8
XFILLER_31_847 VPWR VGND sg13g2_decap_8
XFILLER_11_560 VPWR VGND sg13g2_decap_8
XFILLER_30_357 VPWR VGND sg13g2_decap_8
XFILLER_7_586 VPWR VGND sg13g2_decap_8
XFILLER_3_781 VPWR VGND sg13g2_decap_8
XFILLER_2_280 VPWR VGND sg13g2_decap_8
XFILLER_39_903 VPWR VGND sg13g2_decap_8
XFILLER_38_413 VPWR VGND sg13g2_decap_8
XFILLER_47_980 VPWR VGND sg13g2_decap_8
XFILLER_19_671 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
XFILLER_18_192 VPWR VGND sg13g2_decap_8
XFILLER_34_630 VPWR VGND sg13g2_decap_8
XFILLER_22_814 VPWR VGND sg13g2_decap_8
XFILLER_33_140 VPWR VGND sg13g2_decap_8
XFILLER_21_346 VPWR VGND sg13g2_decap_8
Xoutput18 net18 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_707 VPWR VGND sg13g2_decap_8
XFILLER_0_217 VPWR VGND sg13g2_decap_8
XFILLER_5_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_424 VPWR VGND sg13g2_decap_8
XFILLER_45_917 VPWR VGND sg13g2_decap_8
XFILLER_17_619 VPWR VGND sg13g2_decap_8
XFILLER_44_427 VPWR VGND sg13g2_decap_8
XFILLER_16_118 VPWR VGND sg13g2_decap_8
XFILLER_38_980 VPWR VGND sg13g2_decap_8
XFILLER_25_641 VPWR VGND sg13g2_decap_8
XFILLER_37_490 VPWR VGND sg13g2_decap_8
XFILLER_13_825 VPWR VGND sg13g2_decap_8
XFILLER_24_151 VPWR VGND sg13g2_decap_8
XFILLER_9_818 VPWR VGND sg13g2_decap_8
XFILLER_12_324 VPWR VGND sg13g2_decap_8
XFILLER_40_644 VPWR VGND sg13g2_decap_8
XFILLER_8_317 VPWR VGND sg13g2_decap_8
XFILLER_4_512 VPWR VGND sg13g2_decap_8
XFILLER_4_589 VPWR VGND sg13g2_decap_8
XFILLER_48_700 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_48_777 VPWR VGND sg13g2_decap_8
XFILLER_36_917 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_29_991 VPWR VGND sg13g2_decap_8
XFILLER_35_427 VPWR VGND sg13g2_decap_8
XFILLER_44_994 VPWR VGND sg13g2_decap_8
XFILLER_15_162 VPWR VGND sg13g2_decap_8
XFILLER_16_685 VPWR VGND sg13g2_decap_8
XFILLER_31_644 VPWR VGND sg13g2_decap_8
XFILLER_30_154 VPWR VGND sg13g2_decap_8
XFILLER_12_891 VPWR VGND sg13g2_decap_8
XFILLER_11_1008 VPWR VGND sg13g2_decap_8
XFILLER_8_884 VPWR VGND sg13g2_decap_8
XFILLER_7_383 VPWR VGND sg13g2_decap_8
XFILLER_7_75 VPWR VGND sg13g2_decap_8
XFILLER_39_700 VPWR VGND sg13g2_decap_8
XFILLER_38_210 VPWR VGND sg13g2_decap_8
XFILLER_39_777 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_fill_2
XFILLER_26_438 VPWR VGND sg13g2_decap_8
XFILLER_38_287 VPWR VGND sg13g2_decap_8
XFILLER_22_611 VPWR VGND sg13g2_decap_8
XFILLER_35_994 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_21_143 VPWR VGND sg13g2_decap_8
XFILLER_10_828 VPWR VGND sg13g2_decap_8
XFILLER_22_688 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_29_221 VPWR VGND sg13g2_decap_8
XFILLER_18_906 VPWR VGND sg13g2_decap_8
XFILLER_45_714 VPWR VGND sg13g2_decap_8
XFILLER_17_416 VPWR VGND sg13g2_decap_8
XFILLER_44_224 VPWR VGND sg13g2_decap_8
XFILLER_29_298 VPWR VGND sg13g2_decap_8
XFILLER_16_51 VPWR VGND sg13g2_decap_8
XFILLER_41_931 VPWR VGND sg13g2_decap_8
XFILLER_13_622 VPWR VGND sg13g2_decap_8
XFILLER_9_615 VPWR VGND sg13g2_decap_8
XFILLER_34_1008 VPWR VGND sg13g2_decap_8
XFILLER_40_441 VPWR VGND sg13g2_decap_8
XFILLER_13_699 VPWR VGND sg13g2_decap_8
XFILLER_12_198 VPWR VGND sg13g2_decap_8
XFILLER_5_843 VPWR VGND sg13g2_decap_8
XFILLER_4_386 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_48_574 VPWR VGND sg13g2_decap_8
XFILLER_36_714 VPWR VGND sg13g2_decap_8
XFILLER_35_224 VPWR VGND sg13g2_decap_8
XFILLER_17_983 VPWR VGND sg13g2_decap_8
XFILLER_44_791 VPWR VGND sg13g2_decap_8
XFILLER_16_482 VPWR VGND sg13g2_decap_8
XFILLER_32_931 VPWR VGND sg13g2_decap_8
XFILLER_31_441 VPWR VGND sg13g2_decap_8
X_56__23 VPWR VGND net22 sg13g2_tiehi
XFILLER_8_681 VPWR VGND sg13g2_decap_8
XFILLER_7_180 VPWR VGND sg13g2_decap_8
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_39_574 VPWR VGND sg13g2_decap_8
XFILLER_26_235 VPWR VGND sg13g2_decap_8
XFILLER_27_758 VPWR VGND sg13g2_decap_8
XFILLER_42_728 VPWR VGND sg13g2_decap_8
XFILLER_14_408 VPWR VGND sg13g2_decap_8
XFILLER_23_942 VPWR VGND sg13g2_decap_8
XFILLER_35_791 VPWR VGND sg13g2_decap_8
XFILLER_41_238 VPWR VGND sg13g2_decap_8
XFILLER_10_625 VPWR VGND sg13g2_decap_8
XFILLER_22_485 VPWR VGND sg13g2_decap_8
XFILLER_6_607 VPWR VGND sg13g2_decap_8
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_2_868 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_40_1001 VPWR VGND sg13g2_decap_8
XFILLER_45_511 VPWR VGND sg13g2_decap_8
XFILLER_18_703 VPWR VGND sg13g2_decap_8
XFILLER_17_213 VPWR VGND sg13g2_decap_8
XFILLER_27_72 VPWR VGND sg13g2_decap_8
XFILLER_45_588 VPWR VGND sg13g2_decap_8
XFILLER_33_728 VPWR VGND sg13g2_decap_8
XFILLER_32_238 VPWR VGND sg13g2_decap_8
XFILLER_14_975 VPWR VGND sg13g2_decap_8
XFILLER_9_412 VPWR VGND sg13g2_decap_8
XFILLER_13_496 VPWR VGND sg13g2_decap_8
XFILLER_9_489 VPWR VGND sg13g2_decap_8
XFILLER_5_640 VPWR VGND sg13g2_decap_8
XFILLER_4_183 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_4
XFILLER_49_872 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_36_511 VPWR VGND sg13g2_decap_8
XFILLER_36_588 VPWR VGND sg13g2_decap_8
XFILLER_17_780 VPWR VGND sg13g2_decap_8
XFILLER_24_739 VPWR VGND sg13g2_decap_8
XFILLER_23_249 VPWR VGND sg13g2_decap_8
XFILLER_17_1025 VPWR VGND sg13g2_decap_4
XFILLER_20_945 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_39_371 VPWR VGND sg13g2_decap_8
XFILLER_27_555 VPWR VGND sg13g2_decap_8
XFILLER_42_525 VPWR VGND sg13g2_decap_8
XFILLER_14_205 VPWR VGND sg13g2_decap_8
XFILLER_10_422 VPWR VGND sg13g2_decap_8
XFILLER_11_945 VPWR VGND sg13g2_decap_8
XFILLER_22_282 VPWR VGND sg13g2_decap_8
XFILLER_6_404 VPWR VGND sg13g2_decap_8
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_10_499 VPWR VGND sg13g2_decap_8
XFILLER_2_665 VPWR VGND sg13g2_decap_8
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_18_500 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_decap_8
XFILLER_46_875 VPWR VGND sg13g2_decap_8
XFILLER_18_577 VPWR VGND sg13g2_decap_8
XFILLER_45_385 VPWR VGND sg13g2_decap_8
XFILLER_33_525 VPWR VGND sg13g2_decap_8
XFILLER_14_772 VPWR VGND sg13g2_decap_8
XFILLER_13_293 VPWR VGND sg13g2_decap_8
XFILLER_9_286 VPWR VGND sg13g2_decap_8
XFILLER_6_971 VPWR VGND sg13g2_decap_8
XFILLER_29_809 VPWR VGND sg13g2_decap_8
XFILLER_28_319 VPWR VGND sg13g2_decap_8
XFILLER_37_875 VPWR VGND sg13g2_decap_8
XFILLER_24_536 VPWR VGND sg13g2_decap_8
XFILLER_36_385 VPWR VGND sg13g2_decap_8
XFILLER_12_709 VPWR VGND sg13g2_decap_8
XFILLER_20_742 VPWR VGND sg13g2_decap_8
XFILLER_30_1022 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_43_812 VPWR VGND sg13g2_decap_8
XFILLER_27_352 VPWR VGND sg13g2_decap_8
XFILLER_28_886 VPWR VGND sg13g2_decap_8
XFILLER_42_322 VPWR VGND sg13g2_decap_8
XFILLER_15_547 VPWR VGND sg13g2_decap_8
XFILLER_43_889 VPWR VGND sg13g2_decap_8
XFILLER_42_399 VPWR VGND sg13g2_decap_8
XFILLER_11_742 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_decap_8
XFILLER_6_201 VPWR VGND sg13g2_decap_8
XFILLER_24_95 VPWR VGND sg13g2_decap_8
XFILLER_7_768 VPWR VGND sg13g2_decap_8
XFILLER_10_296 VPWR VGND sg13g2_decap_8
XFILLER_6_278 VPWR VGND sg13g2_decap_8
XFILLER_3_963 VPWR VGND sg13g2_decap_8
XFILLER_2_462 VPWR VGND sg13g2_decap_8
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_19_853 VPWR VGND sg13g2_decap_8
XFILLER_46_672 VPWR VGND sg13g2_decap_8
XFILLER_18_374 VPWR VGND sg13g2_decap_8
XFILLER_34_812 VPWR VGND sg13g2_decap_8
XFILLER_45_182 VPWR VGND sg13g2_decap_8
XFILLER_33_322 VPWR VGND sg13g2_decap_8
XFILLER_21_528 VPWR VGND sg13g2_decap_8
XFILLER_34_889 VPWR VGND sg13g2_decap_8
XFILLER_33_399 VPWR VGND sg13g2_decap_8
XFILLER_14_1017 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_18 VPWR VGND sg13g2_decap_8
XFILLER_29_606 VPWR VGND sg13g2_decap_8
XFILLER_28_116 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_44_609 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_25_823 VPWR VGND sg13g2_decap_8
XFILLER_37_672 VPWR VGND sg13g2_decap_8
XFILLER_24_333 VPWR VGND sg13g2_decap_8
XFILLER_36_182 VPWR VGND sg13g2_decap_8
XFILLER_12_506 VPWR VGND sg13g2_decap_8
XFILLER_40_826 VPWR VGND sg13g2_decap_8
XFILLER_10_64 VPWR VGND sg13g2_fill_1
XFILLER_10_53 VPWR VGND sg13g2_decap_8
XFILLER_10_86 VPWR VGND sg13g2_decap_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_48_959 VPWR VGND sg13g2_decap_8
Xheichips25_template VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_35_609 VPWR VGND sg13g2_decap_8
XFILLER_28_683 VPWR VGND sg13g2_decap_8
XFILLER_34_119 VPWR VGND sg13g2_decap_8
XFILLER_15_344 VPWR VGND sg13g2_decap_8
XFILLER_16_867 VPWR VGND sg13g2_decap_8
XFILLER_43_686 VPWR VGND sg13g2_decap_8
XFILLER_31_826 VPWR VGND sg13g2_decap_8
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_30_336 VPWR VGND sg13g2_decap_8
XFILLER_7_565 VPWR VGND sg13g2_decap_8
XFILLER_3_760 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_39_959 VPWR VGND sg13g2_decap_8
XFILLER_19_650 VPWR VGND sg13g2_decap_8
XFILLER_38_469 VPWR VGND sg13g2_decap_8
XFILLER_18_171 VPWR VGND sg13g2_decap_8
XFILLER_34_686 VPWR VGND sg13g2_decap_8
XFILLER_21_325 VPWR VGND sg13g2_decap_8
XFILLER_33_196 VPWR VGND sg13g2_decap_8
XFILLER_5_1004 VPWR VGND sg13g2_decap_8
XFILLER_29_403 VPWR VGND sg13g2_decap_8
XFILLER_44_406 VPWR VGND sg13g2_decap_8
XFILLER_25_620 VPWR VGND sg13g2_decap_8
XFILLER_12_303 VPWR VGND sg13g2_decap_8
XFILLER_13_804 VPWR VGND sg13g2_decap_8
XFILLER_24_130 VPWR VGND sg13g2_decap_8
XFILLER_25_697 VPWR VGND sg13g2_decap_8
XFILLER_40_623 VPWR VGND sg13g2_decap_8
XFILLER_21_892 VPWR VGND sg13g2_decap_8
XFILLER_4_568 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_29_970 VPWR VGND sg13g2_decap_8
XFILLER_35_406 VPWR VGND sg13g2_decap_8
XFILLER_28_480 VPWR VGND sg13g2_decap_8
XFILLER_44_973 VPWR VGND sg13g2_decap_8
XFILLER_15_141 VPWR VGND sg13g2_decap_8
XFILLER_16_664 VPWR VGND sg13g2_decap_8
XFILLER_43_483 VPWR VGND sg13g2_decap_8
XFILLER_31_623 VPWR VGND sg13g2_decap_8
XFILLER_30_133 VPWR VGND sg13g2_decap_8
XFILLER_12_870 VPWR VGND sg13g2_decap_8
XFILLER_8_863 VPWR VGND sg13g2_decap_8
XFILLER_7_54 VPWR VGND sg13g2_decap_8
XFILLER_7_32 VPWR VGND sg13g2_decap_8
XFILLER_7_362 VPWR VGND sg13g2_decap_8
XFILLER_39_756 VPWR VGND sg13g2_decap_8
XFILLER_26_417 VPWR VGND sg13g2_decap_8
XFILLER_38_266 VPWR VGND sg13g2_decap_8
XFILLER_35_973 VPWR VGND sg13g2_decap_8
XFILLER_34_483 VPWR VGND sg13g2_decap_8
XFILLER_10_807 VPWR VGND sg13g2_decap_8
XFILLER_21_122 VPWR VGND sg13g2_decap_8
XFILLER_22_667 VPWR VGND sg13g2_decap_8
XFILLER_21_199 VPWR VGND sg13g2_decap_8
XFILLER_29_200 VPWR VGND sg13g2_decap_8
XFILLER_44_203 VPWR VGND sg13g2_decap_8
XFILLER_29_277 VPWR VGND sg13g2_decap_8
XFILLER_41_910 VPWR VGND sg13g2_decap_8
XFILLER_13_601 VPWR VGND sg13g2_decap_8
XFILLER_26_984 VPWR VGND sg13g2_decap_8
XFILLER_25_494 VPWR VGND sg13g2_decap_8
XFILLER_40_420 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_fill_1
XFILLER_41_987 VPWR VGND sg13g2_decap_8
XFILLER_12_177 VPWR VGND sg13g2_decap_8
XFILLER_13_678 VPWR VGND sg13g2_decap_8
XFILLER_40_497 VPWR VGND sg13g2_decap_8
XFILLER_5_822 VPWR VGND sg13g2_decap_8
XFILLER_32_84 VPWR VGND sg13g2_decap_8
XFILLER_5_899 VPWR VGND sg13g2_decap_8
XFILLER_4_365 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_17_962 VPWR VGND sg13g2_decap_8
XFILLER_32_910 VPWR VGND sg13g2_decap_8
XFILLER_44_770 VPWR VGND sg13g2_decap_8
XFILLER_16_461 VPWR VGND sg13g2_decap_8
XFILLER_31_420 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
XFILLER_32_987 VPWR VGND sg13g2_decap_8
XFILLER_31_497 VPWR VGND sg13g2_decap_8
XFILLER_8_660 VPWR VGND sg13g2_decap_8
XFILLER_39_553 VPWR VGND sg13g2_decap_8
XFILLER_26_214 VPWR VGND sg13g2_decap_8
XFILLER_27_737 VPWR VGND sg13g2_decap_8
XFILLER_42_707 VPWR VGND sg13g2_decap_8
XFILLER_23_921 VPWR VGND sg13g2_decap_8
XFILLER_35_770 VPWR VGND sg13g2_decap_8
XFILLER_41_217 VPWR VGND sg13g2_decap_8
XFILLER_34_280 VPWR VGND sg13g2_decap_8
XFILLER_10_604 VPWR VGND sg13g2_decap_8
XFILLER_22_464 VPWR VGND sg13g2_decap_8
XFILLER_23_998 VPWR VGND sg13g2_decap_8
XFILLER_5_129 VPWR VGND sg13g2_decap_8
XFILLER_2_847 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_18_759 VPWR VGND sg13g2_decap_8
XFILLER_45_567 VPWR VGND sg13g2_decap_8
XFILLER_17_269 VPWR VGND sg13g2_decap_8
XFILLER_33_707 VPWR VGND sg13g2_decap_8
XFILLER_26_781 VPWR VGND sg13g2_decap_8
XFILLER_32_217 VPWR VGND sg13g2_decap_8
XFILLER_14_954 VPWR VGND sg13g2_decap_8
XFILLER_25_291 VPWR VGND sg13g2_decap_8
XFILLER_41_784 VPWR VGND sg13g2_decap_8
XFILLER_13_475 VPWR VGND sg13g2_decap_8
XFILLER_9_468 VPWR VGND sg13g2_decap_8
XFILLER_40_294 VPWR VGND sg13g2_decap_8
XFILLER_5_696 VPWR VGND sg13g2_decap_8
XFILLER_4_162 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_77 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_fill_2
XFILLER_49_851 VPWR VGND sg13g2_decap_8
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_24_718 VPWR VGND sg13g2_decap_8
XFILLER_36_567 VPWR VGND sg13g2_decap_8
XFILLER_23_228 VPWR VGND sg13g2_decap_8
XFILLER_17_1004 VPWR VGND sg13g2_decap_8
XFILLER_20_924 VPWR VGND sg13g2_decap_8
XFILLER_32_784 VPWR VGND sg13g2_decap_8
XFILLER_31_294 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_24_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_350 VPWR VGND sg13g2_decap_8
XFILLER_27_534 VPWR VGND sg13g2_decap_8
XFILLER_42_504 VPWR VGND sg13g2_decap_8
XFILLER_15_729 VPWR VGND sg13g2_decap_8
XFILLER_10_401 VPWR VGND sg13g2_decap_8
XFILLER_11_924 VPWR VGND sg13g2_decap_8
XFILLER_22_261 VPWR VGND sg13g2_decap_8
XFILLER_23_795 VPWR VGND sg13g2_decap_8
XFILLER_10_478 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_2_644 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_46_854 VPWR VGND sg13g2_decap_8
XFILLER_18_556 VPWR VGND sg13g2_decap_8
XFILLER_33_504 VPWR VGND sg13g2_decap_8
XFILLER_45_364 VPWR VGND sg13g2_decap_8
XFILLER_14_751 VPWR VGND sg13g2_decap_8
XFILLER_41_581 VPWR VGND sg13g2_decap_8
XFILLER_13_272 VPWR VGND sg13g2_decap_8
XFILLER_9_265 VPWR VGND sg13g2_decap_8
XFILLER_6_950 VPWR VGND sg13g2_decap_8
XFILLER_47_1008 VPWR VGND sg13g2_decap_8
XFILLER_5_493 VPWR VGND sg13g2_decap_8
XFILLER_37_854 VPWR VGND sg13g2_decap_8
XFILLER_24_515 VPWR VGND sg13g2_decap_8
XFILLER_36_364 VPWR VGND sg13g2_decap_8
XFILLER_20_721 VPWR VGND sg13g2_decap_8
XFILLER_32_581 VPWR VGND sg13g2_decap_8
XFILLER_30_1001 VPWR VGND sg13g2_decap_8
XFILLER_20_798 VPWR VGND sg13g2_decap_8
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
XFILLER_27_331 VPWR VGND sg13g2_decap_8
XFILLER_28_865 VPWR VGND sg13g2_decap_8
XFILLER_42_301 VPWR VGND sg13g2_decap_8
XFILLER_15_526 VPWR VGND sg13g2_decap_8
XFILLER_43_868 VPWR VGND sg13g2_decap_8
XFILLER_42_378 VPWR VGND sg13g2_decap_8
XFILLER_30_518 VPWR VGND sg13g2_decap_8
XFILLER_11_721 VPWR VGND sg13g2_decap_8
XFILLER_23_592 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_decap_8
XFILLER_10_275 VPWR VGND sg13g2_decap_8
XFILLER_7_747 VPWR VGND sg13g2_decap_8
XFILLER_11_798 VPWR VGND sg13g2_decap_8
XFILLER_6_257 VPWR VGND sg13g2_decap_8
XFILLER_40_84 VPWR VGND sg13g2_decap_8
XFILLER_3_942 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_8
XFILLER_49_60 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_832 VPWR VGND sg13g2_decap_8
XFILLER_46_651 VPWR VGND sg13g2_decap_8
XFILLER_18_353 VPWR VGND sg13g2_decap_8
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_33_301 VPWR VGND sg13g2_decap_8
XFILLER_34_868 VPWR VGND sg13g2_decap_8
XFILLER_21_507 VPWR VGND sg13g2_decap_8
XFILLER_33_378 VPWR VGND sg13g2_decap_8
XFILLER_46_0 VPWR VGND sg13g2_decap_8
XFILLER_5_290 VPWR VGND sg13g2_decap_8
XFILLER_25_802 VPWR VGND sg13g2_decap_8
XFILLER_37_651 VPWR VGND sg13g2_decap_8
XFILLER_36_161 VPWR VGND sg13g2_decap_8
XFILLER_24_312 VPWR VGND sg13g2_decap_8
XFILLER_25_879 VPWR VGND sg13g2_decap_8
XFILLER_40_805 VPWR VGND sg13g2_decap_8
XFILLER_24_389 VPWR VGND sg13g2_decap_8
XFILLER_20_595 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_decap_8
XFILLER_3_249 VPWR VGND sg13g2_decap_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
XFILLER_48_938 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_19_85 VPWR VGND sg13g2_fill_1
XFILLER_19_139 VPWR VGND sg13g2_decap_8
XFILLER_28_662 VPWR VGND sg13g2_decap_8
XFILLER_15_323 VPWR VGND sg13g2_decap_8
XFILLER_16_846 VPWR VGND sg13g2_decap_8
XFILLER_43_665 VPWR VGND sg13g2_decap_8
XFILLER_31_805 VPWR VGND sg13g2_decap_8
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_42_175 VPWR VGND sg13g2_decap_8
XFILLER_30_315 VPWR VGND sg13g2_decap_8
XFILLER_7_544 VPWR VGND sg13g2_decap_8
XFILLER_11_595 VPWR VGND sg13g2_decap_8
XFILLER_18_4 VPWR VGND sg13g2_decap_8
XFILLER_39_938 VPWR VGND sg13g2_decap_8
XFILLER_20_1022 VPWR VGND sg13g2_decap_8
XFILLER_38_448 VPWR VGND sg13g2_decap_8
XFILLER_25_109 VPWR VGND sg13g2_decap_8
XFILLER_34_665 VPWR VGND sg13g2_decap_8
XFILLER_15_890 VPWR VGND sg13g2_decap_8
XFILLER_21_304 VPWR VGND sg13g2_decap_8
XFILLER_22_849 VPWR VGND sg13g2_decap_8
XFILLER_33_175 VPWR VGND sg13g2_decap_8
XFILLER_30_882 VPWR VGND sg13g2_decap_8
XFILLER_29_459 VPWR VGND sg13g2_decap_8
XFILLER_25_676 VPWR VGND sg13g2_decap_8
XFILLER_40_602 VPWR VGND sg13g2_decap_8
XFILLER_24_186 VPWR VGND sg13g2_decap_8
XFILLER_12_359 VPWR VGND sg13g2_decap_8
XFILLER_40_679 VPWR VGND sg13g2_decap_8
XFILLER_21_871 VPWR VGND sg13g2_decap_8
XFILLER_20_392 VPWR VGND sg13g2_decap_8
XFILLER_21_53 VPWR VGND sg13g2_decap_8
XFILLER_4_547 VPWR VGND sg13g2_decap_8
XFILLER_43_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_48_735 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_44_952 VPWR VGND sg13g2_decap_8
XFILLER_16_643 VPWR VGND sg13g2_decap_8
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_15_120 VPWR VGND sg13g2_decap_8
XFILLER_31_602 VPWR VGND sg13g2_decap_8
XFILLER_30_112 VPWR VGND sg13g2_decap_8
XFILLER_15_197 VPWR VGND sg13g2_decap_8
XFILLER_31_679 VPWR VGND sg13g2_decap_8
XFILLER_8_842 VPWR VGND sg13g2_decap_8
XFILLER_7_341 VPWR VGND sg13g2_decap_8
XFILLER_11_392 VPWR VGND sg13g2_decap_8
XFILLER_30_189 VPWR VGND sg13g2_decap_8
XFILLER_39_735 VPWR VGND sg13g2_decap_8
XFILLER_27_919 VPWR VGND sg13g2_decap_8
XFILLER_38_245 VPWR VGND sg13g2_decap_8
XFILLER_35_952 VPWR VGND sg13g2_decap_8
XFILLER_21_101 VPWR VGND sg13g2_decap_8
XFILLER_34_462 VPWR VGND sg13g2_decap_8
XFILLER_22_646 VPWR VGND sg13g2_decap_8
XFILLER_21_178 VPWR VGND sg13g2_decap_8
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_27_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_256 VPWR VGND sg13g2_decap_8
XFILLER_45_749 VPWR VGND sg13g2_decap_8
XFILLER_44_259 VPWR VGND sg13g2_decap_8
XFILLER_26_963 VPWR VGND sg13g2_decap_8
XFILLER_16_86 VPWR VGND sg13g2_decap_8
XFILLER_25_473 VPWR VGND sg13g2_decap_8
XFILLER_41_966 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_decap_8
XFILLER_13_657 VPWR VGND sg13g2_decap_8
XFILLER_16_97 VPWR VGND sg13g2_fill_2
XFILLER_12_156 VPWR VGND sg13g2_decap_8
XFILLER_40_476 VPWR VGND sg13g2_decap_8
XFILLER_8_149 VPWR VGND sg13g2_decap_8
XFILLER_32_63 VPWR VGND sg13g2_decap_8
XFILLER_5_801 VPWR VGND sg13g2_decap_8
XFILLER_10_1010 VPWR VGND sg13g2_decap_8
XFILLER_5_878 VPWR VGND sg13g2_decap_8
XFILLER_4_344 VPWR VGND sg13g2_decap_8
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_17_941 VPWR VGND sg13g2_decap_8
XFILLER_36_749 VPWR VGND sg13g2_decap_8
XFILLER_16_440 VPWR VGND sg13g2_decap_8
XFILLER_35_259 VPWR VGND sg13g2_decap_8
XFILLER_32_966 VPWR VGND sg13g2_decap_8
XFILLER_31_476 VPWR VGND sg13g2_decap_8
XFILLER_39_532 VPWR VGND sg13g2_decap_8
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
XFILLER_27_716 VPWR VGND sg13g2_decap_8
XFILLER_23_900 VPWR VGND sg13g2_decap_8
XFILLER_22_443 VPWR VGND sg13g2_decap_8
XFILLER_23_977 VPWR VGND sg13g2_decap_8
XFILLER_5_108 VPWR VGND sg13g2_decap_8
XFILLER_2_826 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_45_546 VPWR VGND sg13g2_decap_8
XFILLER_18_738 VPWR VGND sg13g2_decap_8
XFILLER_17_248 VPWR VGND sg13g2_decap_8
XFILLER_14_933 VPWR VGND sg13g2_decap_8
XFILLER_26_760 VPWR VGND sg13g2_decap_8
XFILLER_25_270 VPWR VGND sg13g2_decap_8
XFILLER_41_763 VPWR VGND sg13g2_decap_8
XFILLER_13_454 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_9_447 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_decap_8
XFILLER_5_675 VPWR VGND sg13g2_decap_8
XFILLER_4_141 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_4_45 VPWR VGND sg13g2_fill_2
XFILLER_49_830 VPWR VGND sg13g2_decap_8
XFILLER_36_546 VPWR VGND sg13g2_decap_8
XFILLER_23_207 VPWR VGND sg13g2_decap_8
XFILLER_20_903 VPWR VGND sg13g2_decap_8
XFILLER_32_763 VPWR VGND sg13g2_decap_8
XFILLER_31_273 VPWR VGND sg13g2_decap_8
XFILLER_27_513 VPWR VGND sg13g2_decap_8
XFILLER_15_708 VPWR VGND sg13g2_decap_8
XFILLER_11_903 VPWR VGND sg13g2_decap_8
XFILLER_22_240 VPWR VGND sg13g2_decap_8
XFILLER_23_774 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
XFILLER_10_457 VPWR VGND sg13g2_decap_8
XFILLER_7_929 VPWR VGND sg13g2_decap_8
XFILLER_6_439 VPWR VGND sg13g2_decap_8
XFILLER_2_623 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_46_833 VPWR VGND sg13g2_decap_8
XFILLER_18_535 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_14_730 VPWR VGND sg13g2_decap_8
XFILLER_41_560 VPWR VGND sg13g2_decap_8
XFILLER_13_251 VPWR VGND sg13g2_decap_8
XFILLER_9_244 VPWR VGND sg13g2_decap_8
XFILLER_5_472 VPWR VGND sg13g2_decap_8
XFILLER_37_833 VPWR VGND sg13g2_decap_8
XFILLER_36_343 VPWR VGND sg13g2_decap_8
XFILLER_20_700 VPWR VGND sg13g2_decap_8
XFILLER_32_560 VPWR VGND sg13g2_decap_8
XFILLER_20_777 VPWR VGND sg13g2_decap_8
XFILLER_8_1003 VPWR VGND sg13g2_decap_8
XFILLER_27_310 VPWR VGND sg13g2_decap_8
XFILLER_28_844 VPWR VGND sg13g2_decap_8
XFILLER_15_505 VPWR VGND sg13g2_decap_8
XFILLER_27_387 VPWR VGND sg13g2_decap_8
XFILLER_43_847 VPWR VGND sg13g2_decap_8
XFILLER_42_357 VPWR VGND sg13g2_decap_8
XFILLER_11_700 VPWR VGND sg13g2_decap_8
XFILLER_23_571 VPWR VGND sg13g2_decap_8
XFILLER_24_53 VPWR VGND sg13g2_decap_8
XFILLER_10_254 VPWR VGND sg13g2_decap_8
XFILLER_7_726 VPWR VGND sg13g2_decap_8
XFILLER_11_777 VPWR VGND sg13g2_decap_8
XFILLER_6_236 VPWR VGND sg13g2_decap_8
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_3_921 VPWR VGND sg13g2_decap_8
XFILLER_2_420 VPWR VGND sg13g2_decap_8
XFILLER_3_998 VPWR VGND sg13g2_decap_8
XFILLER_2_497 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_19_811 VPWR VGND sg13g2_decap_8
XFILLER_46_630 VPWR VGND sg13g2_decap_8
XFILLER_18_332 VPWR VGND sg13g2_decap_8
XFILLER_45_140 VPWR VGND sg13g2_decap_8
XFILLER_19_888 VPWR VGND sg13g2_decap_8
XFILLER_34_847 VPWR VGND sg13g2_decap_8
XFILLER_33_357 VPWR VGND sg13g2_decap_8
XFILLER_39_0 VPWR VGND sg13g2_decap_8
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
XFILLER_37_630 VPWR VGND sg13g2_decap_8
XFILLER_36_140 VPWR VGND sg13g2_decap_8
XFILLER_25_858 VPWR VGND sg13g2_decap_8
XFILLER_24_368 VPWR VGND sg13g2_decap_8
XFILLER_20_574 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_4
XFILLER_4_729 VPWR VGND sg13g2_decap_8
XFILLER_3_228 VPWR VGND sg13g2_decap_8
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_48_917 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_8
XFILLER_19_118 VPWR VGND sg13g2_decap_8
XFILLER_28_641 VPWR VGND sg13g2_decap_8
XFILLER_15_302 VPWR VGND sg13g2_decap_8
XFILLER_16_825 VPWR VGND sg13g2_decap_8
XFILLER_43_644 VPWR VGND sg13g2_decap_8
XFILLER_27_184 VPWR VGND sg13g2_decap_8
XFILLER_42_154 VPWR VGND sg13g2_decap_8
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_37_1008 VPWR VGND sg13g2_decap_8
XFILLER_15_379 VPWR VGND sg13g2_decap_8
XFILLER_7_523 VPWR VGND sg13g2_decap_8
XFILLER_11_574 VPWR VGND sg13g2_decap_8
XFILLER_3_795 VPWR VGND sg13g2_decap_8
XFILLER_32_7 VPWR VGND sg13g2_decap_8
XFILLER_2_294 VPWR VGND sg13g2_decap_8
XFILLER_39_917 VPWR VGND sg13g2_decap_8
XFILLER_38_427 VPWR VGND sg13g2_decap_8
XFILLER_20_1001 VPWR VGND sg13g2_decap_8
XFILLER_47_994 VPWR VGND sg13g2_decap_8
XFILLER_19_685 VPWR VGND sg13g2_decap_8
XFILLER_34_644 VPWR VGND sg13g2_decap_8
XFILLER_33_154 VPWR VGND sg13g2_decap_8
XFILLER_22_828 VPWR VGND sg13g2_decap_8
XFILLER_30_861 VPWR VGND sg13g2_decap_8
XFILLER_29_438 VPWR VGND sg13g2_decap_8
XFILLER_38_994 VPWR VGND sg13g2_decap_8
XFILLER_25_655 VPWR VGND sg13g2_decap_8
XFILLER_13_839 VPWR VGND sg13g2_decap_8
XFILLER_24_165 VPWR VGND sg13g2_decap_8
XFILLER_12_338 VPWR VGND sg13g2_decap_8
XFILLER_21_850 VPWR VGND sg13g2_decap_8
XFILLER_40_658 VPWR VGND sg13g2_decap_8
XFILLER_20_371 VPWR VGND sg13g2_decap_8
XFILLER_21_32 VPWR VGND sg13g2_decap_8
XFILLER_4_526 VPWR VGND sg13g2_decap_8
XFILLER_21_87 VPWR VGND sg13g2_decap_4
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_43_1001 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_44_931 VPWR VGND sg13g2_decap_8
XFILLER_16_622 VPWR VGND sg13g2_decap_8
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_15_176 VPWR VGND sg13g2_decap_8
XFILLER_16_699 VPWR VGND sg13g2_decap_8
XFILLER_31_658 VPWR VGND sg13g2_decap_8
XFILLER_8_821 VPWR VGND sg13g2_decap_8
XFILLER_30_168 VPWR VGND sg13g2_decap_8
XFILLER_7_320 VPWR VGND sg13g2_decap_8
XFILLER_11_371 VPWR VGND sg13g2_decap_8
XFILLER_8_898 VPWR VGND sg13g2_decap_8
XFILLER_7_397 VPWR VGND sg13g2_decap_8
XFILLER_7_89 VPWR VGND sg13g2_decap_8
XFILLER_3_592 VPWR VGND sg13g2_decap_8
XFILLER_39_714 VPWR VGND sg13g2_decap_8
XFILLER_38_224 VPWR VGND sg13g2_decap_8
XFILLER_47_791 VPWR VGND sg13g2_decap_8
XFILLER_19_482 VPWR VGND sg13g2_decap_8
XFILLER_35_931 VPWR VGND sg13g2_decap_8
XFILLER_34_441 VPWR VGND sg13g2_decap_8
XFILLER_22_625 VPWR VGND sg13g2_decap_8
XFILLER_21_157 VPWR VGND sg13g2_decap_8
XFILLER_1_518 VPWR VGND sg13g2_decap_8
XFILLER_29_235 VPWR VGND sg13g2_decap_8
XFILLER_45_728 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_decap_8
XFILLER_26_942 VPWR VGND sg13g2_decap_8
XFILLER_38_791 VPWR VGND sg13g2_decap_8
XFILLER_25_452 VPWR VGND sg13g2_decap_8
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_16_65 VPWR VGND sg13g2_decap_8
XFILLER_41_945 VPWR VGND sg13g2_decap_8
XFILLER_13_636 VPWR VGND sg13g2_decap_8
XFILLER_9_629 VPWR VGND sg13g2_decap_8
XFILLER_40_455 VPWR VGND sg13g2_decap_8
XFILLER_32_42 VPWR VGND sg13g2_decap_8
XFILLER_5_857 VPWR VGND sg13g2_decap_8
XFILLER_4_323 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_588 VPWR VGND sg13g2_decap_8
XFILLER_36_728 VPWR VGND sg13g2_decap_8
XFILLER_17_920 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_decap_8
XFILLER_17_997 VPWR VGND sg13g2_decap_8
XFILLER_16_496 VPWR VGND sg13g2_decap_8
XFILLER_32_945 VPWR VGND sg13g2_decap_8
XFILLER_31_455 VPWR VGND sg13g2_decap_8
XFILLER_8_695 VPWR VGND sg13g2_decap_8
XFILLER_7_194 VPWR VGND sg13g2_decap_8
XFILLER_4_890 VPWR VGND sg13g2_decap_8
XFILLER_39_511 VPWR VGND sg13g2_decap_8
XFILLER_39_588 VPWR VGND sg13g2_decap_8
XFILLER_26_249 VPWR VGND sg13g2_decap_8
XFILLER_22_422 VPWR VGND sg13g2_decap_8
XFILLER_23_956 VPWR VGND sg13g2_decap_8
XFILLER_10_639 VPWR VGND sg13g2_decap_8
XFILLER_22_499 VPWR VGND sg13g2_decap_8
XFILLER_33_1022 VPWR VGND sg13g2_decap_8
XFILLER_2_805 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_18_717 VPWR VGND sg13g2_decap_8
XFILLER_40_1015 VPWR VGND sg13g2_decap_8
XFILLER_45_525 VPWR VGND sg13g2_decap_8
XFILLER_17_227 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_fill_2
XFILLER_27_86 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_decap_8
XFILLER_41_742 VPWR VGND sg13g2_decap_8
XFILLER_13_433 VPWR VGND sg13g2_decap_8
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_9_426 VPWR VGND sg13g2_decap_8
XFILLER_14_989 VPWR VGND sg13g2_decap_8
XFILLER_40_252 VPWR VGND sg13g2_decap_8
XFILLER_5_654 VPWR VGND sg13g2_decap_8
XFILLER_4_120 VPWR VGND sg13g2_decap_8
XFILLER_4_197 VPWR VGND sg13g2_decap_8
XFILLER_1_882 VPWR VGND sg13g2_decap_8
XFILLER_49_886 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_36_525 VPWR VGND sg13g2_decap_8
XFILLER_16_293 VPWR VGND sg13g2_decap_8
XFILLER_17_794 VPWR VGND sg13g2_decap_8
XFILLER_32_742 VPWR VGND sg13g2_decap_8
XFILLER_31_252 VPWR VGND sg13g2_decap_8
XFILLER_20_959 VPWR VGND sg13g2_decap_8
XFILLER_9_993 VPWR VGND sg13g2_decap_8
XFILLER_8_492 VPWR VGND sg13g2_decap_8
XFILLER_39_385 VPWR VGND sg13g2_decap_8
XFILLER_27_569 VPWR VGND sg13g2_decap_8
XFILLER_14_219 VPWR VGND sg13g2_decap_8
XFILLER_42_539 VPWR VGND sg13g2_decap_8
XFILLER_23_753 VPWR VGND sg13g2_decap_8
XFILLER_7_908 VPWR VGND sg13g2_decap_8
XFILLER_11_959 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
XFILLER_10_436 VPWR VGND sg13g2_decap_8
XFILLER_22_296 VPWR VGND sg13g2_decap_8
XFILLER_6_418 VPWR VGND sg13g2_decap_8
XFILLER_13_88 VPWR VGND sg13g2_fill_1
XFILLER_13_99 VPWR VGND sg13g2_decap_8
XFILLER_2_602 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_2_679 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
XFILLER_46_812 VPWR VGND sg13g2_decap_8
XFILLER_18_514 VPWR VGND sg13g2_decap_8
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_46_889 VPWR VGND sg13g2_decap_8
XFILLER_45_399 VPWR VGND sg13g2_decap_8
XFILLER_33_539 VPWR VGND sg13g2_decap_8
XFILLER_13_230 VPWR VGND sg13g2_decap_8
XFILLER_9_223 VPWR VGND sg13g2_decap_8
XFILLER_14_786 VPWR VGND sg13g2_decap_8
XFILLER_6_985 VPWR VGND sg13g2_decap_8
XFILLER_5_451 VPWR VGND sg13g2_decap_8
XFILLER_49_683 VPWR VGND sg13g2_decap_8
XFILLER_37_812 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_37_889 VPWR VGND sg13g2_decap_8
XFILLER_17_591 VPWR VGND sg13g2_decap_8
XFILLER_36_399 VPWR VGND sg13g2_decap_8
XFILLER_20_756 VPWR VGND sg13g2_decap_8
XFILLER_9_790 VPWR VGND sg13g2_decap_8
XFILLER_47_609 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_28_823 VPWR VGND sg13g2_decap_8
XFILLER_39_182 VPWR VGND sg13g2_decap_8
XFILLER_43_826 VPWR VGND sg13g2_decap_8
XFILLER_27_366 VPWR VGND sg13g2_decap_8
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_23_550 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_10_233 VPWR VGND sg13g2_decap_8
XFILLER_7_705 VPWR VGND sg13g2_decap_8
XFILLER_11_756 VPWR VGND sg13g2_decap_8
XFILLER_6_215 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_decap_8
XFILLER_3_900 VPWR VGND sg13g2_decap_8
XFILLER_3_977 VPWR VGND sg13g2_decap_8
XFILLER_2_476 VPWR VGND sg13g2_decap_8
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_38_609 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_18_311 VPWR VGND sg13g2_decap_8
XFILLER_19_867 VPWR VGND sg13g2_decap_8
XFILLER_46_686 VPWR VGND sg13g2_decap_8
XFILLER_34_826 VPWR VGND sg13g2_decap_8
XFILLER_45_196 VPWR VGND sg13g2_decap_8
XFILLER_18_388 VPWR VGND sg13g2_decap_8
XFILLER_33_336 VPWR VGND sg13g2_decap_8
XFILLER_14_583 VPWR VGND sg13g2_decap_8
XFILLER_6_782 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
XFILLER_49_480 VPWR VGND sg13g2_decap_8
X_79_ net4 net12 VPWR VGND sg13g2_buf_1
XFILLER_37_686 VPWR VGND sg13g2_decap_8
XFILLER_25_837 VPWR VGND sg13g2_decap_8
XFILLER_36_196 VPWR VGND sg13g2_decap_8
XFILLER_24_347 VPWR VGND sg13g2_decap_8
XFILLER_20_553 VPWR VGND sg13g2_decap_8
XFILLER_4_708 VPWR VGND sg13g2_decap_8
XFILLER_3_207 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_19_32 VPWR VGND sg13g2_decap_8
XFILLER_28_620 VPWR VGND sg13g2_decap_8
XFILLER_16_804 VPWR VGND sg13g2_decap_8
XFILLER_43_623 VPWR VGND sg13g2_decap_8
XFILLER_27_163 VPWR VGND sg13g2_decap_8
XFILLER_28_697 VPWR VGND sg13g2_decap_8
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_15_358 VPWR VGND sg13g2_decap_8
XFILLER_7_502 VPWR VGND sg13g2_decap_8
XFILLER_11_553 VPWR VGND sg13g2_decap_8
XFILLER_7_579 VPWR VGND sg13g2_decap_8
XFILLER_3_774 VPWR VGND sg13g2_decap_8
XFILLER_2_273 VPWR VGND sg13g2_decap_8
XFILLER_38_406 VPWR VGND sg13g2_decap_8
XFILLER_47_973 VPWR VGND sg13g2_decap_8
XFILLER_19_664 VPWR VGND sg13g2_decap_8
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_18_185 VPWR VGND sg13g2_decap_8
XFILLER_34_623 VPWR VGND sg13g2_decap_8
XFILLER_22_807 VPWR VGND sg13g2_decap_8
XFILLER_33_133 VPWR VGND sg13g2_decap_8
XFILLER_14_380 VPWR VGND sg13g2_decap_8
XFILLER_21_339 VPWR VGND sg13g2_decap_8
XFILLER_30_840 VPWR VGND sg13g2_decap_8
XFILLER_5_1018 VPWR VGND sg13g2_decap_8
XFILLER_29_417 VPWR VGND sg13g2_decap_8
XFILLER_38_973 VPWR VGND sg13g2_decap_8
XFILLER_25_634 VPWR VGND sg13g2_decap_8
XFILLER_37_483 VPWR VGND sg13g2_decap_8
XFILLER_24_144 VPWR VGND sg13g2_decap_8
XFILLER_12_317 VPWR VGND sg13g2_decap_8
XFILLER_13_818 VPWR VGND sg13g2_decap_8
XFILLER_40_637 VPWR VGND sg13g2_decap_8
XFILLER_20_350 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_4_505 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_29_984 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_44_910 VPWR VGND sg13g2_decap_8
XFILLER_16_601 VPWR VGND sg13g2_decap_8
XFILLER_28_494 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_44_987 VPWR VGND sg13g2_decap_8
XFILLER_15_155 VPWR VGND sg13g2_decap_8
XFILLER_16_678 VPWR VGND sg13g2_decap_8
XFILLER_43_497 VPWR VGND sg13g2_decap_8
XFILLER_31_637 VPWR VGND sg13g2_decap_8
XFILLER_8_800 VPWR VGND sg13g2_decap_8
XFILLER_11_350 VPWR VGND sg13g2_decap_8
XFILLER_30_147 VPWR VGND sg13g2_decap_8
XFILLER_12_884 VPWR VGND sg13g2_decap_8
XFILLER_8_877 VPWR VGND sg13g2_decap_8
XFILLER_7_68 VPWR VGND sg13g2_decap_8
XFILLER_7_376 VPWR VGND sg13g2_decap_8
XFILLER_3_571 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_19_461 VPWR VGND sg13g2_decap_8
XFILLER_35_910 VPWR VGND sg13g2_decap_8
XFILLER_46_280 VPWR VGND sg13g2_decap_8
XFILLER_34_420 VPWR VGND sg13g2_decap_8
XFILLER_22_604 VPWR VGND sg13g2_decap_8
XFILLER_35_987 VPWR VGND sg13g2_decap_8
XFILLER_21_136 VPWR VGND sg13g2_decap_8
XFILLER_34_497 VPWR VGND sg13g2_decap_8
X_59__24 VPWR VGND net23 sg13g2_tiehi
XFILLER_29_214 VPWR VGND sg13g2_decap_8
XFILLER_45_707 VPWR VGND sg13g2_decap_8
XFILLER_17_409 VPWR VGND sg13g2_decap_8
XFILLER_44_217 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_26_921 VPWR VGND sg13g2_decap_8
XFILLER_38_770 VPWR VGND sg13g2_decap_8
XFILLER_16_22 VPWR VGND sg13g2_fill_2
XFILLER_16_44 VPWR VGND sg13g2_decap_8
XFILLER_25_431 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_41_924 VPWR VGND sg13g2_decap_8
XFILLER_13_615 VPWR VGND sg13g2_decap_8
XFILLER_26_998 VPWR VGND sg13g2_decap_8
XFILLER_9_608 VPWR VGND sg13g2_decap_8
XFILLER_40_434 VPWR VGND sg13g2_decap_8
XFILLER_32_21 VPWR VGND sg13g2_decap_8
XFILLER_32_98 VPWR VGND sg13g2_decap_8
XFILLER_5_836 VPWR VGND sg13g2_decap_8
XFILLER_4_302 VPWR VGND sg13g2_decap_8
XFILLER_4_379 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_decap_8
XFILLER_36_707 VPWR VGND sg13g2_decap_8
XFILLER_29_781 VPWR VGND sg13g2_decap_8
XFILLER_35_217 VPWR VGND sg13g2_decap_8
XFILLER_28_291 VPWR VGND sg13g2_decap_8
XFILLER_44_784 VPWR VGND sg13g2_decap_8
XFILLER_16_475 VPWR VGND sg13g2_decap_8
XFILLER_17_976 VPWR VGND sg13g2_decap_8
XFILLER_32_924 VPWR VGND sg13g2_decap_8
XFILLER_43_294 VPWR VGND sg13g2_decap_8
XFILLER_31_434 VPWR VGND sg13g2_decap_8
XFILLER_12_681 VPWR VGND sg13g2_decap_8
XFILLER_8_674 VPWR VGND sg13g2_decap_8
XFILLER_7_173 VPWR VGND sg13g2_decap_8
XFILLER_39_567 VPWR VGND sg13g2_decap_8
XFILLER_26_228 VPWR VGND sg13g2_decap_8
XFILLER_22_401 VPWR VGND sg13g2_decap_8
XFILLER_35_784 VPWR VGND sg13g2_decap_8
XFILLER_23_935 VPWR VGND sg13g2_decap_8
XFILLER_34_294 VPWR VGND sg13g2_decap_8
XFILLER_10_618 VPWR VGND sg13g2_decap_8
XFILLER_33_1001 VPWR VGND sg13g2_decap_8
XFILLER_22_478 VPWR VGND sg13g2_decap_8
XFILLER_45_504 VPWR VGND sg13g2_decap_8
XFILLER_17_206 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_41_721 VPWR VGND sg13g2_decap_8
XFILLER_13_412 VPWR VGND sg13g2_decap_8
XFILLER_26_795 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_9_405 VPWR VGND sg13g2_decap_8
XFILLER_14_968 VPWR VGND sg13g2_decap_8
XFILLER_40_231 VPWR VGND sg13g2_decap_8
XFILLER_41_798 VPWR VGND sg13g2_decap_8
XFILLER_13_489 VPWR VGND sg13g2_decap_8
XFILLER_5_633 VPWR VGND sg13g2_decap_8
XFILLER_4_176 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_49_865 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_36_504 VPWR VGND sg13g2_decap_8
XFILLER_17_773 VPWR VGND sg13g2_decap_8
XFILLER_44_581 VPWR VGND sg13g2_decap_8
XFILLER_16_272 VPWR VGND sg13g2_decap_8
XFILLER_32_721 VPWR VGND sg13g2_decap_8
XFILLER_17_1018 VPWR VGND sg13g2_decap_8
XFILLER_31_231 VPWR VGND sg13g2_decap_8
XFILLER_20_938 VPWR VGND sg13g2_decap_8
XFILLER_32_798 VPWR VGND sg13g2_decap_8
XFILLER_9_972 VPWR VGND sg13g2_decap_8
XFILLER_8_471 VPWR VGND sg13g2_decap_8
XFILLER_39_364 VPWR VGND sg13g2_decap_8
XFILLER_27_548 VPWR VGND sg13g2_decap_8
XFILLER_42_518 VPWR VGND sg13g2_decap_8
XFILLER_23_732 VPWR VGND sg13g2_decap_8
XFILLER_35_581 VPWR VGND sg13g2_decap_8
XFILLER_10_415 VPWR VGND sg13g2_decap_8
XFILLER_11_938 VPWR VGND sg13g2_decap_8
XFILLER_22_275 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_2_658 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_46_868 VPWR VGND sg13g2_decap_8
XFILLER_45_378 VPWR VGND sg13g2_decap_8
XFILLER_33_518 VPWR VGND sg13g2_decap_8
XFILLER_26_592 VPWR VGND sg13g2_decap_8
XFILLER_14_765 VPWR VGND sg13g2_decap_8
XFILLER_9_202 VPWR VGND sg13g2_decap_8
XFILLER_41_595 VPWR VGND sg13g2_decap_8
XFILLER_13_286 VPWR VGND sg13g2_decap_8
XFILLER_9_279 VPWR VGND sg13g2_decap_8
XFILLER_10_982 VPWR VGND sg13g2_decap_8
XFILLER_6_964 VPWR VGND sg13g2_decap_8
XFILLER_5_430 VPWR VGND sg13g2_decap_8
XFILLER_49_662 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_37_868 VPWR VGND sg13g2_decap_8
XFILLER_36_378 VPWR VGND sg13g2_decap_8
XFILLER_17_570 VPWR VGND sg13g2_decap_8
XFILLER_24_529 VPWR VGND sg13g2_decap_8
XFILLER_20_735 VPWR VGND sg13g2_decap_8
XFILLER_32_595 VPWR VGND sg13g2_decap_8
XFILLER_30_1015 VPWR VGND sg13g2_decap_8
XFILLER_28_802 VPWR VGND sg13g2_decap_8
XFILLER_39_161 VPWR VGND sg13g2_decap_8
XFILLER_43_805 VPWR VGND sg13g2_decap_8
XFILLER_27_345 VPWR VGND sg13g2_decap_8
XFILLER_28_879 VPWR VGND sg13g2_decap_8
XFILLER_42_315 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_10_212 VPWR VGND sg13g2_decap_8
XFILLER_11_735 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_10_289 VPWR VGND sg13g2_decap_8
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_3_956 VPWR VGND sg13g2_decap_8
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_46_1022 VPWR VGND sg13g2_decap_8
XFILLER_2_455 VPWR VGND sg13g2_decap_8
XFILLER_49_74 VPWR VGND sg13g2_decap_8
XFILLER_19_846 VPWR VGND sg13g2_decap_8
XFILLER_46_665 VPWR VGND sg13g2_decap_8
XFILLER_18_367 VPWR VGND sg13g2_decap_8
XFILLER_34_805 VPWR VGND sg13g2_decap_8
XFILLER_45_175 VPWR VGND sg13g2_decap_8
XFILLER_33_315 VPWR VGND sg13g2_decap_8
XFILLER_42_882 VPWR VGND sg13g2_decap_8
XFILLER_14_562 VPWR VGND sg13g2_decap_8
XFILLER_41_392 VPWR VGND sg13g2_decap_8
XFILLER_6_761 VPWR VGND sg13g2_decap_8
XFILLER_28_109 VPWR VGND sg13g2_decap_8
X_78_ net3 net11 VPWR VGND sg13g2_buf_1
XFILLER_25_816 VPWR VGND sg13g2_decap_8
XFILLER_37_665 VPWR VGND sg13g2_decap_8
XFILLER_24_326 VPWR VGND sg13g2_decap_8
XFILLER_36_175 VPWR VGND sg13g2_decap_8
XFILLER_40_819 VPWR VGND sg13g2_decap_8
XFILLER_33_882 VPWR VGND sg13g2_decap_8
XFILLER_20_532 VPWR VGND sg13g2_decap_8
XFILLER_32_392 VPWR VGND sg13g2_decap_8
XFILLER_10_46 VPWR VGND sg13g2_decap_8
XFILLER_10_79 VPWR VGND sg13g2_decap_8
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_43_602 VPWR VGND sg13g2_decap_8
XFILLER_27_142 VPWR VGND sg13g2_decap_8
XFILLER_28_676 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_15_337 VPWR VGND sg13g2_decap_8
XFILLER_43_679 VPWR VGND sg13g2_decap_8
XFILLER_31_819 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_11_532 VPWR VGND sg13g2_decap_8
XFILLER_24_893 VPWR VGND sg13g2_decap_8
XFILLER_30_329 VPWR VGND sg13g2_decap_8
XFILLER_7_558 VPWR VGND sg13g2_decap_8
XFILLER_13_1021 VPWR VGND sg13g2_decap_8
XFILLER_3_753 VPWR VGND sg13g2_decap_8
XFILLER_2_252 VPWR VGND sg13g2_decap_8
XFILLER_47_952 VPWR VGND sg13g2_decap_8
XFILLER_19_643 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
XFILLER_18_164 VPWR VGND sg13g2_decap_8
XFILLER_34_602 VPWR VGND sg13g2_decap_8
XFILLER_33_112 VPWR VGND sg13g2_decap_8
XFILLER_21_318 VPWR VGND sg13g2_decap_8
XFILLER_34_679 VPWR VGND sg13g2_decap_8
XFILLER_33_189 VPWR VGND sg13g2_decap_8
XFILLER_30_896 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_8
XFILLER_38_952 VPWR VGND sg13g2_decap_8
XFILLER_25_613 VPWR VGND sg13g2_decap_8
XFILLER_37_462 VPWR VGND sg13g2_decap_8
XFILLER_24_123 VPWR VGND sg13g2_decap_8
XFILLER_40_616 VPWR VGND sg13g2_decap_8
XFILLER_21_885 VPWR VGND sg13g2_decap_8
XFILLER_21_67 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_48_749 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_29_963 VPWR VGND sg13g2_decap_8
XFILLER_28_473 VPWR VGND sg13g2_decap_8
XFILLER_44_966 VPWR VGND sg13g2_decap_8
XFILLER_15_134 VPWR VGND sg13g2_decap_8
XFILLER_16_657 VPWR VGND sg13g2_decap_8
XFILLER_43_476 VPWR VGND sg13g2_decap_8
XFILLER_31_616 VPWR VGND sg13g2_decap_8
XFILLER_24_690 VPWR VGND sg13g2_decap_8
XFILLER_30_126 VPWR VGND sg13g2_decap_8
XFILLER_12_863 VPWR VGND sg13g2_decap_8
XFILLER_8_856 VPWR VGND sg13g2_decap_8
XFILLER_7_25 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_7_355 VPWR VGND sg13g2_decap_8
XFILLER_7_47 VPWR VGND sg13g2_decap_8
XFILLER_3_550 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_39_749 VPWR VGND sg13g2_decap_8
XFILLER_19_440 VPWR VGND sg13g2_decap_8
XFILLER_38_259 VPWR VGND sg13g2_decap_8
XFILLER_35_966 VPWR VGND sg13g2_decap_8
XFILLER_34_476 VPWR VGND sg13g2_decap_8
XFILLER_21_115 VPWR VGND sg13g2_decap_8
XFILLER_30_693 VPWR VGND sg13g2_decap_8
XFILLER_26_900 VPWR VGND sg13g2_decap_8
XFILLER_25_410 VPWR VGND sg13g2_decap_8
XFILLER_41_903 VPWR VGND sg13g2_decap_8
XFILLER_26_977 VPWR VGND sg13g2_decap_8
XFILLER_25_487 VPWR VGND sg13g2_decap_8
XFILLER_40_413 VPWR VGND sg13g2_decap_8
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_21_682 VPWR VGND sg13g2_decap_8
XFILLER_5_815 VPWR VGND sg13g2_decap_8
XFILLER_32_77 VPWR VGND sg13g2_decap_8
XFILLER_10_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_358 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_29_760 VPWR VGND sg13g2_decap_8
XFILLER_17_955 VPWR VGND sg13g2_decap_8
XFILLER_28_270 VPWR VGND sg13g2_decap_8
XFILLER_44_763 VPWR VGND sg13g2_decap_8
XFILLER_16_454 VPWR VGND sg13g2_decap_8
XFILLER_32_903 VPWR VGND sg13g2_decap_8
XFILLER_43_273 VPWR VGND sg13g2_decap_8
XFILLER_31_413 VPWR VGND sg13g2_decap_8
XFILLER_12_660 VPWR VGND sg13g2_decap_8
XFILLER_40_980 VPWR VGND sg13g2_decap_8
XFILLER_8_653 VPWR VGND sg13g2_decap_8
XFILLER_7_152 VPWR VGND sg13g2_decap_8
XFILLER_39_546 VPWR VGND sg13g2_decap_8
XFILLER_26_207 VPWR VGND sg13g2_decap_8
XFILLER_23_914 VPWR VGND sg13g2_decap_8
XFILLER_35_763 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_decap_8
XFILLER_22_457 VPWR VGND sg13g2_decap_8
XFILLER_31_980 VPWR VGND sg13g2_decap_8
XFILLER_30_490 VPWR VGND sg13g2_decap_8
XFILLER_27_44 VPWR VGND sg13g2_fill_1
XFILLER_41_700 VPWR VGND sg13g2_decap_8
XFILLER_26_774 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_14_947 VPWR VGND sg13g2_decap_8
XFILLER_25_284 VPWR VGND sg13g2_decap_8
XFILLER_40_210 VPWR VGND sg13g2_decap_8
XFILLER_41_777 VPWR VGND sg13g2_decap_8
XFILLER_13_468 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_5_612 VPWR VGND sg13g2_decap_8
XFILLER_5_689 VPWR VGND sg13g2_decap_8
XFILLER_4_155 VPWR VGND sg13g2_decap_8
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_49_844 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
XFILLER_44_560 VPWR VGND sg13g2_decap_8
XFILLER_16_251 VPWR VGND sg13g2_decap_8
XFILLER_17_752 VPWR VGND sg13g2_decap_8
XFILLER_32_700 VPWR VGND sg13g2_decap_8
XFILLER_31_210 VPWR VGND sg13g2_decap_8
XFILLER_20_917 VPWR VGND sg13g2_decap_8
XFILLER_32_777 VPWR VGND sg13g2_decap_8
XFILLER_9_951 VPWR VGND sg13g2_decap_8
XFILLER_31_287 VPWR VGND sg13g2_decap_8
XFILLER_8_450 VPWR VGND sg13g2_decap_8
XFILLER_39_343 VPWR VGND sg13g2_decap_8
XFILLER_27_527 VPWR VGND sg13g2_decap_8
XFILLER_23_711 VPWR VGND sg13g2_decap_8
XFILLER_35_560 VPWR VGND sg13g2_decap_8
XFILLER_11_917 VPWR VGND sg13g2_decap_8
XFILLER_22_254 VPWR VGND sg13g2_decap_8
XFILLER_23_788 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_2_637 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_46_847 VPWR VGND sg13g2_decap_8
XFILLER_18_549 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_45_357 VPWR VGND sg13g2_decap_8
XFILLER_26_571 VPWR VGND sg13g2_decap_8
XFILLER_14_744 VPWR VGND sg13g2_decap_8
XFILLER_41_574 VPWR VGND sg13g2_decap_8
XFILLER_13_265 VPWR VGND sg13g2_decap_8
XFILLER_9_258 VPWR VGND sg13g2_decap_8
XFILLER_10_961 VPWR VGND sg13g2_decap_8
XFILLER_6_943 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_486 VPWR VGND sg13g2_decap_8
XFILLER_49_641 VPWR VGND sg13g2_decap_8
XFILLER_23_1012 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_37_847 VPWR VGND sg13g2_decap_8
XFILLER_24_508 VPWR VGND sg13g2_decap_8
XFILLER_36_357 VPWR VGND sg13g2_decap_8
XFILLER_20_714 VPWR VGND sg13g2_decap_8
XFILLER_32_574 VPWR VGND sg13g2_decap_8
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_1017 VPWR VGND sg13g2_decap_8
XFILLER_39_140 VPWR VGND sg13g2_decap_8
XFILLER_27_324 VPWR VGND sg13g2_decap_8
XFILLER_28_858 VPWR VGND sg13g2_decap_8
XFILLER_15_519 VPWR VGND sg13g2_decap_8
XFILLER_11_714 VPWR VGND sg13g2_decap_8
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_23_585 VPWR VGND sg13g2_decap_8
XFILLER_10_268 VPWR VGND sg13g2_decap_8
XFILLER_40_77 VPWR VGND sg13g2_decap_8
XFILLER_3_935 VPWR VGND sg13g2_decap_8
XFILLER_46_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_434 VPWR VGND sg13g2_decap_8
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_19_825 VPWR VGND sg13g2_decap_8
XFILLER_46_644 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_18_346 VPWR VGND sg13g2_decap_8
XFILLER_27_891 VPWR VGND sg13g2_decap_8
XFILLER_14_541 VPWR VGND sg13g2_decap_8
XFILLER_42_861 VPWR VGND sg13g2_decap_8
XFILLER_41_371 VPWR VGND sg13g2_decap_8
XFILLER_6_740 VPWR VGND sg13g2_decap_8
XFILLER_5_283 VPWR VGND sg13g2_decap_8
XFILLER_37_644 VPWR VGND sg13g2_decap_8
XFILLER_24_305 VPWR VGND sg13g2_decap_8
XFILLER_36_154 VPWR VGND sg13g2_decap_8
XFILLER_33_861 VPWR VGND sg13g2_decap_8
XFILLER_20_511 VPWR VGND sg13g2_decap_8
XFILLER_32_371 VPWR VGND sg13g2_decap_8
XFILLER_20_588 VPWR VGND sg13g2_decap_8
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_0_938 VPWR VGND sg13g2_decap_8
XFILLER_19_67 VPWR VGND sg13g2_decap_8
XFILLER_27_121 VPWR VGND sg13g2_decap_8
XFILLER_28_655 VPWR VGND sg13g2_decap_8
XFILLER_15_316 VPWR VGND sg13g2_decap_8
XFILLER_16_839 VPWR VGND sg13g2_decap_8
XFILLER_43_658 VPWR VGND sg13g2_decap_8
XFILLER_27_198 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_decap_8
XFILLER_24_872 VPWR VGND sg13g2_decap_8
XFILLER_30_308 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_11_511 VPWR VGND sg13g2_decap_8
XFILLER_23_382 VPWR VGND sg13g2_decap_8
XFILLER_13_1000 VPWR VGND sg13g2_decap_8
XFILLER_7_537 VPWR VGND sg13g2_decap_8
XFILLER_11_588 VPWR VGND sg13g2_decap_8
XFILLER_3_732 VPWR VGND sg13g2_decap_8
XFILLER_2_231 VPWR VGND sg13g2_decap_8
XFILLER_47_931 VPWR VGND sg13g2_decap_8
XFILLER_19_622 VPWR VGND sg13g2_decap_8
XFILLER_46_441 VPWR VGND sg13g2_decap_8
XFILLER_20_1015 VPWR VGND sg13g2_decap_8
XFILLER_19_699 VPWR VGND sg13g2_decap_8
XFILLER_34_658 VPWR VGND sg13g2_decap_8
XFILLER_33_168 VPWR VGND sg13g2_decap_8
XFILLER_15_883 VPWR VGND sg13g2_decap_8
XFILLER_30_875 VPWR VGND sg13g2_decap_8
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_38_931 VPWR VGND sg13g2_decap_8
XFILLER_37_441 VPWR VGND sg13g2_decap_8
XFILLER_24_102 VPWR VGND sg13g2_decap_8
XFILLER_25_669 VPWR VGND sg13g2_decap_8
XFILLER_24_179 VPWR VGND sg13g2_decap_8
XFILLER_36_1022 VPWR VGND sg13g2_decap_8
XFILLER_21_864 VPWR VGND sg13g2_decap_8
XFILLER_20_385 VPWR VGND sg13g2_decap_8
XFILLER_21_46 VPWR VGND sg13g2_decap_8
XFILLER_43_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_29_942 VPWR VGND sg13g2_decap_8
XFILLER_28_452 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_44_945 VPWR VGND sg13g2_decap_8
XFILLER_16_636 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_30_105 VPWR VGND sg13g2_decap_8
XFILLER_12_842 VPWR VGND sg13g2_decap_8
XFILLER_8_835 VPWR VGND sg13g2_decap_8
XFILLER_7_334 VPWR VGND sg13g2_decap_8
XFILLER_11_385 VPWR VGND sg13g2_decap_8
XFILLER_30_7 VPWR VGND sg13g2_decap_8
XFILLER_39_728 VPWR VGND sg13g2_decap_8
XFILLER_38_238 VPWR VGND sg13g2_decap_8
XFILLER_19_496 VPWR VGND sg13g2_decap_8
XFILLER_35_945 VPWR VGND sg13g2_decap_8
XFILLER_34_455 VPWR VGND sg13g2_decap_8
XFILLER_15_680 VPWR VGND sg13g2_decap_8
XFILLER_22_639 VPWR VGND sg13g2_decap_8
XFILLER_30_672 VPWR VGND sg13g2_decap_8
XFILLER_29_249 VPWR VGND sg13g2_decap_8
XFILLER_26_956 VPWR VGND sg13g2_decap_8
XFILLER_25_466 VPWR VGND sg13g2_decap_8
XFILLER_41_959 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_decap_8
XFILLER_16_79 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_4
XFILLER_12_149 VPWR VGND sg13g2_decap_8
XFILLER_40_469 VPWR VGND sg13g2_decap_8
XFILLER_21_661 VPWR VGND sg13g2_decap_8
XFILLER_32_56 VPWR VGND sg13g2_decap_8
XFILLER_20_182 VPWR VGND sg13g2_decap_8
XFILLER_10_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_337 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_44_742 VPWR VGND sg13g2_decap_8
XFILLER_16_433 VPWR VGND sg13g2_decap_8
XFILLER_17_934 VPWR VGND sg13g2_decap_8
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_32_959 VPWR VGND sg13g2_decap_8
XFILLER_31_469 VPWR VGND sg13g2_decap_8
XFILLER_8_632 VPWR VGND sg13g2_decap_8
XFILLER_7_131 VPWR VGND sg13g2_decap_8
XFILLER_11_182 VPWR VGND sg13g2_decap_8
XFILLER_39_525 VPWR VGND sg13g2_decap_8
XFILLER_27_709 VPWR VGND sg13g2_decap_8
XFILLER_19_293 VPWR VGND sg13g2_decap_8
XFILLER_35_742 VPWR VGND sg13g2_decap_8
XFILLER_34_252 VPWR VGND sg13g2_decap_8
XFILLER_22_436 VPWR VGND sg13g2_decap_8
XFILLER_2_819 VPWR VGND sg13g2_decap_8
XFILLER_1_329 VPWR VGND sg13g2_decap_8
XFILLER_45_539 VPWR VGND sg13g2_decap_8
XFILLER_26_753 VPWR VGND sg13g2_decap_8
XFILLER_14_926 VPWR VGND sg13g2_decap_8
XFILLER_25_263 VPWR VGND sg13g2_decap_8
XFILLER_41_756 VPWR VGND sg13g2_decap_8
XFILLER_13_447 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_5_668 VPWR VGND sg13g2_decap_8
XFILLER_4_134 VPWR VGND sg13g2_decap_8
XFILLER_49_823 VPWR VGND sg13g2_decap_8
XFILLER_1_896 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_731 VPWR VGND sg13g2_decap_8
XFILLER_36_539 VPWR VGND sg13g2_decap_8
XFILLER_16_230 VPWR VGND sg13g2_decap_8
XFILLER_32_756 VPWR VGND sg13g2_decap_8
XFILLER_9_930 VPWR VGND sg13g2_decap_8
XFILLER_31_266 VPWR VGND sg13g2_decap_8
XFILLER_39_322 VPWR VGND sg13g2_decap_8
XFILLER_27_506 VPWR VGND sg13g2_decap_8
XFILLER_39_399 VPWR VGND sg13g2_decap_8
XFILLER_22_233 VPWR VGND sg13g2_decap_8
XFILLER_23_767 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_2_616 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_46_826 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_45_336 VPWR VGND sg13g2_decap_8
XFILLER_18_528 VPWR VGND sg13g2_decap_8
XFILLER_26_550 VPWR VGND sg13g2_decap_8
XFILLER_14_723 VPWR VGND sg13g2_decap_8
XFILLER_41_553 VPWR VGND sg13g2_decap_8
XFILLER_13_244 VPWR VGND sg13g2_decap_8
XFILLER_9_237 VPWR VGND sg13g2_decap_8
XFILLER_6_922 VPWR VGND sg13g2_decap_8
XFILLER_10_940 VPWR VGND sg13g2_decap_8
XFILLER_5_465 VPWR VGND sg13g2_decap_8
XFILLER_6_999 VPWR VGND sg13g2_decap_8
XFILLER_49_620 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_37_826 VPWR VGND sg13g2_decap_8
XFILLER_49_697 VPWR VGND sg13g2_decap_8
XFILLER_36_336 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_32_553 VPWR VGND sg13g2_decap_8
XFILLER_5_70 VPWR VGND sg13g2_decap_8
XFILLER_27_303 VPWR VGND sg13g2_decap_8
XFILLER_28_837 VPWR VGND sg13g2_decap_8
XFILLER_39_196 VPWR VGND sg13g2_decap_8
XFILLER_23_564 VPWR VGND sg13g2_decap_8
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_10_247 VPWR VGND sg13g2_decap_8
XFILLER_7_719 VPWR VGND sg13g2_decap_8
XFILLER_6_229 VPWR VGND sg13g2_decap_8
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_3_914 VPWR VGND sg13g2_decap_8
XFILLER_2_413 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_19_804 VPWR VGND sg13g2_decap_8
XFILLER_46_623 VPWR VGND sg13g2_decap_8
XFILLER_18_325 VPWR VGND sg13g2_decap_8
XFILLER_45_133 VPWR VGND sg13g2_decap_8
XFILLER_27_870 VPWR VGND sg13g2_decap_8
XFILLER_42_840 VPWR VGND sg13g2_decap_8
XFILLER_14_520 VPWR VGND sg13g2_decap_8
XFILLER_41_350 VPWR VGND sg13g2_decap_8
XFILLER_14_597 VPWR VGND sg13g2_decap_8
XFILLER_14_90 VPWR VGND sg13g2_decap_4
XFILLER_6_796 VPWR VGND sg13g2_decap_8
XFILLER_5_262 VPWR VGND sg13g2_decap_8
XFILLER_2_980 VPWR VGND sg13g2_decap_8
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_49_494 VPWR VGND sg13g2_decap_8
XFILLER_37_623 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_18_892 VPWR VGND sg13g2_decap_8
XFILLER_33_840 VPWR VGND sg13g2_decap_8
XFILLER_32_350 VPWR VGND sg13g2_decap_8
XFILLER_20_567 VPWR VGND sg13g2_decap_8
XFILLER_10_15 VPWR VGND sg13g2_fill_2
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_27_100 VPWR VGND sg13g2_decap_8
XFILLER_28_634 VPWR VGND sg13g2_decap_8
XFILLER_16_818 VPWR VGND sg13g2_decap_8
XFILLER_27_177 VPWR VGND sg13g2_decap_8
XFILLER_43_637 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_24_851 VPWR VGND sg13g2_decap_8
XFILLER_23_361 VPWR VGND sg13g2_decap_8
XFILLER_11_567 VPWR VGND sg13g2_decap_8
XFILLER_7_516 VPWR VGND sg13g2_decap_8
XFILLER_3_711 VPWR VGND sg13g2_decap_8
XFILLER_2_210 VPWR VGND sg13g2_decap_8
XFILLER_3_788 VPWR VGND sg13g2_decap_8
XFILLER_2_287 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_decap_8
XFILLER_19_601 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_47_987 VPWR VGND sg13g2_decap_8
XFILLER_19_678 VPWR VGND sg13g2_decap_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
XFILLER_18_199 VPWR VGND sg13g2_decap_8
XFILLER_34_637 VPWR VGND sg13g2_decap_8
XFILLER_15_862 VPWR VGND sg13g2_decap_8
XFILLER_33_147 VPWR VGND sg13g2_decap_8
XFILLER_14_394 VPWR VGND sg13g2_decap_8
XFILLER_30_854 VPWR VGND sg13g2_decap_8
XFILLER_6_593 VPWR VGND sg13g2_decap_8
XFILLER_38_910 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
XFILLER_2_93 VPWR VGND sg13g2_fill_1
XFILLER_37_420 VPWR VGND sg13g2_decap_8
X_59_ net23 VGND VPWR _05_ net5 clknet_1_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_987 VPWR VGND sg13g2_decap_8
XFILLER_25_648 VPWR VGND sg13g2_decap_8
XFILLER_37_497 VPWR VGND sg13g2_decap_8
XFILLER_24_158 VPWR VGND sg13g2_decap_8
XFILLER_36_1001 VPWR VGND sg13g2_decap_8
XFILLER_21_843 VPWR VGND sg13g2_decap_8
XFILLER_20_364 VPWR VGND sg13g2_decap_8
XFILLER_21_25 VPWR VGND sg13g2_decap_8
XFILLER_4_519 VPWR VGND sg13g2_decap_8
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_29_921 VPWR VGND sg13g2_decap_8
XFILLER_28_431 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_44_924 VPWR VGND sg13g2_decap_8
XFILLER_16_615 VPWR VGND sg13g2_decap_8
XFILLER_29_998 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_15_169 VPWR VGND sg13g2_decap_8
XFILLER_12_821 VPWR VGND sg13g2_decap_8
XFILLER_8_814 VPWR VGND sg13g2_decap_8
XFILLER_7_313 VPWR VGND sg13g2_decap_8
XFILLER_11_364 VPWR VGND sg13g2_decap_8
XFILLER_12_898 VPWR VGND sg13g2_decap_8
XFILLER_3_585 VPWR VGND sg13g2_decap_8
XFILLER_39_707 VPWR VGND sg13g2_decap_8
XFILLER_38_217 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_19_475 VPWR VGND sg13g2_decap_8
XFILLER_35_924 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
XFILLER_34_434 VPWR VGND sg13g2_decap_8
XFILLER_22_618 VPWR VGND sg13g2_decap_8
XFILLER_14_191 VPWR VGND sg13g2_decap_8
XFILLER_30_651 VPWR VGND sg13g2_decap_8
XFILLER_7_880 VPWR VGND sg13g2_decap_8
XFILLER_6_390 VPWR VGND sg13g2_decap_8
XFILLER_29_228 VPWR VGND sg13g2_decap_8
XFILLER_38_784 VPWR VGND sg13g2_decap_8
XFILLER_26_935 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_decap_8
XFILLER_16_58 VPWR VGND sg13g2_decap_8
XFILLER_25_445 VPWR VGND sg13g2_decap_8
XFILLER_41_938 VPWR VGND sg13g2_decap_8
XFILLER_13_629 VPWR VGND sg13g2_decap_8
XFILLER_21_640 VPWR VGND sg13g2_decap_8
XFILLER_40_448 VPWR VGND sg13g2_decap_8
XFILLER_32_35 VPWR VGND sg13g2_decap_8
XFILLER_20_161 VPWR VGND sg13g2_decap_8
XFILLER_4_316 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_17_913 VPWR VGND sg13g2_decap_8
XFILLER_44_721 VPWR VGND sg13g2_decap_8
XFILLER_16_412 VPWR VGND sg13g2_decap_8
XFILLER_29_795 VPWR VGND sg13g2_decap_8
XFILLER_43_231 VPWR VGND sg13g2_decap_8
XFILLER_44_798 VPWR VGND sg13g2_decap_8
XFILLER_16_489 VPWR VGND sg13g2_decap_8
XFILLER_32_938 VPWR VGND sg13g2_decap_8
XFILLER_31_448 VPWR VGND sg13g2_decap_8
XFILLER_8_611 VPWR VGND sg13g2_decap_8
XFILLER_7_110 VPWR VGND sg13g2_decap_8
XFILLER_11_161 VPWR VGND sg13g2_decap_8
XFILLER_12_695 VPWR VGND sg13g2_decap_8
XFILLER_8_688 VPWR VGND sg13g2_decap_8
XFILLER_7_187 VPWR VGND sg13g2_decap_8
XFILLER_4_883 VPWR VGND sg13g2_decap_8
XFILLER_3_382 VPWR VGND sg13g2_decap_8
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_39_504 VPWR VGND sg13g2_decap_8
XFILLER_47_581 VPWR VGND sg13g2_decap_8
XFILLER_19_272 VPWR VGND sg13g2_decap_8
XFILLER_35_721 VPWR VGND sg13g2_decap_8
XFILLER_34_231 VPWR VGND sg13g2_decap_8
XFILLER_22_415 VPWR VGND sg13g2_decap_8
XFILLER_23_949 VPWR VGND sg13g2_decap_8
XFILLER_35_798 VPWR VGND sg13g2_decap_8
XFILLER_33_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_81 VPWR VGND sg13g2_decap_8
XFILLER_1_308 VPWR VGND sg13g2_decap_8
XFILLER_40_1008 VPWR VGND sg13g2_decap_8
XFILLER_45_518 VPWR VGND sg13g2_decap_8
XFILLER_27_35 VPWR VGND sg13g2_decap_8
XFILLER_26_732 VPWR VGND sg13g2_decap_8
XFILLER_38_581 VPWR VGND sg13g2_decap_8
XFILLER_14_905 VPWR VGND sg13g2_decap_8
XFILLER_25_242 VPWR VGND sg13g2_decap_8
XFILLER_27_79 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_41_735 VPWR VGND sg13g2_decap_8
XFILLER_13_426 VPWR VGND sg13g2_decap_8
XFILLER_9_419 VPWR VGND sg13g2_decap_8
XFILLER_40_245 VPWR VGND sg13g2_decap_8
XFILLER_22_982 VPWR VGND sg13g2_decap_8
XFILLER_5_647 VPWR VGND sg13g2_decap_8
XFILLER_4_113 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_fill_2
X_61__22 VPWR VGND net21 sg13g2_tiehi
XFILLER_49_802 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_1_875 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_49_879 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_36_518 VPWR VGND sg13g2_decap_8
XFILLER_17_710 VPWR VGND sg13g2_decap_8
XFILLER_29_592 VPWR VGND sg13g2_decap_8
XFILLER_17_787 VPWR VGND sg13g2_decap_8
XFILLER_44_595 VPWR VGND sg13g2_decap_8
XFILLER_16_286 VPWR VGND sg13g2_decap_8
XFILLER_32_735 VPWR VGND sg13g2_decap_8
XFILLER_31_245 VPWR VGND sg13g2_decap_8
XFILLER_13_993 VPWR VGND sg13g2_decap_8
XFILLER_9_986 VPWR VGND sg13g2_decap_8
XFILLER_12_492 VPWR VGND sg13g2_decap_8
XFILLER_8_485 VPWR VGND sg13g2_decap_8
XFILLER_4_680 VPWR VGND sg13g2_decap_8
XFILLER_39_301 VPWR VGND sg13g2_decap_8
XFILLER_39_378 VPWR VGND sg13g2_decap_8
XFILLER_22_212 VPWR VGND sg13g2_decap_8
XFILLER_23_746 VPWR VGND sg13g2_decap_8
XFILLER_35_595 VPWR VGND sg13g2_decap_8
XFILLER_10_429 VPWR VGND sg13g2_decap_8
XFILLER_22_289 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_46_805 VPWR VGND sg13g2_decap_8
XFILLER_18_507 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_14_702 VPWR VGND sg13g2_decap_8
XFILLER_41_532 VPWR VGND sg13g2_decap_8
XFILLER_13_223 VPWR VGND sg13g2_decap_8
XFILLER_9_216 VPWR VGND sg13g2_decap_8
XFILLER_14_779 VPWR VGND sg13g2_decap_8
XFILLER_16_1021 VPWR VGND sg13g2_decap_8
XFILLER_6_901 VPWR VGND sg13g2_decap_8
XFILLER_10_996 VPWR VGND sg13g2_decap_8
XFILLER_6_978 VPWR VGND sg13g2_decap_8
XFILLER_5_444 VPWR VGND sg13g2_decap_8
XFILLER_1_672 VPWR VGND sg13g2_decap_8
XFILLER_49_676 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_37_805 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_45_882 VPWR VGND sg13g2_decap_8
XFILLER_44_392 VPWR VGND sg13g2_decap_8
XFILLER_17_584 VPWR VGND sg13g2_decap_8
XFILLER_32_532 VPWR VGND sg13g2_decap_8
XFILLER_20_749 VPWR VGND sg13g2_decap_8
XFILLER_13_790 VPWR VGND sg13g2_decap_8
XFILLER_8_282 VPWR VGND sg13g2_decap_8
XFILLER_9_783 VPWR VGND sg13g2_decap_8
XFILLER_28_816 VPWR VGND sg13g2_decap_8
XFILLER_39_175 VPWR VGND sg13g2_decap_8
XFILLER_27_359 VPWR VGND sg13g2_decap_8
XFILLER_43_819 VPWR VGND sg13g2_decap_8
XFILLER_36_882 VPWR VGND sg13g2_decap_8
XFILLER_42_329 VPWR VGND sg13g2_decap_8
XFILLER_35_392 VPWR VGND sg13g2_decap_8
XFILLER_23_543 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_11_749 VPWR VGND sg13g2_decap_8
XFILLER_10_226 VPWR VGND sg13g2_decap_8
XFILLER_6_208 VPWR VGND sg13g2_decap_8
XFILLER_40_35 VPWR VGND sg13g2_decap_8
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_2_469 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_46_602 VPWR VGND sg13g2_decap_8
XFILLER_18_304 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_46_679 VPWR VGND sg13g2_decap_8
XFILLER_34_819 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
XFILLER_33_329 VPWR VGND sg13g2_decap_8
XFILLER_42_896 VPWR VGND sg13g2_decap_8
XFILLER_14_576 VPWR VGND sg13g2_decap_8
XFILLER_10_793 VPWR VGND sg13g2_decap_8
XFILLER_6_775 VPWR VGND sg13g2_decap_8
XFILLER_5_241 VPWR VGND sg13g2_decap_8
XFILLER_49_473 VPWR VGND sg13g2_decap_8
XFILLER_37_602 VPWR VGND sg13g2_decap_8
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_18_871 VPWR VGND sg13g2_decap_8
XFILLER_37_679 VPWR VGND sg13g2_decap_8
XFILLER_17_381 VPWR VGND sg13g2_decap_8
XFILLER_36_189 VPWR VGND sg13g2_decap_8
XFILLER_33_896 VPWR VGND sg13g2_decap_8
XFILLER_20_546 VPWR VGND sg13g2_decap_8
XFILLER_9_580 VPWR VGND sg13g2_decap_8
XFILLER_19_25 VPWR VGND sg13g2_decap_8
XFILLER_28_613 VPWR VGND sg13g2_decap_8
XFILLER_43_616 VPWR VGND sg13g2_decap_8
XFILLER_27_156 VPWR VGND sg13g2_decap_8
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_24_830 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
XFILLER_23_340 VPWR VGND sg13g2_decap_8
XFILLER_11_546 VPWR VGND sg13g2_decap_8
XFILLER_3_767 VPWR VGND sg13g2_decap_8
XFILLER_2_266 VPWR VGND sg13g2_decap_8
XFILLER_47_966 VPWR VGND sg13g2_decap_8
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_19_657 VPWR VGND sg13g2_decap_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_34_616 VPWR VGND sg13g2_decap_8
XFILLER_18_178 VPWR VGND sg13g2_decap_8
XFILLER_33_126 VPWR VGND sg13g2_decap_8
XFILLER_15_841 VPWR VGND sg13g2_decap_8
XFILLER_14_373 VPWR VGND sg13g2_decap_8
XFILLER_42_693 VPWR VGND sg13g2_decap_8
XFILLER_30_833 VPWR VGND sg13g2_decap_8
XFILLER_10_590 VPWR VGND sg13g2_decap_8
XFILLER_6_572 VPWR VGND sg13g2_decap_8
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_2_72 VPWR VGND sg13g2_decap_8
XFILLER_38_966 VPWR VGND sg13g2_decap_8
X_58_ net VGND VPWR _04_ net4 clknet_1_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_37_476 VPWR VGND sg13g2_decap_8
XFILLER_25_627 VPWR VGND sg13g2_decap_8
XFILLER_24_137 VPWR VGND sg13g2_decap_8
XFILLER_21_822 VPWR VGND sg13g2_decap_8
XFILLER_33_693 VPWR VGND sg13g2_decap_8
XFILLER_20_343 VPWR VGND sg13g2_decap_8
XFILLER_21_899 VPWR VGND sg13g2_decap_8
XFILLER_29_900 VPWR VGND sg13g2_decap_8
XFILLER_28_410 VPWR VGND sg13g2_decap_8
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_44_903 VPWR VGND sg13g2_decap_8
XFILLER_29_977 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_28_487 VPWR VGND sg13g2_decap_8
XFILLER_15_148 VPWR VGND sg13g2_decap_8
XFILLER_12_800 VPWR VGND sg13g2_decap_8
XFILLER_11_343 VPWR VGND sg13g2_decap_8
XFILLER_12_877 VPWR VGND sg13g2_decap_8
XFILLER_7_39 VPWR VGND sg13g2_decap_4
XFILLER_7_369 VPWR VGND sg13g2_decap_8
XFILLER_3_564 VPWR VGND sg13g2_decap_8
XFILLER_11_81 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_19_454 VPWR VGND sg13g2_decap_8
XFILLER_35_903 VPWR VGND sg13g2_decap_8
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_34_413 VPWR VGND sg13g2_decap_8
XFILLER_43_980 VPWR VGND sg13g2_decap_8
XFILLER_42_490 VPWR VGND sg13g2_decap_8
XFILLER_14_170 VPWR VGND sg13g2_decap_8
XFILLER_21_129 VPWR VGND sg13g2_decap_8
XFILLER_30_630 VPWR VGND sg13g2_decap_8
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_29_207 VPWR VGND sg13g2_decap_8
XFILLER_26_914 VPWR VGND sg13g2_decap_8
XFILLER_38_763 VPWR VGND sg13g2_decap_8
XFILLER_25_424 VPWR VGND sg13g2_decap_8
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_41_917 VPWR VGND sg13g2_decap_8
XFILLER_13_608 VPWR VGND sg13g2_decap_8
XFILLER_16_37 VPWR VGND sg13g2_decap_8
XFILLER_34_980 VPWR VGND sg13g2_decap_8
XFILLER_40_427 VPWR VGND sg13g2_decap_8
XFILLER_33_490 VPWR VGND sg13g2_decap_8
XFILLER_20_140 VPWR VGND sg13g2_decap_8
XFILLER_32_14 VPWR VGND sg13g2_decap_8
XFILLER_21_696 VPWR VGND sg13g2_decap_8
XFILLER_5_829 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_44_700 VPWR VGND sg13g2_decap_8
XFILLER_29_774 VPWR VGND sg13g2_decap_8
XFILLER_43_210 VPWR VGND sg13g2_decap_8
XFILLER_28_284 VPWR VGND sg13g2_decap_8
XFILLER_17_969 VPWR VGND sg13g2_decap_8
XFILLER_44_777 VPWR VGND sg13g2_decap_8
XFILLER_16_468 VPWR VGND sg13g2_decap_8
XFILLER_32_917 VPWR VGND sg13g2_decap_8
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_25_991 VPWR VGND sg13g2_decap_8
XFILLER_31_427 VPWR VGND sg13g2_decap_8
XFILLER_11_140 VPWR VGND sg13g2_decap_8
XFILLER_12_674 VPWR VGND sg13g2_decap_8
XFILLER_40_994 VPWR VGND sg13g2_decap_8
XFILLER_8_667 VPWR VGND sg13g2_decap_8
XFILLER_7_166 VPWR VGND sg13g2_decap_8
XFILLER_4_862 VPWR VGND sg13g2_decap_8
XFILLER_3_361 VPWR VGND sg13g2_decap_8
XFILLER_26_1012 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_19_251 VPWR VGND sg13g2_decap_8
XFILLER_35_700 VPWR VGND sg13g2_decap_8
XFILLER_34_210 VPWR VGND sg13g2_decap_8
XFILLER_23_928 VPWR VGND sg13g2_decap_8
XFILLER_35_777 VPWR VGND sg13g2_decap_8
XFILLER_34_287 VPWR VGND sg13g2_decap_8
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_31_994 VPWR VGND sg13g2_decap_8
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_26_711 VPWR VGND sg13g2_decap_8
XFILLER_38_560 VPWR VGND sg13g2_decap_8
XFILLER_25_221 VPWR VGND sg13g2_decap_8
XFILLER_41_714 VPWR VGND sg13g2_decap_8
XFILLER_13_405 VPWR VGND sg13g2_decap_8
XFILLER_26_788 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_25_298 VPWR VGND sg13g2_decap_8
XFILLER_40_224 VPWR VGND sg13g2_decap_8
XFILLER_22_961 VPWR VGND sg13g2_decap_8
XFILLER_21_493 VPWR VGND sg13g2_decap_8
XFILLER_5_626 VPWR VGND sg13g2_decap_8
XFILLER_49_1012 VPWR VGND sg13g2_decap_8
XFILLER_4_169 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_fill_2
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_49_858 VPWR VGND sg13g2_decap_8
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_29_571 VPWR VGND sg13g2_decap_8
XFILLER_44_574 VPWR VGND sg13g2_decap_8
XFILLER_16_265 VPWR VGND sg13g2_decap_8
XFILLER_17_91 VPWR VGND sg13g2_decap_8
XFILLER_17_766 VPWR VGND sg13g2_decap_8
XFILLER_32_714 VPWR VGND sg13g2_decap_8
XFILLER_31_224 VPWR VGND sg13g2_decap_8
XFILLER_13_972 VPWR VGND sg13g2_decap_8
XFILLER_12_471 VPWR VGND sg13g2_decap_8
XFILLER_40_791 VPWR VGND sg13g2_decap_8
XFILLER_8_464 VPWR VGND sg13g2_decap_8
XFILLER_9_965 VPWR VGND sg13g2_decap_8
XFILLER_39_357 VPWR VGND sg13g2_decap_8
XFILLER_35_574 VPWR VGND sg13g2_decap_8
XFILLER_23_725 VPWR VGND sg13g2_decap_8
XFILLER_10_408 VPWR VGND sg13g2_decap_8
XFILLER_22_268 VPWR VGND sg13g2_decap_8
XFILLER_31_791 VPWR VGND sg13g2_decap_8
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_41_511 VPWR VGND sg13g2_decap_8
XFILLER_13_202 VPWR VGND sg13g2_decap_8
XFILLER_26_585 VPWR VGND sg13g2_decap_8
XFILLER_14_758 VPWR VGND sg13g2_decap_8
XFILLER_16_1000 VPWR VGND sg13g2_decap_8
XFILLER_41_588 VPWR VGND sg13g2_decap_8
XFILLER_13_279 VPWR VGND sg13g2_decap_8
XFILLER_21_290 VPWR VGND sg13g2_decap_8
XFILLER_10_975 VPWR VGND sg13g2_decap_8
XFILLER_6_957 VPWR VGND sg13g2_decap_8
XFILLER_5_423 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_49_655 VPWR VGND sg13g2_decap_8
XFILLER_23_1026 VPWR VGND sg13g2_fill_2
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_45_861 VPWR VGND sg13g2_decap_8
XFILLER_17_563 VPWR VGND sg13g2_decap_8
XFILLER_44_371 VPWR VGND sg13g2_decap_8
XFILLER_32_511 VPWR VGND sg13g2_decap_8
XFILLER_20_728 VPWR VGND sg13g2_decap_8
XFILLER_32_588 VPWR VGND sg13g2_decap_8
XFILLER_9_762 VPWR VGND sg13g2_decap_8
XFILLER_30_1008 VPWR VGND sg13g2_decap_8
XFILLER_8_261 VPWR VGND sg13g2_decap_8
XFILLER_5_990 VPWR VGND sg13g2_decap_8
XFILLER_5_94 VPWR VGND sg13g2_decap_8
XFILLER_39_154 VPWR VGND sg13g2_decap_8
XFILLER_27_338 VPWR VGND sg13g2_decap_8
XFILLER_42_308 VPWR VGND sg13g2_decap_8
XFILLER_36_861 VPWR VGND sg13g2_decap_8
XFILLER_23_522 VPWR VGND sg13g2_decap_8
XFILLER_35_371 VPWR VGND sg13g2_decap_8
XFILLER_39_1022 VPWR VGND sg13g2_decap_8
XFILLER_10_205 VPWR VGND sg13g2_decap_8
XFILLER_11_728 VPWR VGND sg13g2_decap_8
XFILLER_23_599 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_46_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_949 VPWR VGND sg13g2_decap_8
XFILLER_2_448 VPWR VGND sg13g2_decap_8
XFILLER_49_67 VPWR VGND sg13g2_decap_8
XFILLER_19_839 VPWR VGND sg13g2_decap_8
XFILLER_46_658 VPWR VGND sg13g2_decap_8
XFILLER_45_168 VPWR VGND sg13g2_decap_8
XFILLER_33_308 VPWR VGND sg13g2_decap_8
XFILLER_26_382 VPWR VGND sg13g2_decap_8
XFILLER_42_875 VPWR VGND sg13g2_decap_8
XFILLER_14_555 VPWR VGND sg13g2_decap_8
XFILLER_41_385 VPWR VGND sg13g2_decap_8
XFILLER_10_772 VPWR VGND sg13g2_decap_8
XFILLER_6_754 VPWR VGND sg13g2_decap_8
XFILLER_5_220 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_5_297 VPWR VGND sg13g2_decap_8
XFILLER_30_91 VPWR VGND sg13g2_decap_8
XFILLER_7_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_452 VPWR VGND sg13g2_decap_8
XFILLER_37_658 VPWR VGND sg13g2_decap_8
XFILLER_18_850 VPWR VGND sg13g2_decap_8
XFILLER_25_809 VPWR VGND sg13g2_decap_8
XFILLER_36_168 VPWR VGND sg13g2_decap_8
XFILLER_17_360 VPWR VGND sg13g2_decap_8
XFILLER_24_319 VPWR VGND sg13g2_decap_8
XFILLER_33_875 VPWR VGND sg13g2_decap_8
XFILLER_20_525 VPWR VGND sg13g2_decap_8
XFILLER_32_385 VPWR VGND sg13g2_decap_8
XFILLER_10_39 VPWR VGND sg13g2_decap_8
XFILLER_27_135 VPWR VGND sg13g2_decap_8
XFILLER_28_669 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_decap_8
XFILLER_24_886 VPWR VGND sg13g2_decap_8
XFILLER_11_525 VPWR VGND sg13g2_decap_8
XFILLER_23_396 VPWR VGND sg13g2_decap_8
XFILLER_13_1014 VPWR VGND sg13g2_decap_8
XFILLER_3_746 VPWR VGND sg13g2_decap_8
XFILLER_2_245 VPWR VGND sg13g2_decap_8
XFILLER_47_945 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_decap_8
XFILLER_19_636 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_18_157 VPWR VGND sg13g2_decap_8
XFILLER_15_820 VPWR VGND sg13g2_decap_8
XFILLER_33_105 VPWR VGND sg13g2_decap_8
XFILLER_42_672 VPWR VGND sg13g2_decap_8
XFILLER_14_352 VPWR VGND sg13g2_decap_8
XFILLER_15_897 VPWR VGND sg13g2_decap_8
XFILLER_30_812 VPWR VGND sg13g2_decap_8
XFILLER_41_182 VPWR VGND sg13g2_decap_8
XFILLER_30_889 VPWR VGND sg13g2_decap_8
XFILLER_6_551 VPWR VGND sg13g2_decap_8
XFILLER_38_945 VPWR VGND sg13g2_decap_8
XFILLER_25_606 VPWR VGND sg13g2_decap_8
X_57_ net20 VGND VPWR _03_ net3 clknet_1_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_37_455 VPWR VGND sg13g2_decap_8
XFILLER_24_116 VPWR VGND sg13g2_decap_8
XFILLER_40_609 VPWR VGND sg13g2_decap_8
XFILLER_21_801 VPWR VGND sg13g2_decap_8
XFILLER_33_672 VPWR VGND sg13g2_decap_8
XFILLER_20_322 VPWR VGND sg13g2_decap_8
XFILLER_32_182 VPWR VGND sg13g2_decap_8
XFILLER_21_878 VPWR VGND sg13g2_decap_8
XFILLER_20_399 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_29_956 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_28_466 VPWR VGND sg13g2_decap_8
XFILLER_44_959 VPWR VGND sg13g2_decap_8
XFILLER_15_127 VPWR VGND sg13g2_decap_8
XFILLER_31_609 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_30_119 VPWR VGND sg13g2_decap_8
XFILLER_11_322 VPWR VGND sg13g2_decap_8
XFILLER_12_856 VPWR VGND sg13g2_decap_8
XFILLER_24_683 VPWR VGND sg13g2_decap_8
XFILLER_23_193 VPWR VGND sg13g2_decap_8
XFILLER_8_849 VPWR VGND sg13g2_decap_8
XFILLER_7_348 VPWR VGND sg13g2_decap_8
XFILLER_11_399 VPWR VGND sg13g2_decap_8
XFILLER_11_60 VPWR VGND sg13g2_decap_8
XFILLER_3_543 VPWR VGND sg13g2_decap_8
XFILLER_4_1023 VPWR VGND sg13g2_decap_4
XFILLER_19_433 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_35_959 VPWR VGND sg13g2_decap_8
XFILLER_21_108 VPWR VGND sg13g2_decap_8
XFILLER_34_469 VPWR VGND sg13g2_decap_8
XFILLER_15_694 VPWR VGND sg13g2_decap_8
XFILLER_30_686 VPWR VGND sg13g2_decap_8
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_38_742 VPWR VGND sg13g2_decap_8
XFILLER_25_403 VPWR VGND sg13g2_decap_8
XFILLER_37_252 VPWR VGND sg13g2_decap_8
XFILLER_40_406 VPWR VGND sg13g2_decap_8
XFILLER_21_675 VPWR VGND sg13g2_decap_8
XFILLER_5_808 VPWR VGND sg13g2_decap_8
XFILLER_20_196 VPWR VGND sg13g2_decap_8
XFILLER_10_1017 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_29_753 VPWR VGND sg13g2_decap_8
XFILLER_17_948 VPWR VGND sg13g2_decap_8
XFILLER_28_263 VPWR VGND sg13g2_decap_8
XFILLER_44_756 VPWR VGND sg13g2_decap_8
XFILLER_16_447 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_decap_8
XFILLER_25_970 VPWR VGND sg13g2_decap_8
XFILLER_31_406 VPWR VGND sg13g2_decap_8
XFILLER_24_480 VPWR VGND sg13g2_decap_8
XFILLER_12_653 VPWR VGND sg13g2_decap_8
XFILLER_40_973 VPWR VGND sg13g2_decap_8
XFILLER_8_646 VPWR VGND sg13g2_decap_8
XFILLER_7_145 VPWR VGND sg13g2_decap_8
XFILLER_11_196 VPWR VGND sg13g2_decap_8
XFILLER_4_841 VPWR VGND sg13g2_decap_8
XFILLER_3_340 VPWR VGND sg13g2_decap_8
XFILLER_39_539 VPWR VGND sg13g2_decap_8
XFILLER_19_230 VPWR VGND sg13g2_decap_8
XFILLER_23_907 VPWR VGND sg13g2_decap_8
XFILLER_35_756 VPWR VGND sg13g2_decap_8
XFILLER_34_266 VPWR VGND sg13g2_decap_8
XFILLER_15_491 VPWR VGND sg13g2_decap_8
XFILLER_31_973 VPWR VGND sg13g2_decap_8
XFILLER_30_483 VPWR VGND sg13g2_decap_8
XFILLER_25_200 VPWR VGND sg13g2_decap_8
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_26_767 VPWR VGND sg13g2_decap_8
XFILLER_25_277 VPWR VGND sg13g2_decap_8
XFILLER_40_203 VPWR VGND sg13g2_decap_8
XFILLER_22_940 VPWR VGND sg13g2_decap_8
XFILLER_21_472 VPWR VGND sg13g2_decap_8
XFILLER_5_605 VPWR VGND sg13g2_decap_8
XFILLER_4_148 VPWR VGND sg13g2_decap_8
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_49_837 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_550 VPWR VGND sg13g2_decap_8
XFILLER_17_745 VPWR VGND sg13g2_decap_8
XFILLER_44_553 VPWR VGND sg13g2_decap_8
XFILLER_16_244 VPWR VGND sg13g2_decap_8
XFILLER_17_70 VPWR VGND sg13g2_decap_8
XFILLER_31_203 VPWR VGND sg13g2_decap_8
XFILLER_13_951 VPWR VGND sg13g2_decap_8
XFILLER_9_944 VPWR VGND sg13g2_decap_8
XFILLER_12_450 VPWR VGND sg13g2_decap_8
XFILLER_40_770 VPWR VGND sg13g2_decap_8
XFILLER_8_443 VPWR VGND sg13g2_decap_8
XFILLER_33_91 VPWR VGND sg13g2_decap_8
XFILLER_39_336 VPWR VGND sg13g2_decap_8
XFILLER_23_704 VPWR VGND sg13g2_decap_8
XFILLER_35_553 VPWR VGND sg13g2_decap_8
XFILLER_22_247 VPWR VGND sg13g2_decap_8
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_31_770 VPWR VGND sg13g2_decap_8
XFILLER_30_280 VPWR VGND sg13g2_decap_8
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_26_564 VPWR VGND sg13g2_decap_8
XFILLER_14_737 VPWR VGND sg13g2_decap_8
XFILLER_41_567 VPWR VGND sg13g2_decap_8
XFILLER_13_258 VPWR VGND sg13g2_decap_8
XFILLER_10_954 VPWR VGND sg13g2_decap_8
XFILLER_6_936 VPWR VGND sg13g2_decap_8
XFILLER_5_402 VPWR VGND sg13g2_decap_8
XFILLER_5_479 VPWR VGND sg13g2_decap_8
XFILLER_1_630 VPWR VGND sg13g2_decap_8
XFILLER_49_634 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_23_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_45_840 VPWR VGND sg13g2_decap_8
XFILLER_44_350 VPWR VGND sg13g2_decap_8
XFILLER_17_542 VPWR VGND sg13g2_decap_8
XFILLER_20_707 VPWR VGND sg13g2_decap_8
XFILLER_32_567 VPWR VGND sg13g2_decap_8
XFILLER_9_741 VPWR VGND sg13g2_decap_8
XFILLER_8_240 VPWR VGND sg13g2_decap_8
XFILLER_5_84 VPWR VGND sg13g2_decap_4
XFILLER_39_133 VPWR VGND sg13g2_decap_8
XFILLER_27_317 VPWR VGND sg13g2_decap_8
XFILLER_36_840 VPWR VGND sg13g2_decap_8
XFILLER_35_350 VPWR VGND sg13g2_decap_8
XFILLER_39_1001 VPWR VGND sg13g2_decap_8
XFILLER_23_501 VPWR VGND sg13g2_decap_8
XFILLER_11_707 VPWR VGND sg13g2_decap_8
XFILLER_23_578 VPWR VGND sg13g2_decap_8
XFILLER_3_928 VPWR VGND sg13g2_decap_8
XFILLER_2_427 VPWR VGND sg13g2_decap_8
XFILLER_49_46 VPWR VGND sg13g2_decap_8
XFILLER_19_818 VPWR VGND sg13g2_decap_8
XFILLER_46_637 VPWR VGND sg13g2_decap_8
XFILLER_18_339 VPWR VGND sg13g2_decap_8
XFILLER_45_147 VPWR VGND sg13g2_decap_8
XFILLER_26_361 VPWR VGND sg13g2_decap_8
XFILLER_27_884 VPWR VGND sg13g2_decap_8
XFILLER_42_854 VPWR VGND sg13g2_decap_8
XFILLER_14_534 VPWR VGND sg13g2_decap_8
XFILLER_41_364 VPWR VGND sg13g2_decap_8
XFILLER_14_71 VPWR VGND sg13g2_decap_8
XFILLER_10_751 VPWR VGND sg13g2_decap_8
XFILLER_6_733 VPWR VGND sg13g2_decap_8
XFILLER_5_276 VPWR VGND sg13g2_decap_8
XFILLER_30_70 VPWR VGND sg13g2_decap_8
XFILLER_2_994 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_431 VPWR VGND sg13g2_decap_8
XFILLER_37_637 VPWR VGND sg13g2_decap_8
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_33_854 VPWR VGND sg13g2_decap_8
XFILLER_20_504 VPWR VGND sg13g2_decap_8
XFILLER_32_364 VPWR VGND sg13g2_decap_8
XFILLER_27_114 VPWR VGND sg13g2_decap_8
XFILLER_28_648 VPWR VGND sg13g2_decap_8
XFILLER_15_309 VPWR VGND sg13g2_decap_8
XFILLER_24_865 VPWR VGND sg13g2_decap_8
XFILLER_11_504 VPWR VGND sg13g2_decap_8
XFILLER_23_375 VPWR VGND sg13g2_decap_8
XFILLER_3_725 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_2_224 VPWR VGND sg13g2_decap_8
XFILLER_47_924 VPWR VGND sg13g2_decap_8
XFILLER_19_615 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_20_1008 VPWR VGND sg13g2_decap_8
XFILLER_27_681 VPWR VGND sg13g2_decap_8
XFILLER_14_331 VPWR VGND sg13g2_decap_8
XFILLER_42_651 VPWR VGND sg13g2_decap_8
XFILLER_15_876 VPWR VGND sg13g2_decap_8
XFILLER_25_81 VPWR VGND sg13g2_decap_8
XFILLER_41_161 VPWR VGND sg13g2_decap_8
XFILLER_30_868 VPWR VGND sg13g2_decap_8
XFILLER_6_530 VPWR VGND sg13g2_decap_8
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_2_791 VPWR VGND sg13g2_decap_8
XFILLER_38_924 VPWR VGND sg13g2_decap_8
XFILLER_37_434 VPWR VGND sg13g2_decap_8
X_56_ net22 VGND VPWR net37 net10 clknet_1_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_651 VPWR VGND sg13g2_decap_8
XFILLER_36_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_301 VPWR VGND sg13g2_decap_8
XFILLER_32_161 VPWR VGND sg13g2_decap_8
XFILLER_21_857 VPWR VGND sg13g2_decap_8
XFILLER_20_378 VPWR VGND sg13g2_decap_8
XFILLER_21_39 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_43_1008 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_29_935 VPWR VGND sg13g2_decap_8
XFILLER_28_445 VPWR VGND sg13g2_decap_8
XFILLER_44_938 VPWR VGND sg13g2_decap_8
XFILLER_16_629 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_24_662 VPWR VGND sg13g2_decap_8
XFILLER_11_301 VPWR VGND sg13g2_decap_8
XFILLER_12_835 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_decap_8
XFILLER_8_828 VPWR VGND sg13g2_decap_8
XFILLER_7_327 VPWR VGND sg13g2_decap_8
XFILLER_11_378 VPWR VGND sg13g2_decap_8
XFILLER_3_522 VPWR VGND sg13g2_decap_8
XFILLER_3_599 VPWR VGND sg13g2_decap_8
XFILLER_47_721 VPWR VGND sg13g2_decap_8
XFILLER_4_1002 VPWR VGND sg13g2_decap_8
XFILLER_19_412 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_19_489 VPWR VGND sg13g2_decap_8
XFILLER_35_938 VPWR VGND sg13g2_decap_8
XFILLER_34_448 VPWR VGND sg13g2_decap_8
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_15_673 VPWR VGND sg13g2_decap_8
XFILLER_30_665 VPWR VGND sg13g2_decap_8
XFILLER_7_894 VPWR VGND sg13g2_decap_8
Xclkbuf_1_0__f_clk clknet_1_0__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_38_721 VPWR VGND sg13g2_decap_8
XFILLER_37_231 VPWR VGND sg13g2_decap_8
X_39_ net38 net8 _10_ _11_ _15_ VPWR VGND sg13g2_and4_1
XFILLER_38_798 VPWR VGND sg13g2_decap_8
XFILLER_26_949 VPWR VGND sg13g2_decap_8
XFILLER_12_109 VPWR VGND sg13g2_decap_8
XFILLER_25_459 VPWR VGND sg13g2_decap_8
XFILLER_21_654 VPWR VGND sg13g2_decap_8
XFILLER_20_175 VPWR VGND sg13g2_decap_8
XFILLER_32_49 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_29_732 VPWR VGND sg13g2_decap_8
XFILLER_17_927 VPWR VGND sg13g2_decap_8
XFILLER_28_242 VPWR VGND sg13g2_decap_8
XFILLER_44_735 VPWR VGND sg13g2_decap_8
XFILLER_16_426 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_12_632 VPWR VGND sg13g2_decap_8
XFILLER_40_952 VPWR VGND sg13g2_decap_8
XFILLER_8_625 VPWR VGND sg13g2_decap_8
XFILLER_7_124 VPWR VGND sg13g2_decap_8
XFILLER_11_175 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
XFILLER_4_820 VPWR VGND sg13g2_decap_8
XFILLER_22_71 VPWR VGND sg13g2_fill_2
XFILLER_4_897 VPWR VGND sg13g2_decap_8
XFILLER_3_396 VPWR VGND sg13g2_decap_8
XFILLER_39_518 VPWR VGND sg13g2_decap_8
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_19_286 VPWR VGND sg13g2_decap_8
XFILLER_35_735 VPWR VGND sg13g2_decap_8
XFILLER_34_245 VPWR VGND sg13g2_decap_8
XFILLER_15_470 VPWR VGND sg13g2_decap_8
XFILLER_16_993 VPWR VGND sg13g2_decap_8
XFILLER_22_429 VPWR VGND sg13g2_decap_8
XFILLER_31_952 VPWR VGND sg13g2_decap_8
XFILLER_30_462 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_7_691 VPWR VGND sg13g2_decap_8
XFILLER_26_746 VPWR VGND sg13g2_decap_8
XFILLER_38_595 VPWR VGND sg13g2_decap_8
XFILLER_14_919 VPWR VGND sg13g2_decap_8
XFILLER_25_256 VPWR VGND sg13g2_decap_8
XFILLER_41_749 VPWR VGND sg13g2_decap_8
XFILLER_40_259 VPWR VGND sg13g2_decap_8
XFILLER_21_451 VPWR VGND sg13g2_decap_8
XFILLER_22_996 VPWR VGND sg13g2_decap_8
XFILLER_4_127 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_49_816 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_44_532 VPWR VGND sg13g2_decap_8
XFILLER_16_223 VPWR VGND sg13g2_decap_8
XFILLER_17_724 VPWR VGND sg13g2_decap_8
XFILLER_32_749 VPWR VGND sg13g2_decap_8
XFILLER_13_930 VPWR VGND sg13g2_decap_8
XFILLER_31_259 VPWR VGND sg13g2_decap_8
XFILLER_8_422 VPWR VGND sg13g2_decap_8
XFILLER_9_923 VPWR VGND sg13g2_decap_8
XFILLER_33_70 VPWR VGND sg13g2_decap_8
XFILLER_8_499 VPWR VGND sg13g2_decap_8
XFILLER_4_694 VPWR VGND sg13g2_decap_8
XFILLER_3_193 VPWR VGND sg13g2_decap_8
XFILLER_39_315 VPWR VGND sg13g2_decap_8
XFILLER_48_882 VPWR VGND sg13g2_decap_8
XFILLER_47_392 VPWR VGND sg13g2_decap_8
XFILLER_35_532 VPWR VGND sg13g2_decap_8
XFILLER_16_790 VPWR VGND sg13g2_decap_8
XFILLER_22_226 VPWR VGND sg13g2_decap_8
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_2_609 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_46_819 VPWR VGND sg13g2_decap_8
XFILLER_45_329 VPWR VGND sg13g2_decap_8
XFILLER_39_882 VPWR VGND sg13g2_decap_8
XFILLER_26_543 VPWR VGND sg13g2_decap_8
XFILLER_38_392 VPWR VGND sg13g2_decap_8
XFILLER_14_716 VPWR VGND sg13g2_decap_8
XFILLER_41_546 VPWR VGND sg13g2_decap_8
XFILLER_13_237 VPWR VGND sg13g2_decap_8
XFILLER_10_933 VPWR VGND sg13g2_decap_8
XFILLER_22_793 VPWR VGND sg13g2_decap_8
XFILLER_6_915 VPWR VGND sg13g2_decap_8
XFILLER_5_458 VPWR VGND sg13g2_decap_8
XFILLER_49_613 VPWR VGND sg13g2_decap_8
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_819 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_17_521 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_36_329 VPWR VGND sg13g2_decap_8
XFILLER_45_896 VPWR VGND sg13g2_decap_8
XFILLER_17_598 VPWR VGND sg13g2_decap_8
XFILLER_32_546 VPWR VGND sg13g2_decap_8
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_9_720 VPWR VGND sg13g2_decap_8
XFILLER_8_296 VPWR VGND sg13g2_decap_8
XFILLER_9_797 VPWR VGND sg13g2_decap_8
XFILLER_5_63 VPWR VGND sg13g2_decap_8
XFILLER_4_491 VPWR VGND sg13g2_decap_8
XFILLER_39_112 VPWR VGND sg13g2_decap_8
XFILLER_39_189 VPWR VGND sg13g2_decap_8
XFILLER_36_896 VPWR VGND sg13g2_decap_8
XFILLER_23_557 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_3_907 VPWR VGND sg13g2_decap_8
XFILLER_2_406 VPWR VGND sg13g2_decap_8
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_46_616 VPWR VGND sg13g2_decap_8
XFILLER_45_126 VPWR VGND sg13g2_decap_8
XFILLER_18_318 VPWR VGND sg13g2_decap_8
XFILLER_26_340 VPWR VGND sg13g2_decap_8
XFILLER_27_863 VPWR VGND sg13g2_decap_8
XFILLER_14_513 VPWR VGND sg13g2_decap_8
XFILLER_42_833 VPWR VGND sg13g2_decap_8
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_10_730 VPWR VGND sg13g2_decap_8
XFILLER_14_50 VPWR VGND sg13g2_decap_8
XFILLER_6_712 VPWR VGND sg13g2_decap_8
XFILLER_22_590 VPWR VGND sg13g2_decap_8
XFILLER_5_255 VPWR VGND sg13g2_decap_8
XFILLER_6_789 VPWR VGND sg13g2_decap_8
XFILLER_2_973 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_37_616 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XFILLER_18_885 VPWR VGND sg13g2_decap_8
XFILLER_45_693 VPWR VGND sg13g2_decap_8
XFILLER_17_395 VPWR VGND sg13g2_decap_8
XFILLER_33_833 VPWR VGND sg13g2_decap_8
XFILLER_32_343 VPWR VGND sg13g2_decap_8
XFILLER_9_594 VPWR VGND sg13g2_decap_8
XFILLER_19_39 VPWR VGND sg13g2_decap_8
XFILLER_28_627 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_decap_8
XFILLER_24_844 VPWR VGND sg13g2_decap_8
XFILLER_36_693 VPWR VGND sg13g2_decap_8
XFILLER_23_354 VPWR VGND sg13g2_decap_8
XFILLER_7_509 VPWR VGND sg13g2_decap_8
XFILLER_3_704 VPWR VGND sg13g2_decap_8
XFILLER_2_203 VPWR VGND sg13g2_decap_8
XFILLER_47_903 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_27_660 VPWR VGND sg13g2_decap_8
XFILLER_42_630 VPWR VGND sg13g2_decap_8
XFILLER_14_310 VPWR VGND sg13g2_decap_8
XFILLER_15_855 VPWR VGND sg13g2_decap_8
XFILLER_25_60 VPWR VGND sg13g2_decap_8
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_14_387 VPWR VGND sg13g2_decap_8
XFILLER_30_847 VPWR VGND sg13g2_decap_8
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_6_586 VPWR VGND sg13g2_decap_8
XFILLER_29_1012 VPWR VGND sg13g2_decap_8
XFILLER_2_770 VPWR VGND sg13g2_decap_8
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_2_20 VPWR VGND sg13g2_fill_1
XFILLER_38_903 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_2_86 VPWR VGND sg13g2_decap_8
XFILLER_37_413 VPWR VGND sg13g2_decap_8
X_55_ net24 VGND VPWR net40 net9 clknet_1_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_46_980 VPWR VGND sg13g2_decap_8
XFILLER_45_490 VPWR VGND sg13g2_decap_8
XFILLER_18_682 VPWR VGND sg13g2_decap_8
XFILLER_33_630 VPWR VGND sg13g2_decap_8
XFILLER_17_192 VPWR VGND sg13g2_decap_8
XFILLER_32_140 VPWR VGND sg13g2_decap_8
XFILLER_21_836 VPWR VGND sg13g2_decap_8
XFILLER_20_357 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_9_391 VPWR VGND sg13g2_decap_8
XFILLER_0_707 VPWR VGND sg13g2_decap_8
XFILLER_29_914 VPWR VGND sg13g2_decap_8
XFILLER_28_424 VPWR VGND sg13g2_decap_8
XFILLER_44_917 VPWR VGND sg13g2_decap_8
XFILLER_16_608 VPWR VGND sg13g2_decap_8
XFILLER_37_980 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
XFILLER_36_490 VPWR VGND sg13g2_decap_8
XFILLER_24_641 VPWR VGND sg13g2_decap_8
XFILLER_12_814 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_8_807 VPWR VGND sg13g2_decap_8
XFILLER_7_306 VPWR VGND sg13g2_decap_8
XFILLER_11_357 VPWR VGND sg13g2_decap_8
XFILLER_3_501 VPWR VGND sg13g2_decap_8
XFILLER_3_578 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_decap_4
XFILLER_47_700 VPWR VGND sg13g2_decap_8
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_19_468 VPWR VGND sg13g2_decap_8
XFILLER_35_917 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
XFILLER_28_991 VPWR VGND sg13g2_decap_8
XFILLER_34_427 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_15_652 VPWR VGND sg13g2_decap_8
XFILLER_43_994 VPWR VGND sg13g2_decap_8
XFILLER_14_184 VPWR VGND sg13g2_decap_8
XFILLER_30_644 VPWR VGND sg13g2_decap_8
XFILLER_7_873 VPWR VGND sg13g2_decap_8
XFILLER_6_383 VPWR VGND sg13g2_decap_8
XFILLER_38_700 VPWR VGND sg13g2_decap_8
XFILLER_37_210 VPWR VGND sg13g2_decap_8
X_38_ VGND VPWR net8 _12_ _14_ net38 sg13g2_a21oi_1
XFILLER_26_928 VPWR VGND sg13g2_decap_8
XFILLER_38_777 VPWR VGND sg13g2_decap_8
XFILLER_16_18 VPWR VGND sg13g2_decap_4
XFILLER_25_438 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_decap_8
XFILLER_34_994 VPWR VGND sg13g2_decap_8
XFILLER_21_633 VPWR VGND sg13g2_decap_8
XFILLER_32_28 VPWR VGND sg13g2_decap_8
XFILLER_20_154 VPWR VGND sg13g2_decap_8
XFILLER_4_309 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_711 VPWR VGND sg13g2_decap_8
XFILLER_28_221 VPWR VGND sg13g2_decap_8
XFILLER_44_714 VPWR VGND sg13g2_decap_8
XFILLER_16_405 VPWR VGND sg13g2_decap_8
XFILLER_17_906 VPWR VGND sg13g2_decap_8
XFILLER_29_788 VPWR VGND sg13g2_decap_8
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_28_298 VPWR VGND sg13g2_decap_8
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_12_611 VPWR VGND sg13g2_decap_8
XFILLER_40_931 VPWR VGND sg13g2_decap_8
XFILLER_8_604 VPWR VGND sg13g2_decap_8
XFILLER_7_103 VPWR VGND sg13g2_decap_8
XFILLER_11_154 VPWR VGND sg13g2_decap_8
XFILLER_12_688 VPWR VGND sg13g2_decap_8
XFILLER_4_876 VPWR VGND sg13g2_decap_8
XFILLER_3_375 VPWR VGND sg13g2_decap_8
XFILLER_26_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_574 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
XFILLER_19_265 VPWR VGND sg13g2_decap_8
XFILLER_35_714 VPWR VGND sg13g2_decap_8
XFILLER_34_224 VPWR VGND sg13g2_decap_8
XFILLER_22_408 VPWR VGND sg13g2_decap_8
XFILLER_16_972 VPWR VGND sg13g2_decap_8
XFILLER_43_791 VPWR VGND sg13g2_decap_8
XFILLER_31_931 VPWR VGND sg13g2_decap_8
XFILLER_33_1008 VPWR VGND sg13g2_decap_8
XFILLER_30_441 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_decap_8
XFILLER_7_670 VPWR VGND sg13g2_decap_8
XFILLER_6_180 VPWR VGND sg13g2_decap_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_38_574 VPWR VGND sg13g2_decap_8
XFILLER_26_725 VPWR VGND sg13g2_decap_8
XFILLER_25_235 VPWR VGND sg13g2_decap_8
XFILLER_41_728 VPWR VGND sg13g2_decap_8
XFILLER_13_419 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
XFILLER_21_430 VPWR VGND sg13g2_decap_8
XFILLER_34_791 VPWR VGND sg13g2_decap_8
XFILLER_40_238 VPWR VGND sg13g2_decap_8
XFILLER_22_975 VPWR VGND sg13g2_decap_8
XFILLER_49_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_868 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_17_703 VPWR VGND sg13g2_decap_8
XFILLER_44_511 VPWR VGND sg13g2_decap_8
XFILLER_16_202 VPWR VGND sg13g2_decap_8
XFILLER_29_585 VPWR VGND sg13g2_decap_8
XFILLER_44_588 VPWR VGND sg13g2_decap_8
XFILLER_16_279 VPWR VGND sg13g2_decap_8
XFILLER_32_728 VPWR VGND sg13g2_decap_8
XFILLER_9_902 VPWR VGND sg13g2_decap_8
XFILLER_31_238 VPWR VGND sg13g2_decap_8
XFILLER_8_401 VPWR VGND sg13g2_decap_8
XFILLER_13_986 VPWR VGND sg13g2_decap_8
XFILLER_9_979 VPWR VGND sg13g2_decap_8
XFILLER_12_485 VPWR VGND sg13g2_decap_8
XFILLER_8_478 VPWR VGND sg13g2_decap_8
XFILLER_4_673 VPWR VGND sg13g2_decap_8
XFILLER_3_172 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_8
XFILLER_48_861 VPWR VGND sg13g2_decap_8
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_35_511 VPWR VGND sg13g2_decap_8
XFILLER_22_205 VPWR VGND sg13g2_decap_8
XFILLER_23_739 VPWR VGND sg13g2_decap_8
XFILLER_35_588 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_39_861 VPWR VGND sg13g2_decap_8
XFILLER_26_522 VPWR VGND sg13g2_decap_8
XFILLER_38_371 VPWR VGND sg13g2_decap_8
XFILLER_41_525 VPWR VGND sg13g2_decap_8
XFILLER_13_216 VPWR VGND sg13g2_decap_8
XFILLER_26_599 VPWR VGND sg13g2_decap_8
XFILLER_9_209 VPWR VGND sg13g2_decap_8
XFILLER_10_912 VPWR VGND sg13g2_decap_8
XFILLER_16_1014 VPWR VGND sg13g2_decap_8
XFILLER_22_772 VPWR VGND sg13g2_decap_8
XFILLER_5_437 VPWR VGND sg13g2_decap_8
XFILLER_10_989 VPWR VGND sg13g2_decap_8
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_49_669 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_17_500 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_29_382 VPWR VGND sg13g2_decap_8
XFILLER_45_875 VPWR VGND sg13g2_decap_8
XFILLER_17_577 VPWR VGND sg13g2_decap_8
XFILLER_44_385 VPWR VGND sg13g2_decap_8
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_32_525 VPWR VGND sg13g2_decap_8
XFILLER_13_783 VPWR VGND sg13g2_decap_8
XFILLER_9_776 VPWR VGND sg13g2_decap_8
XFILLER_12_282 VPWR VGND sg13g2_decap_8
XFILLER_8_275 VPWR VGND sg13g2_decap_8
XFILLER_5_20 VPWR VGND sg13g2_fill_1
XFILLER_5_42 VPWR VGND sg13g2_decap_8
XFILLER_4_470 VPWR VGND sg13g2_decap_8
XFILLER_28_809 VPWR VGND sg13g2_decap_8
XFILLER_39_168 VPWR VGND sg13g2_decap_8
XFILLER_36_875 VPWR VGND sg13g2_decap_8
XFILLER_23_536 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_35_385 VPWR VGND sg13g2_decap_8
XFILLER_10_219 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_27_842 VPWR VGND sg13g2_decap_8
XFILLER_42_812 VPWR VGND sg13g2_decap_8
XFILLER_26_396 VPWR VGND sg13g2_decap_8
XFILLER_41_322 VPWR VGND sg13g2_decap_8
XFILLER_42_889 VPWR VGND sg13g2_decap_8
XFILLER_14_569 VPWR VGND sg13g2_decap_8
XFILLER_41_399 VPWR VGND sg13g2_decap_8
XFILLER_10_786 VPWR VGND sg13g2_decap_8
XFILLER_6_768 VPWR VGND sg13g2_decap_8
XFILLER_5_234 VPWR VGND sg13g2_decap_8
XFILLER_2_952 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_39_70 VPWR VGND sg13g2_decap_8
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_45_672 VPWR VGND sg13g2_decap_8
XFILLER_18_864 VPWR VGND sg13g2_decap_8
XFILLER_33_812 VPWR VGND sg13g2_decap_8
XFILLER_44_182 VPWR VGND sg13g2_decap_8
XFILLER_17_374 VPWR VGND sg13g2_decap_8
XFILLER_32_322 VPWR VGND sg13g2_decap_8
XFILLER_33_889 VPWR VGND sg13g2_decap_8
XFILLER_13_580 VPWR VGND sg13g2_decap_8
XFILLER_20_539 VPWR VGND sg13g2_decap_8
XFILLER_32_399 VPWR VGND sg13g2_decap_8
XFILLER_9_573 VPWR VGND sg13g2_decap_8
XFILLER_19_18 VPWR VGND sg13g2_decap_8
XFILLER_28_606 VPWR VGND sg13g2_decap_8
XFILLER_27_149 VPWR VGND sg13g2_decap_8
XFILLER_43_609 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_36_672 VPWR VGND sg13g2_decap_8
XFILLER_42_119 VPWR VGND sg13g2_decap_8
XFILLER_24_823 VPWR VGND sg13g2_decap_8
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_23_333 VPWR VGND sg13g2_decap_8
XFILLER_11_539 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_259 VPWR VGND sg13g2_decap_8
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_47_959 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_34_609 VPWR VGND sg13g2_decap_8
XFILLER_15_834 VPWR VGND sg13g2_decap_8
XFILLER_33_119 VPWR VGND sg13g2_decap_8
XFILLER_26_193 VPWR VGND sg13g2_decap_8
XFILLER_42_686 VPWR VGND sg13g2_decap_8
XFILLER_14_366 VPWR VGND sg13g2_decap_8
XFILLER_30_826 VPWR VGND sg13g2_decap_8
XFILLER_41_196 VPWR VGND sg13g2_decap_8
XFILLER_10_583 VPWR VGND sg13g2_decap_8
XFILLER_6_565 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_2_65 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
X_54_ net25 VGND VPWR _00_ net8 clknet_1_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_959 VPWR VGND sg13g2_decap_8
XFILLER_18_661 VPWR VGND sg13g2_decap_8
XFILLER_37_469 VPWR VGND sg13g2_decap_8
XFILLER_17_171 VPWR VGND sg13g2_decap_8
XFILLER_21_815 VPWR VGND sg13g2_decap_8
XFILLER_33_686 VPWR VGND sg13g2_decap_8
XFILLER_20_336 VPWR VGND sg13g2_decap_8
XFILLER_32_196 VPWR VGND sg13g2_decap_8
XFILLER_9_370 VPWR VGND sg13g2_decap_8
XFILLER_28_403 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
XFILLER_24_620 VPWR VGND sg13g2_decap_8
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_24_697 VPWR VGND sg13g2_decap_8
XFILLER_11_336 VPWR VGND sg13g2_decap_8
XFILLER_11_74 VPWR VGND sg13g2_decap_8
XFILLER_3_557 VPWR VGND sg13g2_decap_8
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_19_447 VPWR VGND sg13g2_decap_8
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_28_970 VPWR VGND sg13g2_decap_8
XFILLER_34_406 VPWR VGND sg13g2_decap_8
XFILLER_43_973 VPWR VGND sg13g2_decap_8
XFILLER_15_631 VPWR VGND sg13g2_decap_8
XFILLER_14_163 VPWR VGND sg13g2_decap_8
XFILLER_30_623 VPWR VGND sg13g2_decap_8
XFILLER_42_483 VPWR VGND sg13g2_decap_8
XFILLER_10_380 VPWR VGND sg13g2_decap_8
XFILLER_7_852 VPWR VGND sg13g2_decap_8
XFILLER_6_362 VPWR VGND sg13g2_decap_8
XFILLER_38_756 VPWR VGND sg13g2_decap_8
X_37_ VGND VPWR net46 _12_ _00_ _13_ sg13g2_a21oi_1
XFILLER_26_907 VPWR VGND sg13g2_decap_8
XFILLER_37_266 VPWR VGND sg13g2_decap_8
XFILLER_25_417 VPWR VGND sg13g2_decap_8
XFILLER_21_612 VPWR VGND sg13g2_decap_8
XFILLER_34_973 VPWR VGND sg13g2_decap_8
XFILLER_33_483 VPWR VGND sg13g2_decap_8
XFILLER_20_133 VPWR VGND sg13g2_decap_8
XFILLER_21_689 VPWR VGND sg13g2_decap_8
XFILLER_28_200 VPWR VGND sg13g2_decap_8
XFILLER_29_767 VPWR VGND sg13g2_decap_8
XFILLER_43_203 VPWR VGND sg13g2_decap_8
XFILLER_28_277 VPWR VGND sg13g2_decap_8
XFILLER_25_984 VPWR VGND sg13g2_decap_8
XFILLER_40_910 VPWR VGND sg13g2_decap_8
XFILLER_24_494 VPWR VGND sg13g2_decap_8
XFILLER_11_133 VPWR VGND sg13g2_decap_8
XFILLER_12_667 VPWR VGND sg13g2_decap_8
XFILLER_40_987 VPWR VGND sg13g2_decap_8
XFILLER_7_159 VPWR VGND sg13g2_decap_8
XFILLER_4_855 VPWR VGND sg13g2_decap_8
XFILLER_3_354 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_26_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_19_244 VPWR VGND sg13g2_decap_8
XFILLER_34_203 VPWR VGND sg13g2_decap_8
XFILLER_16_951 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_decap_8
XFILLER_31_910 VPWR VGND sg13g2_decap_8
XFILLER_42_280 VPWR VGND sg13g2_decap_8
XFILLER_30_420 VPWR VGND sg13g2_decap_8
XFILLER_31_987 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_30_497 VPWR VGND sg13g2_decap_8
XFILLER_33_0 VPWR VGND sg13g2_decap_8
XFILLER_26_704 VPWR VGND sg13g2_decap_8
XFILLER_38_553 VPWR VGND sg13g2_decap_8
XFILLER_25_214 VPWR VGND sg13g2_decap_8
XFILLER_41_707 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_34_770 VPWR VGND sg13g2_decap_8
XFILLER_40_217 VPWR VGND sg13g2_decap_8
XFILLER_22_954 VPWR VGND sg13g2_decap_8
XFILLER_33_280 VPWR VGND sg13g2_decap_8
XFILLER_21_486 VPWR VGND sg13g2_decap_8
XFILLER_5_619 VPWR VGND sg13g2_decap_8
XFILLER_49_1005 VPWR VGND sg13g2_decap_8
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_29_564 VPWR VGND sg13g2_decap_8
XFILLER_17_759 VPWR VGND sg13g2_decap_8
XFILLER_32_707 VPWR VGND sg13g2_decap_8
XFILLER_44_567 VPWR VGND sg13g2_decap_8
XFILLER_16_258 VPWR VGND sg13g2_decap_8
XFILLER_17_84 VPWR VGND sg13g2_decap_8
XFILLER_31_217 VPWR VGND sg13g2_decap_8
XFILLER_25_781 VPWR VGND sg13g2_decap_8
XFILLER_12_464 VPWR VGND sg13g2_decap_8
XFILLER_13_965 VPWR VGND sg13g2_decap_8
XFILLER_24_291 VPWR VGND sg13g2_decap_8
XFILLER_9_958 VPWR VGND sg13g2_decap_8
XFILLER_40_784 VPWR VGND sg13g2_decap_8
XFILLER_8_457 VPWR VGND sg13g2_decap_8
XFILLER_4_652 VPWR VGND sg13g2_decap_8
XFILLER_3_151 VPWR VGND sg13g2_decap_8
XFILLER_48_840 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
XFILLER_23_718 VPWR VGND sg13g2_decap_8
XFILLER_35_567 VPWR VGND sg13g2_decap_8
XFILLER_31_784 VPWR VGND sg13g2_decap_8
XFILLER_30_294 VPWR VGND sg13g2_decap_8
XFILLER_38_28 VPWR VGND sg13g2_decap_8
XFILLER_39_840 VPWR VGND sg13g2_decap_8
XFILLER_26_501 VPWR VGND sg13g2_decap_8
XFILLER_38_350 VPWR VGND sg13g2_decap_8
XFILLER_41_504 VPWR VGND sg13g2_decap_8
XFILLER_26_578 VPWR VGND sg13g2_decap_8
XFILLER_22_751 VPWR VGND sg13g2_decap_8
XFILLER_10_968 VPWR VGND sg13g2_decap_8
XFILLER_21_283 VPWR VGND sg13g2_decap_8
XFILLER_5_416 VPWR VGND sg13g2_decap_8
XFILLER_1_644 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_49_648 VPWR VGND sg13g2_decap_8
XFILLER_23_1019 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_29_361 VPWR VGND sg13g2_decap_8
XFILLER_45_854 VPWR VGND sg13g2_decap_8
XFILLER_17_556 VPWR VGND sg13g2_decap_8
XFILLER_44_364 VPWR VGND sg13g2_decap_8
XFILLER_32_504 VPWR VGND sg13g2_decap_8
XFILLER_13_762 VPWR VGND sg13g2_decap_8
XFILLER_12_261 VPWR VGND sg13g2_decap_8
XFILLER_40_581 VPWR VGND sg13g2_decap_8
XFILLER_8_254 VPWR VGND sg13g2_decap_8
XFILLER_9_755 VPWR VGND sg13g2_decap_8
XFILLER_5_983 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_fill_1
XFILLER_39_147 VPWR VGND sg13g2_decap_8
XFILLER_36_854 VPWR VGND sg13g2_decap_8
XFILLER_23_515 VPWR VGND sg13g2_decap_8
XFILLER_35_364 VPWR VGND sg13g2_decap_8
XFILLER_39_1015 VPWR VGND sg13g2_decap_8
XFILLER_31_581 VPWR VGND sg13g2_decap_8
XFILLER_46_1008 VPWR VGND sg13g2_decap_8
XFILLER_27_821 VPWR VGND sg13g2_decap_8
XFILLER_14_548 VPWR VGND sg13g2_decap_8
XFILLER_26_375 VPWR VGND sg13g2_decap_8
XFILLER_27_898 VPWR VGND sg13g2_decap_8
XFILLER_41_301 VPWR VGND sg13g2_decap_8
XFILLER_42_868 VPWR VGND sg13g2_decap_8
XFILLER_41_378 VPWR VGND sg13g2_decap_8
XFILLER_5_213 VPWR VGND sg13g2_decap_8
XFILLER_10_765 VPWR VGND sg13g2_decap_8
XFILLER_6_747 VPWR VGND sg13g2_decap_8
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_30_84 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_7_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_18_843 VPWR VGND sg13g2_decap_8
XFILLER_45_651 VPWR VGND sg13g2_decap_8
XFILLER_17_353 VPWR VGND sg13g2_decap_8
XFILLER_44_161 VPWR VGND sg13g2_decap_8
XFILLER_32_301 VPWR VGND sg13g2_decap_8
XFILLER_33_868 VPWR VGND sg13g2_decap_8
XFILLER_20_518 VPWR VGND sg13g2_decap_8
XFILLER_32_378 VPWR VGND sg13g2_decap_8
XFILLER_9_552 VPWR VGND sg13g2_decap_8
XFILLER_5_780 VPWR VGND sg13g2_decap_8
XFILLER_27_128 VPWR VGND sg13g2_decap_8
XFILLER_24_802 VPWR VGND sg13g2_decap_8
XFILLER_36_651 VPWR VGND sg13g2_decap_8
XFILLER_23_312 VPWR VGND sg13g2_decap_8
XFILLER_35_161 VPWR VGND sg13g2_decap_8
XFILLER_24_879 VPWR VGND sg13g2_decap_8
XFILLER_11_518 VPWR VGND sg13g2_decap_8
XFILLER_23_389 VPWR VGND sg13g2_decap_8
XFILLER_13_1007 VPWR VGND sg13g2_decap_8
XFILLER_3_739 VPWR VGND sg13g2_decap_8
XFILLER_2_238 VPWR VGND sg13g2_decap_8
XFILLER_47_938 VPWR VGND sg13g2_decap_8
XFILLER_19_629 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_15_813 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_decap_8
XFILLER_27_695 VPWR VGND sg13g2_decap_8
XFILLER_42_665 VPWR VGND sg13g2_decap_8
XFILLER_14_345 VPWR VGND sg13g2_decap_8
XFILLER_30_805 VPWR VGND sg13g2_decap_8
XFILLER_25_95 VPWR VGND sg13g2_decap_8
XFILLER_41_175 VPWR VGND sg13g2_decap_8
XFILLER_10_562 VPWR VGND sg13g2_decap_8
XFILLER_6_544 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
X_53_ VPWR VGND _08_ _09_ _21_ _10_ _07_ _11_ sg13g2_a221oi_1
XFILLER_38_938 VPWR VGND sg13g2_decap_8
XFILLER_37_448 VPWR VGND sg13g2_decap_8
XFILLER_18_640 VPWR VGND sg13g2_decap_8
XFILLER_17_150 VPWR VGND sg13g2_decap_8
XFILLER_24_109 VPWR VGND sg13g2_decap_8
XFILLER_33_665 VPWR VGND sg13g2_decap_8
XFILLER_20_315 VPWR VGND sg13g2_decap_8
XFILLER_32_175 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_29_949 VPWR VGND sg13g2_decap_8
XFILLER_28_459 VPWR VGND sg13g2_decap_8
XFILLER_24_676 VPWR VGND sg13g2_decap_8
XFILLER_11_315 VPWR VGND sg13g2_decap_8
XFILLER_12_849 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_decap_8
XFILLER_20_882 VPWR VGND sg13g2_decap_8
XFILLER_11_20 VPWR VGND sg13g2_fill_1
XFILLER_3_536 VPWR VGND sg13g2_decap_8
XFILLER_11_53 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1016 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_19_426 VPWR VGND sg13g2_decap_8
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_15_610 VPWR VGND sg13g2_decap_8
XFILLER_43_952 VPWR VGND sg13g2_decap_8
XFILLER_27_492 VPWR VGND sg13g2_decap_8
XFILLER_42_462 VPWR VGND sg13g2_decap_8
XFILLER_14_142 VPWR VGND sg13g2_decap_8
XFILLER_15_687 VPWR VGND sg13g2_decap_8
XFILLER_30_602 VPWR VGND sg13g2_decap_8
XFILLER_30_679 VPWR VGND sg13g2_decap_8
XFILLER_7_831 VPWR VGND sg13g2_decap_8
XFILLER_11_882 VPWR VGND sg13g2_decap_8
XFILLER_6_341 VPWR VGND sg13g2_decap_8
XFILLER_42_1022 VPWR VGND sg13g2_decap_8
XFILLER_38_735 VPWR VGND sg13g2_decap_8
X_36_ net1 VPWR _13_ VGND net46 _12_ sg13g2_o21ai_1
XFILLER_37_245 VPWR VGND sg13g2_decap_8
XFILLER_19_993 VPWR VGND sg13g2_decap_8
XFILLER_34_952 VPWR VGND sg13g2_decap_8
XFILLER_33_462 VPWR VGND sg13g2_decap_8
XFILLER_20_112 VPWR VGND sg13g2_decap_8
XFILLER_21_668 VPWR VGND sg13g2_decap_8
XFILLER_20_189 VPWR VGND sg13g2_decap_8
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_29_746 VPWR VGND sg13g2_decap_8
XFILLER_28_256 VPWR VGND sg13g2_decap_8
XFILLER_44_749 VPWR VGND sg13g2_decap_8
XFILLER_43_259 VPWR VGND sg13g2_decap_8
XFILLER_25_963 VPWR VGND sg13g2_decap_8
XFILLER_12_646 VPWR VGND sg13g2_decap_8
XFILLER_24_473 VPWR VGND sg13g2_decap_8
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_8_639 VPWR VGND sg13g2_decap_8
XFILLER_7_138 VPWR VGND sg13g2_decap_8
XFILLER_11_189 VPWR VGND sg13g2_decap_8
XFILLER_4_834 VPWR VGND sg13g2_decap_8
XFILLER_3_333 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_19_223 VPWR VGND sg13g2_decap_8
XFILLER_16_930 VPWR VGND sg13g2_decap_8
XFILLER_35_749 VPWR VGND sg13g2_decap_8
XFILLER_34_259 VPWR VGND sg13g2_decap_8
XFILLER_15_484 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
XFILLER_31_966 VPWR VGND sg13g2_decap_8
XFILLER_30_476 VPWR VGND sg13g2_decap_8
X_55__25 VPWR VGND net24 sg13g2_tiehi
XFILLER_38_532 VPWR VGND sg13g2_decap_8
XFILLER_19_790 VPWR VGND sg13g2_decap_8
XFILLER_22_933 VPWR VGND sg13g2_decap_8
XFILLER_21_465 VPWR VGND sg13g2_decap_8
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_826 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_29_543 VPWR VGND sg13g2_decap_8
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_17_738 VPWR VGND sg13g2_decap_8
XFILLER_44_546 VPWR VGND sg13g2_decap_8
XFILLER_16_237 VPWR VGND sg13g2_decap_8
XFILLER_17_63 VPWR VGND sg13g2_decap_8
XFILLER_25_760 VPWR VGND sg13g2_decap_8
XFILLER_13_944 VPWR VGND sg13g2_decap_8
XFILLER_24_270 VPWR VGND sg13g2_decap_8
XFILLER_12_443 VPWR VGND sg13g2_decap_8
XFILLER_40_763 VPWR VGND sg13g2_decap_8
XFILLER_8_436 VPWR VGND sg13g2_decap_8
XFILLER_9_937 VPWR VGND sg13g2_decap_8
XFILLER_33_84 VPWR VGND sg13g2_decap_8
XFILLER_4_631 VPWR VGND sg13g2_decap_8
XFILLER_3_130 VPWR VGND sg13g2_decap_8
XFILLER_39_329 VPWR VGND sg13g2_decap_8
XFILLER_48_896 VPWR VGND sg13g2_decap_8
XFILLER_35_546 VPWR VGND sg13g2_decap_8
XFILLER_15_281 VPWR VGND sg13g2_decap_8
XFILLER_31_763 VPWR VGND sg13g2_decap_8
XFILLER_30_273 VPWR VGND sg13g2_decap_8
XFILLER_39_896 VPWR VGND sg13g2_decap_8
XFILLER_26_557 VPWR VGND sg13g2_decap_8
XFILLER_22_730 VPWR VGND sg13g2_decap_8
XFILLER_21_262 VPWR VGND sg13g2_decap_8
XFILLER_10_947 VPWR VGND sg13g2_decap_8
XFILLER_6_929 VPWR VGND sg13g2_decap_8
XFILLER_1_623 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_49_627 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_29_340 VPWR VGND sg13g2_decap_8
XFILLER_45_833 VPWR VGND sg13g2_decap_8
XFILLER_17_535 VPWR VGND sg13g2_decap_8
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_44_343 VPWR VGND sg13g2_decap_8
XFILLER_13_741 VPWR VGND sg13g2_decap_8
XFILLER_9_734 VPWR VGND sg13g2_decap_8
XFILLER_12_240 VPWR VGND sg13g2_decap_8
XFILLER_40_560 VPWR VGND sg13g2_decap_8
XFILLER_8_233 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_5_962 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_fill_1
XFILLER_5_77 VPWR VGND sg13g2_decap_8
XFILLER_39_126 VPWR VGND sg13g2_decap_8
XFILLER_48_693 VPWR VGND sg13g2_decap_8
XFILLER_36_833 VPWR VGND sg13g2_decap_8
XFILLER_35_343 VPWR VGND sg13g2_decap_8
XFILLER_31_560 VPWR VGND sg13g2_decap_8
XFILLER_49_39 VPWR VGND sg13g2_decap_8
XFILLER_27_800 VPWR VGND sg13g2_decap_8
XFILLER_39_693 VPWR VGND sg13g2_decap_8
XFILLER_26_354 VPWR VGND sg13g2_decap_8
XFILLER_27_877 VPWR VGND sg13g2_decap_8
XFILLER_42_847 VPWR VGND sg13g2_decap_8
XFILLER_14_527 VPWR VGND sg13g2_decap_8
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_10_744 VPWR VGND sg13g2_decap_8
XFILLER_14_64 VPWR VGND sg13g2_decap_8
XFILLER_6_726 VPWR VGND sg13g2_decap_8
XFILLER_5_269 VPWR VGND sg13g2_decap_8
XFILLER_30_63 VPWR VGND sg13g2_decap_8
XFILLER_2_910 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_49_424 VPWR VGND sg13g2_decap_8
XFILLER_2_987 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_45_630 VPWR VGND sg13g2_decap_8
XFILLER_18_822 VPWR VGND sg13g2_decap_8
XFILLER_44_140 VPWR VGND sg13g2_decap_8
XFILLER_17_332 VPWR VGND sg13g2_decap_8
XFILLER_18_899 VPWR VGND sg13g2_decap_8
XFILLER_33_847 VPWR VGND sg13g2_decap_8
XFILLER_32_357 VPWR VGND sg13g2_decap_8
XFILLER_9_531 VPWR VGND sg13g2_decap_8
XFILLER_27_107 VPWR VGND sg13g2_decap_8
XFILLER_49_991 VPWR VGND sg13g2_decap_8
XFILLER_48_490 VPWR VGND sg13g2_decap_8
XFILLER_36_630 VPWR VGND sg13g2_decap_8
XFILLER_35_140 VPWR VGND sg13g2_decap_8
XFILLER_24_858 VPWR VGND sg13g2_decap_8
XFILLER_23_368 VPWR VGND sg13g2_decap_8
XFILLER_3_718 VPWR VGND sg13g2_decap_8
XFILLER_2_217 VPWR VGND sg13g2_decap_8
XFILLER_47_917 VPWR VGND sg13g2_decap_8
XFILLER_19_608 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_39_490 VPWR VGND sg13g2_decap_8
XFILLER_26_151 VPWR VGND sg13g2_decap_8
XFILLER_27_674 VPWR VGND sg13g2_decap_8
XFILLER_42_644 VPWR VGND sg13g2_decap_8
XFILLER_14_324 VPWR VGND sg13g2_decap_8
XFILLER_15_869 VPWR VGND sg13g2_decap_8
XFILLER_25_74 VPWR VGND sg13g2_decap_8
XFILLER_41_154 VPWR VGND sg13g2_decap_8
XFILLER_10_541 VPWR VGND sg13g2_decap_8
XFILLER_6_523 VPWR VGND sg13g2_decap_8
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_29_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_784 VPWR VGND sg13g2_decap_8
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
X_52_ net42 _22_ _06_ VPWR VGND sg13g2_nor2_1
XFILLER_38_917 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
XFILLER_37_427 VPWR VGND sg13g2_decap_8
XFILLER_46_994 VPWR VGND sg13g2_decap_8
XFILLER_18_696 VPWR VGND sg13g2_decap_8
XFILLER_33_644 VPWR VGND sg13g2_decap_8
XFILLER_36_1008 VPWR VGND sg13g2_decap_8
XFILLER_32_154 VPWR VGND sg13g2_decap_8
XFILLER_14_891 VPWR VGND sg13g2_decap_8
XFILLER_29_928 VPWR VGND sg13g2_decap_8
XFILLER_28_438 VPWR VGND sg13g2_decap_8
XFILLER_37_994 VPWR VGND sg13g2_decap_8
XFILLER_24_655 VPWR VGND sg13g2_decap_8
XFILLER_12_828 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_20_861 VPWR VGND sg13g2_decap_8
XFILLER_11_32 VPWR VGND sg13g2_decap_4
XFILLER_3_515 VPWR VGND sg13g2_decap_8
XFILLER_47_714 VPWR VGND sg13g2_decap_8
XFILLER_19_405 VPWR VGND sg13g2_decap_8
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_27_471 VPWR VGND sg13g2_decap_8
XFILLER_43_931 VPWR VGND sg13g2_decap_8
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_42_441 VPWR VGND sg13g2_decap_8
XFILLER_14_132 VPWR VGND sg13g2_fill_1
XFILLER_15_666 VPWR VGND sg13g2_decap_8
XFILLER_14_198 VPWR VGND sg13g2_decap_8
XFILLER_7_810 VPWR VGND sg13g2_decap_8
XFILLER_11_861 VPWR VGND sg13g2_decap_8
XFILLER_30_658 VPWR VGND sg13g2_decap_8
XFILLER_6_320 VPWR VGND sg13g2_decap_8
XFILLER_7_887 VPWR VGND sg13g2_decap_8
XFILLER_6_397 VPWR VGND sg13g2_decap_8
XFILLER_42_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_581 VPWR VGND sg13g2_decap_8
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_38_714 VPWR VGND sg13g2_decap_8
XFILLER_37_224 VPWR VGND sg13g2_decap_8
X_35_ _10_ _11_ _12_ VPWR VGND sg13g2_and2_1
XFILLER_19_972 VPWR VGND sg13g2_decap_8
XFILLER_46_791 VPWR VGND sg13g2_decap_8
XFILLER_18_493 VPWR VGND sg13g2_decap_8
XFILLER_34_931 VPWR VGND sg13g2_decap_8
XFILLER_33_441 VPWR VGND sg13g2_decap_8
XFILLER_21_647 VPWR VGND sg13g2_decap_8
XFILLER_20_168 VPWR VGND sg13g2_decap_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_29_725 VPWR VGND sg13g2_decap_8
XFILLER_28_235 VPWR VGND sg13g2_decap_8
XFILLER_44_728 VPWR VGND sg13g2_decap_8
XFILLER_16_419 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_25_942 VPWR VGND sg13g2_decap_8
XFILLER_37_791 VPWR VGND sg13g2_decap_8
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_24_452 VPWR VGND sg13g2_decap_8
XFILLER_12_625 VPWR VGND sg13g2_decap_8
XFILLER_40_945 VPWR VGND sg13g2_decap_8
XFILLER_8_618 VPWR VGND sg13g2_decap_8
XFILLER_7_117 VPWR VGND sg13g2_decap_8
XFILLER_11_168 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_4_813 VPWR VGND sg13g2_decap_8
XFILLER_3_312 VPWR VGND sg13g2_decap_8
XFILLER_3_389 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_19_202 VPWR VGND sg13g2_decap_8
XFILLER_47_588 VPWR VGND sg13g2_decap_8
XFILLER_19_279 VPWR VGND sg13g2_decap_8
XFILLER_35_728 VPWR VGND sg13g2_decap_8
XFILLER_34_238 VPWR VGND sg13g2_decap_8
XFILLER_15_463 VPWR VGND sg13g2_decap_8
XFILLER_16_986 VPWR VGND sg13g2_decap_8
XFILLER_31_945 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_30_455 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_decap_8
XFILLER_7_684 VPWR VGND sg13g2_decap_8
XFILLER_6_194 VPWR VGND sg13g2_decap_8
XFILLER_38_511 VPWR VGND sg13g2_decap_8
XFILLER_26_739 VPWR VGND sg13g2_decap_8
XFILLER_38_588 VPWR VGND sg13g2_decap_8
XFILLER_25_249 VPWR VGND sg13g2_decap_8
XFILLER_18_290 VPWR VGND sg13g2_decap_8
XFILLER_22_912 VPWR VGND sg13g2_decap_8
XFILLER_21_444 VPWR VGND sg13g2_decap_8
XFILLER_22_989 VPWR VGND sg13g2_decap_8
XFILLER_1_805 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_49_809 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_29_522 VPWR VGND sg13g2_decap_8
XFILLER_17_717 VPWR VGND sg13g2_decap_8
XFILLER_44_525 VPWR VGND sg13g2_decap_8
XFILLER_16_216 VPWR VGND sg13g2_decap_8
XFILLER_29_599 VPWR VGND sg13g2_decap_8
XFILLER_13_923 VPWR VGND sg13g2_decap_8
XFILLER_9_916 VPWR VGND sg13g2_decap_8
XFILLER_12_422 VPWR VGND sg13g2_decap_8
XFILLER_40_742 VPWR VGND sg13g2_decap_8
XFILLER_8_415 VPWR VGND sg13g2_decap_8
XFILLER_32_1022 VPWR VGND sg13g2_decap_8
XFILLER_33_63 VPWR VGND sg13g2_decap_8
XFILLER_12_499 VPWR VGND sg13g2_decap_8
XFILLER_4_610 VPWR VGND sg13g2_decap_8
XFILLER_4_687 VPWR VGND sg13g2_decap_8
XFILLER_3_186 VPWR VGND sg13g2_decap_8
XFILLER_39_308 VPWR VGND sg13g2_decap_8
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_48_875 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_35_525 VPWR VGND sg13g2_decap_8
XFILLER_15_260 VPWR VGND sg13g2_decap_8
XFILLER_16_783 VPWR VGND sg13g2_decap_8
XFILLER_22_219 VPWR VGND sg13g2_decap_8
XFILLER_31_742 VPWR VGND sg13g2_decap_8
XFILLER_30_252 VPWR VGND sg13g2_decap_8
XFILLER_8_982 VPWR VGND sg13g2_decap_8
XFILLER_7_481 VPWR VGND sg13g2_decap_8
XFILLER_39_875 VPWR VGND sg13g2_decap_8
XFILLER_26_536 VPWR VGND sg13g2_decap_8
XFILLER_38_385 VPWR VGND sg13g2_decap_8
XFILLER_14_709 VPWR VGND sg13g2_decap_8
XFILLER_41_539 VPWR VGND sg13g2_decap_8
XFILLER_10_926 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_241 VPWR VGND sg13g2_decap_8
XFILLER_22_786 VPWR VGND sg13g2_decap_8
XFILLER_6_908 VPWR VGND sg13g2_decap_8
XFILLER_1_602 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_49_606 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_45_812 VPWR VGND sg13g2_decap_8
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_44_322 VPWR VGND sg13g2_decap_8
XFILLER_17_514 VPWR VGND sg13g2_decap_8
XFILLER_29_396 VPWR VGND sg13g2_decap_8
XFILLER_45_889 VPWR VGND sg13g2_decap_8
XFILLER_44_399 VPWR VGND sg13g2_decap_8
XFILLER_13_720 VPWR VGND sg13g2_decap_8
XFILLER_32_539 VPWR VGND sg13g2_decap_8
XFILLER_44_84 VPWR VGND sg13g2_decap_8
XFILLER_8_212 VPWR VGND sg13g2_decap_8
XFILLER_9_713 VPWR VGND sg13g2_decap_8
XFILLER_12_296 VPWR VGND sg13g2_decap_8
XFILLER_13_797 VPWR VGND sg13g2_decap_8
XFILLER_8_289 VPWR VGND sg13g2_decap_8
XFILLER_5_941 VPWR VGND sg13g2_decap_8
XFILLER_5_56 VPWR VGND sg13g2_decap_8
XFILLER_4_484 VPWR VGND sg13g2_decap_8
XFILLER_39_105 VPWR VGND sg13g2_decap_8
XFILLER_48_672 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_36_812 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
XFILLER_35_322 VPWR VGND sg13g2_decap_8
XFILLER_36_889 VPWR VGND sg13g2_decap_8
XFILLER_35_399 VPWR VGND sg13g2_decap_8
XFILLER_16_580 VPWR VGND sg13g2_decap_8
XFILLER_49_18 VPWR VGND sg13g2_decap_8
XFILLER_46_609 VPWR VGND sg13g2_decap_8
XFILLER_22_1010 VPWR VGND sg13g2_decap_8
XFILLER_39_672 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_26_333 VPWR VGND sg13g2_decap_8
XFILLER_27_856 VPWR VGND sg13g2_decap_8
XFILLER_42_826 VPWR VGND sg13g2_decap_8
XFILLER_14_506 VPWR VGND sg13g2_decap_8
XFILLER_41_336 VPWR VGND sg13g2_decap_8
XFILLER_14_43 VPWR VGND sg13g2_decap_8
XFILLER_10_723 VPWR VGND sg13g2_decap_8
XFILLER_22_583 VPWR VGND sg13g2_decap_8
XFILLER_6_705 VPWR VGND sg13g2_decap_8
XFILLER_5_248 VPWR VGND sg13g2_decap_8
XFILLER_30_42 VPWR VGND sg13g2_decap_8
XFILLER_2_966 VPWR VGND sg13g2_decap_8
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_decap_8
XFILLER_18_801 VPWR VGND sg13g2_decap_8
XFILLER_37_609 VPWR VGND sg13g2_decap_8
XFILLER_17_311 VPWR VGND sg13g2_decap_8
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_18_878 VPWR VGND sg13g2_decap_8
XFILLER_29_193 VPWR VGND sg13g2_decap_8
XFILLER_45_686 VPWR VGND sg13g2_decap_8
XFILLER_17_388 VPWR VGND sg13g2_decap_8
XFILLER_33_826 VPWR VGND sg13g2_decap_8
XFILLER_44_196 VPWR VGND sg13g2_decap_8
XFILLER_32_336 VPWR VGND sg13g2_decap_8
XFILLER_9_510 VPWR VGND sg13g2_decap_8
XFILLER_13_594 VPWR VGND sg13g2_decap_8
XFILLER_9_587 VPWR VGND sg13g2_decap_8
XFILLER_4_281 VPWR VGND sg13g2_decap_8
XFILLER_49_970 VPWR VGND sg13g2_decap_8
XFILLER_24_837 VPWR VGND sg13g2_decap_8
XFILLER_36_686 VPWR VGND sg13g2_decap_8
XFILLER_23_347 VPWR VGND sg13g2_decap_8
XFILLER_35_196 VPWR VGND sg13g2_decap_8
XFILLER_46_406 VPWR VGND sg13g2_decap_8
XFILLER_26_130 VPWR VGND sg13g2_decap_8
XFILLER_27_653 VPWR VGND sg13g2_decap_8
XFILLER_14_303 VPWR VGND sg13g2_decap_8
XFILLER_42_623 VPWR VGND sg13g2_decap_8
XFILLER_15_848 VPWR VGND sg13g2_decap_8
XFILLER_25_53 VPWR VGND sg13g2_decap_8
XFILLER_41_133 VPWR VGND sg13g2_decap_8
XFILLER_10_520 VPWR VGND sg13g2_decap_8
XFILLER_22_380 VPWR VGND sg13g2_decap_8
XFILLER_6_502 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_10_597 VPWR VGND sg13g2_decap_8
XFILLER_6_579 VPWR VGND sg13g2_decap_8
XFILLER_29_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_763 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
X_51_ _22_ net1 _21_ VPWR VGND sg13g2_nand2_1
XFILLER_37_406 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_2_79 VPWR VGND sg13g2_decap_8
XFILLER_46_973 VPWR VGND sg13g2_decap_8
XFILLER_18_675 VPWR VGND sg13g2_decap_8
XFILLER_45_483 VPWR VGND sg13g2_decap_8
XFILLER_17_185 VPWR VGND sg13g2_decap_8
XFILLER_33_623 VPWR VGND sg13g2_decap_8
XFILLER_21_829 VPWR VGND sg13g2_decap_8
XFILLER_32_133 VPWR VGND sg13g2_decap_8
XFILLER_14_870 VPWR VGND sg13g2_decap_8
XFILLER_13_391 VPWR VGND sg13g2_decap_8
XFILLER_9_384 VPWR VGND sg13g2_decap_8
XFILLER_29_907 VPWR VGND sg13g2_decap_8
XFILLER_28_417 VPWR VGND sg13g2_decap_8
XFILLER_37_973 VPWR VGND sg13g2_decap_8
XFILLER_24_634 VPWR VGND sg13g2_decap_8
XFILLER_36_483 VPWR VGND sg13g2_decap_8
XFILLER_12_807 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_20_840 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_11_88 VPWR VGND sg13g2_decap_8
XFILLER_11_99 VPWR VGND sg13g2_fill_2
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_43_910 VPWR VGND sg13g2_decap_8
XFILLER_27_450 VPWR VGND sg13g2_decap_8
XFILLER_28_984 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_42_420 VPWR VGND sg13g2_decap_8
XFILLER_15_645 VPWR VGND sg13g2_decap_8
XFILLER_43_987 VPWR VGND sg13g2_decap_8
XFILLER_42_497 VPWR VGND sg13g2_decap_8
XFILLER_14_177 VPWR VGND sg13g2_decap_8
XFILLER_30_637 VPWR VGND sg13g2_decap_8
XFILLER_11_840 VPWR VGND sg13g2_decap_8
XFILLER_10_394 VPWR VGND sg13g2_decap_8
XFILLER_7_866 VPWR VGND sg13g2_decap_8
XFILLER_6_376 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_8
XFILLER_2_560 VPWR VGND sg13g2_decap_8
XFILLER_37_203 VPWR VGND sg13g2_decap_8
X_34_ _11_ net44 net41 net5 VPWR VGND sg13g2_and3_1
XFILLER_19_951 VPWR VGND sg13g2_decap_8
XFILLER_46_770 VPWR VGND sg13g2_decap_8
XFILLER_34_910 VPWR VGND sg13g2_decap_8
XFILLER_45_280 VPWR VGND sg13g2_decap_8
XFILLER_18_472 VPWR VGND sg13g2_decap_8
XFILLER_33_420 VPWR VGND sg13g2_decap_8
XFILLER_34_987 VPWR VGND sg13g2_decap_8
XFILLER_21_626 VPWR VGND sg13g2_decap_8
XFILLER_33_497 VPWR VGND sg13g2_decap_8
XFILLER_20_147 VPWR VGND sg13g2_decap_8
XFILLER_9_181 VPWR VGND sg13g2_decap_8
XFILLER_29_704 VPWR VGND sg13g2_decap_8
XFILLER_28_214 VPWR VGND sg13g2_decap_8
XFILLER_44_707 VPWR VGND sg13g2_decap_8
XFILLER_37_770 VPWR VGND sg13g2_decap_8
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_25_921 VPWR VGND sg13g2_decap_8
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_12_604 VPWR VGND sg13g2_decap_8
XFILLER_24_431 VPWR VGND sg13g2_decap_8
XFILLER_25_998 VPWR VGND sg13g2_decap_8
XFILLER_40_924 VPWR VGND sg13g2_decap_8
XFILLER_11_147 VPWR VGND sg13g2_decap_8
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_4_869 VPWR VGND sg13g2_decap_8
XFILLER_3_368 VPWR VGND sg13g2_decap_8
XFILLER_26_1019 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
XFILLER_19_258 VPWR VGND sg13g2_decap_8
XFILLER_35_707 VPWR VGND sg13g2_decap_8
XFILLER_28_781 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_decap_8
XFILLER_15_442 VPWR VGND sg13g2_decap_8
XFILLER_16_965 VPWR VGND sg13g2_decap_8
XFILLER_43_784 VPWR VGND sg13g2_decap_8
XFILLER_31_924 VPWR VGND sg13g2_decap_8
XFILLER_42_294 VPWR VGND sg13g2_decap_8
XFILLER_30_434 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
XFILLER_10_191 VPWR VGND sg13g2_decap_8
XFILLER_7_663 VPWR VGND sg13g2_decap_8
XFILLER_6_173 VPWR VGND sg13g2_decap_8
XFILLER_26_718 VPWR VGND sg13g2_decap_8
XFILLER_38_567 VPWR VGND sg13g2_decap_8
XFILLER_25_228 VPWR VGND sg13g2_decap_8
XFILLER_34_784 VPWR VGND sg13g2_decap_8
XFILLER_21_423 VPWR VGND sg13g2_decap_8
XFILLER_22_968 VPWR VGND sg13g2_decap_8
XFILLER_33_294 VPWR VGND sg13g2_decap_8
XFILLER_49_1019 VPWR VGND sg13g2_decap_8
XFILLER_29_501 VPWR VGND sg13g2_decap_8
XFILLER_44_504 VPWR VGND sg13g2_decap_8
XFILLER_17_21 VPWR VGND sg13g2_fill_1
XFILLER_29_578 VPWR VGND sg13g2_decap_8
XFILLER_13_902 VPWR VGND sg13g2_decap_8
XFILLER_17_98 VPWR VGND sg13g2_decap_8
XFILLER_12_401 VPWR VGND sg13g2_decap_8
XFILLER_25_795 VPWR VGND sg13g2_decap_8
XFILLER_40_721 VPWR VGND sg13g2_decap_8
XFILLER_33_42 VPWR VGND sg13g2_decap_8
XFILLER_12_478 VPWR VGND sg13g2_decap_8
XFILLER_13_979 VPWR VGND sg13g2_decap_8
XFILLER_32_1001 VPWR VGND sg13g2_decap_8
XFILLER_21_990 VPWR VGND sg13g2_decap_8
XFILLER_40_798 VPWR VGND sg13g2_decap_8
XFILLER_4_666 VPWR VGND sg13g2_decap_8
XFILLER_3_165 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_48_854 VPWR VGND sg13g2_decap_8
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_35_504 VPWR VGND sg13g2_decap_8
XFILLER_16_762 VPWR VGND sg13g2_decap_8
XFILLER_31_721 VPWR VGND sg13g2_decap_8
XFILLER_43_581 VPWR VGND sg13g2_decap_8
XFILLER_30_231 VPWR VGND sg13g2_decap_8
XFILLER_31_798 VPWR VGND sg13g2_decap_8
XFILLER_8_961 VPWR VGND sg13g2_decap_8
XFILLER_7_460 VPWR VGND sg13g2_decap_8
XFILLER_31_0 VPWR VGND sg13g2_decap_8
XFILLER_39_854 VPWR VGND sg13g2_decap_8
XFILLER_38_364 VPWR VGND sg13g2_decap_8
XFILLER_26_515 VPWR VGND sg13g2_decap_8
XFILLER_41_518 VPWR VGND sg13g2_decap_8
XFILLER_13_209 VPWR VGND sg13g2_decap_8
XFILLER_16_1007 VPWR VGND sg13g2_decap_8
XFILLER_21_220 VPWR VGND sg13g2_decap_8
XFILLER_34_581 VPWR VGND sg13g2_decap_8
XFILLER_10_905 VPWR VGND sg13g2_decap_8
XFILLER_22_765 VPWR VGND sg13g2_decap_8
XFILLER_21_297 VPWR VGND sg13g2_decap_8
XFILLER_1_658 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_44_301 VPWR VGND sg13g2_decap_8
XFILLER_29_375 VPWR VGND sg13g2_decap_8
XFILLER_45_868 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_8
XFILLER_32_518 VPWR VGND sg13g2_decap_8
XFILLER_44_63 VPWR VGND sg13g2_decap_8
XFILLER_25_592 VPWR VGND sg13g2_decap_8
XFILLER_13_776 VPWR VGND sg13g2_decap_8
XFILLER_9_769 VPWR VGND sg13g2_decap_8
XFILLER_12_275 VPWR VGND sg13g2_decap_8
XFILLER_40_595 VPWR VGND sg13g2_decap_8
XFILLER_8_268 VPWR VGND sg13g2_decap_8
XFILLER_5_920 VPWR VGND sg13g2_decap_8
XFILLER_5_997 VPWR VGND sg13g2_decap_8
XFILLER_4_463 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_decap_8
XFILLER_36_868 VPWR VGND sg13g2_decap_8
XFILLER_23_529 VPWR VGND sg13g2_decap_8
XFILLER_35_378 VPWR VGND sg13g2_decap_8
XFILLER_31_595 VPWR VGND sg13g2_decap_8
XFILLER_39_651 VPWR VGND sg13g2_decap_8
XFILLER_26_312 VPWR VGND sg13g2_decap_8
XFILLER_27_835 VPWR VGND sg13g2_decap_8
XFILLER_38_161 VPWR VGND sg13g2_decap_8
XFILLER_42_805 VPWR VGND sg13g2_decap_8
XFILLER_26_389 VPWR VGND sg13g2_decap_8
XFILLER_41_315 VPWR VGND sg13g2_decap_8
XFILLER_14_11 VPWR VGND sg13g2_decap_4
XFILLER_10_702 VPWR VGND sg13g2_decap_8
XFILLER_22_562 VPWR VGND sg13g2_decap_8
XFILLER_10_779 VPWR VGND sg13g2_decap_8
XFILLER_5_227 VPWR VGND sg13g2_decap_8
XFILLER_30_21 VPWR VGND sg13g2_decap_8
XFILLER_30_98 VPWR VGND sg13g2_decap_8
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_29_172 VPWR VGND sg13g2_decap_8
XFILLER_18_857 VPWR VGND sg13g2_decap_8
XFILLER_45_665 VPWR VGND sg13g2_decap_8
XFILLER_17_367 VPWR VGND sg13g2_decap_8
XFILLER_33_805 VPWR VGND sg13g2_decap_8
XFILLER_44_175 VPWR VGND sg13g2_decap_8
XFILLER_32_315 VPWR VGND sg13g2_decap_8
XFILLER_41_882 VPWR VGND sg13g2_decap_8
XFILLER_13_573 VPWR VGND sg13g2_decap_8
XFILLER_9_566 VPWR VGND sg13g2_decap_8
XFILLER_40_392 VPWR VGND sg13g2_decap_8
XFILLER_4_260 VPWR VGND sg13g2_decap_8
XFILLER_5_794 VPWR VGND sg13g2_decap_8
XFILLER_45_1022 VPWR VGND sg13g2_decap_8
XFILLER_24_816 VPWR VGND sg13g2_decap_8
XFILLER_36_665 VPWR VGND sg13g2_decap_8
XFILLER_23_326 VPWR VGND sg13g2_decap_8
XFILLER_35_175 VPWR VGND sg13g2_decap_8
XFILLER_32_882 VPWR VGND sg13g2_decap_8
XFILLER_31_392 VPWR VGND sg13g2_decap_8
XFILLER_18_109 VPWR VGND sg13g2_decap_8
XFILLER_27_632 VPWR VGND sg13g2_decap_8
XFILLER_42_602 VPWR VGND sg13g2_decap_8
XFILLER_15_827 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_26_186 VPWR VGND sg13g2_decap_8
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_42_679 VPWR VGND sg13g2_decap_8
XFILLER_14_359 VPWR VGND sg13g2_decap_8
XFILLER_30_819 VPWR VGND sg13g2_decap_8
XFILLER_23_893 VPWR VGND sg13g2_decap_8
XFILLER_41_189 VPWR VGND sg13g2_decap_8
XFILLER_10_576 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_6_558 VPWR VGND sg13g2_decap_8
XFILLER_2_742 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_4
XFILLER_49_256 VPWR VGND sg13g2_decap_8
X_50_ net5 _10_ net41 _21_ VPWR VGND sg13g2_nand3_1
XFILLER_2_58 VPWR VGND sg13g2_decap_8
XFILLER_46_952 VPWR VGND sg13g2_decap_8
XFILLER_18_654 VPWR VGND sg13g2_decap_8
XFILLER_45_462 VPWR VGND sg13g2_decap_8
XFILLER_17_164 VPWR VGND sg13g2_decap_8
XFILLER_33_602 VPWR VGND sg13g2_decap_8
XFILLER_32_112 VPWR VGND sg13g2_decap_8
XFILLER_21_808 VPWR VGND sg13g2_decap_8
XFILLER_33_679 VPWR VGND sg13g2_decap_8
XFILLER_13_370 VPWR VGND sg13g2_decap_8
XFILLER_20_329 VPWR VGND sg13g2_decap_8
XFILLER_32_189 VPWR VGND sg13g2_decap_8
XFILLER_9_363 VPWR VGND sg13g2_decap_8
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
XFILLER_5_591 VPWR VGND sg13g2_decap_8
XFILLER_37_952 VPWR VGND sg13g2_decap_8
XFILLER_36_462 VPWR VGND sg13g2_decap_8
XFILLER_24_613 VPWR VGND sg13g2_decap_8
XFILLER_23_123 VPWR VGND sg13g2_decap_8
XFILLER_11_329 VPWR VGND sg13g2_decap_8
XFILLER_20_896 VPWR VGND sg13g2_decap_8
XFILLER_11_67 VPWR VGND sg13g2_decap_8
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_28_963 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_15_624 VPWR VGND sg13g2_decap_8
XFILLER_43_966 VPWR VGND sg13g2_decap_8
XFILLER_42_476 VPWR VGND sg13g2_decap_8
XFILLER_14_156 VPWR VGND sg13g2_decap_8
XFILLER_30_616 VPWR VGND sg13g2_decap_8
XFILLER_23_690 VPWR VGND sg13g2_decap_8
XFILLER_10_373 VPWR VGND sg13g2_decap_8
XFILLER_7_845 VPWR VGND sg13g2_decap_8
XFILLER_11_896 VPWR VGND sg13g2_decap_8
XFILLER_6_355 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
X_33_ _10_ net2 net34 net3 VPWR VGND sg13g2_and3_1
XFILLER_19_930 VPWR VGND sg13g2_decap_8
XFILLER_38_749 VPWR VGND sg13g2_decap_8
XFILLER_18_451 VPWR VGND sg13g2_decap_8
XFILLER_37_259 VPWR VGND sg13g2_decap_8
XFILLER_34_966 VPWR VGND sg13g2_decap_8
XFILLER_21_605 VPWR VGND sg13g2_decap_8
XFILLER_33_476 VPWR VGND sg13g2_decap_8
XFILLER_20_126 VPWR VGND sg13g2_decap_8
XFILLER_9_160 VPWR VGND sg13g2_decap_8
XFILLER_25_900 VPWR VGND sg13g2_decap_8
XFILLER_24_410 VPWR VGND sg13g2_decap_8
XFILLER_25_977 VPWR VGND sg13g2_decap_8
XFILLER_40_903 VPWR VGND sg13g2_decap_8
XFILLER_24_487 VPWR VGND sg13g2_decap_8
XFILLER_11_126 VPWR VGND sg13g2_decap_8
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_20_693 VPWR VGND sg13g2_decap_8
XFILLER_4_848 VPWR VGND sg13g2_decap_8
XFILLER_3_347 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_19_237 VPWR VGND sg13g2_decap_8
XFILLER_28_760 VPWR VGND sg13g2_decap_8
XFILLER_16_944 VPWR VGND sg13g2_decap_8
XFILLER_43_763 VPWR VGND sg13g2_decap_8
XFILLER_15_421 VPWR VGND sg13g2_decap_8
XFILLER_31_903 VPWR VGND sg13g2_decap_8
XFILLER_42_273 VPWR VGND sg13g2_decap_8
XFILLER_30_413 VPWR VGND sg13g2_decap_8
XFILLER_15_498 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_fill_2
XFILLER_10_170 VPWR VGND sg13g2_decap_8
XFILLER_7_642 VPWR VGND sg13g2_decap_8
XFILLER_11_693 VPWR VGND sg13g2_decap_8
XFILLER_6_152 VPWR VGND sg13g2_decap_8
XFILLER_38_546 VPWR VGND sg13g2_decap_8
XFILLER_25_207 VPWR VGND sg13g2_decap_8
XFILLER_21_402 VPWR VGND sg13g2_decap_8
XFILLER_34_763 VPWR VGND sg13g2_decap_8
XFILLER_22_947 VPWR VGND sg13g2_decap_8
XFILLER_33_273 VPWR VGND sg13g2_decap_8
XFILLER_21_479 VPWR VGND sg13g2_decap_8
XFILLER_30_980 VPWR VGND sg13g2_decap_8
XFILLER_29_557 VPWR VGND sg13g2_decap_8
XFILLER_17_77 VPWR VGND sg13g2_decap_8
XFILLER_25_774 VPWR VGND sg13g2_decap_8
XFILLER_40_700 VPWR VGND sg13g2_decap_8
XFILLER_13_958 VPWR VGND sg13g2_decap_8
XFILLER_24_284 VPWR VGND sg13g2_decap_8
XFILLER_33_21 VPWR VGND sg13g2_decap_8
XFILLER_12_457 VPWR VGND sg13g2_decap_8
XFILLER_40_777 VPWR VGND sg13g2_decap_8
XFILLER_33_98 VPWR VGND sg13g2_decap_8
XFILLER_20_490 VPWR VGND sg13g2_decap_8
XFILLER_4_645 VPWR VGND sg13g2_decap_8
XFILLER_3_144 VPWR VGND sg13g2_decap_8
X_60__20 VPWR VGND net19 sg13g2_tiehi
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_48_833 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_16_741 VPWR VGND sg13g2_decap_8
XFILLER_43_560 VPWR VGND sg13g2_decap_8
XFILLER_31_700 VPWR VGND sg13g2_decap_8
XFILLER_15_295 VPWR VGND sg13g2_decap_8
XFILLER_30_210 VPWR VGND sg13g2_decap_8
XFILLER_31_777 VPWR VGND sg13g2_decap_8
XFILLER_8_940 VPWR VGND sg13g2_decap_8
XFILLER_30_287 VPWR VGND sg13g2_decap_8
XFILLER_11_490 VPWR VGND sg13g2_decap_8
XFILLER_39_833 VPWR VGND sg13g2_decap_8
XFILLER_38_343 VPWR VGND sg13g2_decap_8
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_34_560 VPWR VGND sg13g2_decap_8
XFILLER_22_744 VPWR VGND sg13g2_decap_8
XFILLER_21_276 VPWR VGND sg13g2_decap_8
XFILLER_5_409 VPWR VGND sg13g2_decap_8
XFILLER_1_637 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_clk clknet_1_1__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_354 VPWR VGND sg13g2_decap_8
XFILLER_45_847 VPWR VGND sg13g2_decap_8
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_17_549 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_25_571 VPWR VGND sg13g2_decap_8
XFILLER_12_254 VPWR VGND sg13g2_decap_8
XFILLER_13_755 VPWR VGND sg13g2_decap_8
XFILLER_9_748 VPWR VGND sg13g2_decap_8
XFILLER_40_574 VPWR VGND sg13g2_decap_8
XFILLER_8_247 VPWR VGND sg13g2_decap_8
XFILLER_5_976 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_4_442 VPWR VGND sg13g2_decap_8
XFILLER_48_630 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_36_847 VPWR VGND sg13g2_decap_8
XFILLER_39_1008 VPWR VGND sg13g2_decap_8
XFILLER_23_508 VPWR VGND sg13g2_decap_8
XFILLER_35_357 VPWR VGND sg13g2_decap_8
XFILLER_31_574 VPWR VGND sg13g2_decap_8
XFILLER_39_630 VPWR VGND sg13g2_decap_8
XFILLER_27_814 VPWR VGND sg13g2_decap_8
XFILLER_38_140 VPWR VGND sg13g2_decap_8
XFILLER_26_368 VPWR VGND sg13g2_decap_8
XFILLER_22_541 VPWR VGND sg13g2_decap_8
XFILLER_14_78 VPWR VGND sg13g2_decap_4
XFILLER_10_758 VPWR VGND sg13g2_decap_8
XFILLER_5_206 VPWR VGND sg13g2_decap_8
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_30_77 VPWR VGND sg13g2_decap_8
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_7_1006 VPWR VGND sg13g2_decap_8
XFILLER_39_42 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_18_836 VPWR VGND sg13g2_decap_8
XFILLER_29_151 VPWR VGND sg13g2_decap_8
XFILLER_45_644 VPWR VGND sg13g2_decap_8
XFILLER_17_346 VPWR VGND sg13g2_decap_8
XFILLER_44_154 VPWR VGND sg13g2_decap_8
XFILLER_41_861 VPWR VGND sg13g2_decap_8
XFILLER_13_552 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_decap_8
XFILLER_9_545 VPWR VGND sg13g2_decap_8
XFILLER_5_773 VPWR VGND sg13g2_decap_8
XFILLER_45_1001 VPWR VGND sg13g2_decap_8
XFILLER_36_644 VPWR VGND sg13g2_decap_8
XFILLER_23_305 VPWR VGND sg13g2_decap_8
XFILLER_35_154 VPWR VGND sg13g2_decap_8
XFILLER_32_861 VPWR VGND sg13g2_decap_8
XFILLER_31_371 VPWR VGND sg13g2_decap_8
XFILLER_27_611 VPWR VGND sg13g2_decap_8
XFILLER_15_806 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_27_688 VPWR VGND sg13g2_decap_8
XFILLER_14_338 VPWR VGND sg13g2_decap_8
XFILLER_26_165 VPWR VGND sg13g2_decap_8
XFILLER_42_658 VPWR VGND sg13g2_decap_8
XFILLER_25_88 VPWR VGND sg13g2_decap_8
XFILLER_23_872 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_decap_8
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_10_555 VPWR VGND sg13g2_decap_8
XFILLER_6_537 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_2_721 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_2_798 VPWR VGND sg13g2_decap_8
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_46_931 VPWR VGND sg13g2_decap_8
XFILLER_17_121 VPWR VGND sg13g2_decap_8
XFILLER_18_633 VPWR VGND sg13g2_decap_8
XFILLER_45_441 VPWR VGND sg13g2_decap_8
XFILLER_17_132 VPWR VGND sg13g2_fill_2
XFILLER_17_143 VPWR VGND sg13g2_decap_8
XFILLER_33_658 VPWR VGND sg13g2_decap_8
XFILLER_20_308 VPWR VGND sg13g2_decap_8
XFILLER_32_168 VPWR VGND sg13g2_decap_8
XFILLER_9_342 VPWR VGND sg13g2_decap_8
XFILLER_5_570 VPWR VGND sg13g2_decap_8
XFILLER_37_931 VPWR VGND sg13g2_decap_8
XFILLER_36_441 VPWR VGND sg13g2_decap_8
XFILLER_23_102 VPWR VGND sg13g2_decap_8
XFILLER_24_669 VPWR VGND sg13g2_decap_8
XFILLER_11_308 VPWR VGND sg13g2_decap_8
XFILLER_23_179 VPWR VGND sg13g2_decap_8
XFILLER_20_875 VPWR VGND sg13g2_decap_8
XFILLER_11_46 VPWR VGND sg13g2_decap_8
XFILLER_3_529 VPWR VGND sg13g2_decap_8
XFILLER_47_728 VPWR VGND sg13g2_decap_8
XFILLER_4_1009 VPWR VGND sg13g2_decap_8
XFILLER_19_419 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_28_942 VPWR VGND sg13g2_decap_8
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_15_603 VPWR VGND sg13g2_decap_8
XFILLER_43_945 VPWR VGND sg13g2_decap_8
XFILLER_27_485 VPWR VGND sg13g2_decap_8
XFILLER_42_455 VPWR VGND sg13g2_decap_8
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_35_1022 VPWR VGND sg13g2_decap_8
XFILLER_10_352 VPWR VGND sg13g2_decap_8
XFILLER_7_824 VPWR VGND sg13g2_decap_8
XFILLER_11_875 VPWR VGND sg13g2_decap_8
XFILLER_6_334 VPWR VGND sg13g2_decap_8
XFILLER_42_1015 VPWR VGND sg13g2_decap_8
XFILLER_2_595 VPWR VGND sg13g2_decap_8
X_32_ VPWR _09_ net1 VGND sg13g2_inv_1
XFILLER_38_728 VPWR VGND sg13g2_decap_8
XFILLER_37_238 VPWR VGND sg13g2_decap_8
XFILLER_18_430 VPWR VGND sg13g2_decap_8
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_34_945 VPWR VGND sg13g2_decap_8
XFILLER_33_455 VPWR VGND sg13g2_decap_8
XFILLER_20_105 VPWR VGND sg13g2_decap_8
XFILLER_29_739 VPWR VGND sg13g2_decap_8
XFILLER_28_249 VPWR VGND sg13g2_decap_8
XFILLER_25_956 VPWR VGND sg13g2_decap_8
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_24_466 VPWR VGND sg13g2_decap_8
XFILLER_12_639 VPWR VGND sg13g2_decap_8
XFILLER_40_959 VPWR VGND sg13g2_decap_8
XFILLER_20_672 VPWR VGND sg13g2_decap_8
XFILLER_22_67 VPWR VGND sg13g2_decap_4
XFILLER_4_827 VPWR VGND sg13g2_decap_8
XFILLER_3_326 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_216 VPWR VGND sg13g2_decap_8
XFILLER_15_400 VPWR VGND sg13g2_decap_8
XFILLER_16_923 VPWR VGND sg13g2_decap_8
XFILLER_43_742 VPWR VGND sg13g2_decap_8
XFILLER_27_282 VPWR VGND sg13g2_decap_8
XFILLER_42_252 VPWR VGND sg13g2_decap_8
XFILLER_15_477 VPWR VGND sg13g2_decap_8
XFILLER_31_959 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_30_469 VPWR VGND sg13g2_decap_8
XFILLER_7_621 VPWR VGND sg13g2_decap_8
XFILLER_11_672 VPWR VGND sg13g2_decap_8
XFILLER_6_131 VPWR VGND sg13g2_decap_8
XFILLER_7_698 VPWR VGND sg13g2_decap_8
XFILLER_3_893 VPWR VGND sg13g2_decap_8
XFILLER_2_392 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
XFILLER_38_525 VPWR VGND sg13g2_decap_8
XFILLER_19_783 VPWR VGND sg13g2_decap_8
XFILLER_34_742 VPWR VGND sg13g2_decap_8
XFILLER_22_926 VPWR VGND sg13g2_decap_8
XFILLER_33_252 VPWR VGND sg13g2_decap_8
XFILLER_21_458 VPWR VGND sg13g2_decap_8
XFILLER_1_819 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_29_536 VPWR VGND sg13g2_decap_8
XFILLER_44_539 VPWR VGND sg13g2_decap_8
XFILLER_17_56 VPWR VGND sg13g2_decap_8
XFILLER_25_753 VPWR VGND sg13g2_decap_8
XFILLER_24_263 VPWR VGND sg13g2_decap_8
XFILLER_12_436 VPWR VGND sg13g2_decap_8
XFILLER_13_937 VPWR VGND sg13g2_decap_8
XFILLER_33_77 VPWR VGND sg13g2_decap_8
XFILLER_40_756 VPWR VGND sg13g2_decap_8
XFILLER_8_429 VPWR VGND sg13g2_decap_8
XFILLER_4_624 VPWR VGND sg13g2_decap_8
XFILLER_3_123 VPWR VGND sg13g2_decap_8
XFILLER_48_812 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_48_889 VPWR VGND sg13g2_decap_8
XFILLER_35_539 VPWR VGND sg13g2_decap_8
XFILLER_47_399 VPWR VGND sg13g2_decap_8
XFILLER_16_720 VPWR VGND sg13g2_decap_8
XFILLER_15_274 VPWR VGND sg13g2_decap_8
XFILLER_16_797 VPWR VGND sg13g2_decap_8
XFILLER_31_756 VPWR VGND sg13g2_decap_8
XFILLER_30_266 VPWR VGND sg13g2_decap_8
XFILLER_8_996 VPWR VGND sg13g2_decap_8
XFILLER_7_495 VPWR VGND sg13g2_decap_8
XFILLER_3_690 VPWR VGND sg13g2_decap_8
XFILLER_39_812 VPWR VGND sg13g2_decap_8
XFILLER_38_322 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_889 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_19_580 VPWR VGND sg13g2_decap_8
XFILLER_38_399 VPWR VGND sg13g2_decap_8
XFILLER_22_723 VPWR VGND sg13g2_decap_8
XFILLER_21_255 VPWR VGND sg13g2_decap_8
XFILLER_1_616 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_29_333 VPWR VGND sg13g2_decap_8
XFILLER_45_826 VPWR VGND sg13g2_decap_8
XFILLER_17_528 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_25_550 VPWR VGND sg13g2_decap_8
XFILLER_13_734 VPWR VGND sg13g2_decap_8
XFILLER_44_98 VPWR VGND sg13g2_decap_8
XFILLER_9_727 VPWR VGND sg13g2_decap_8
XFILLER_12_233 VPWR VGND sg13g2_decap_8
XFILLER_40_553 VPWR VGND sg13g2_decap_8
XFILLER_8_226 VPWR VGND sg13g2_decap_8
XFILLER_5_955 VPWR VGND sg13g2_decap_8
XFILLER_4_421 VPWR VGND sg13g2_decap_8
XFILLER_4_498 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_48_686 VPWR VGND sg13g2_decap_8
XFILLER_36_826 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_35_336 VPWR VGND sg13g2_decap_8
XFILLER_16_594 VPWR VGND sg13g2_decap_8
XFILLER_31_553 VPWR VGND sg13g2_decap_8
XFILLER_8_793 VPWR VGND sg13g2_decap_8
XFILLER_7_292 VPWR VGND sg13g2_decap_8
XFILLER_22_1024 VPWR VGND sg13g2_decap_4
XFILLER_39_686 VPWR VGND sg13g2_decap_8
XFILLER_26_347 VPWR VGND sg13g2_decap_8
XFILLER_38_196 VPWR VGND sg13g2_decap_8
XFILLER_22_520 VPWR VGND sg13g2_decap_8
XFILLER_14_57 VPWR VGND sg13g2_decap_8
XFILLER_10_737 VPWR VGND sg13g2_decap_8
XFILLER_22_597 VPWR VGND sg13g2_decap_8
XFILLER_6_719 VPWR VGND sg13g2_decap_8
XFILLER_30_56 VPWR VGND sg13g2_decap_8
XFILLER_2_903 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_29_130 VPWR VGND sg13g2_decap_8
XFILLER_39_98 VPWR VGND sg13g2_decap_8
XFILLER_18_815 VPWR VGND sg13g2_decap_8
XFILLER_45_623 VPWR VGND sg13g2_decap_8
XFILLER_17_325 VPWR VGND sg13g2_decap_8
XFILLER_44_133 VPWR VGND sg13g2_decap_8
XFILLER_41_840 VPWR VGND sg13g2_decap_8
XFILLER_13_531 VPWR VGND sg13g2_decap_8
XFILLER_9_524 VPWR VGND sg13g2_decap_8
XFILLER_40_350 VPWR VGND sg13g2_decap_8
XFILLER_5_752 VPWR VGND sg13g2_decap_8
XFILLER_4_295 VPWR VGND sg13g2_decap_8
XFILLER_1_980 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_49_984 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
XFILLER_36_623 VPWR VGND sg13g2_decap_8
XFILLER_35_133 VPWR VGND sg13g2_decap_8
XFILLER_17_892 VPWR VGND sg13g2_decap_8
XFILLER_16_391 VPWR VGND sg13g2_decap_8
XFILLER_32_840 VPWR VGND sg13g2_decap_8
XFILLER_31_350 VPWR VGND sg13g2_decap_8
XFILLER_8_590 VPWR VGND sg13g2_decap_8
XFILLER_39_483 VPWR VGND sg13g2_decap_8
XFILLER_26_144 VPWR VGND sg13g2_decap_8
XFILLER_27_667 VPWR VGND sg13g2_decap_8
XFILLER_42_637 VPWR VGND sg13g2_decap_8
XFILLER_14_317 VPWR VGND sg13g2_decap_8
XFILLER_23_851 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_decap_8
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_10_534 VPWR VGND sg13g2_decap_8
XFILLER_22_394 VPWR VGND sg13g2_decap_8
XFILLER_6_516 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_2_700 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_29_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_46_910 VPWR VGND sg13g2_decap_8
XFILLER_45_420 VPWR VGND sg13g2_decap_8
XFILLER_18_612 VPWR VGND sg13g2_decap_8
XFILLER_46_987 VPWR VGND sg13g2_decap_8
XFILLER_45_497 VPWR VGND sg13g2_decap_8
XFILLER_18_689 VPWR VGND sg13g2_decap_8
XFILLER_33_637 VPWR VGND sg13g2_decap_8
XFILLER_17_199 VPWR VGND sg13g2_decap_8
XFILLER_32_147 VPWR VGND sg13g2_decap_8
XFILLER_14_884 VPWR VGND sg13g2_decap_8
XFILLER_9_321 VPWR VGND sg13g2_decap_8
XFILLER_9_398 VPWR VGND sg13g2_decap_8
XFILLER_37_910 VPWR VGND sg13g2_decap_8
XFILLER_49_781 VPWR VGND sg13g2_decap_8
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_36_420 VPWR VGND sg13g2_decap_8
XFILLER_37_987 VPWR VGND sg13g2_decap_8
XFILLER_36_497 VPWR VGND sg13g2_decap_8
XFILLER_24_648 VPWR VGND sg13g2_decap_8
XFILLER_23_158 VPWR VGND sg13g2_decap_8
XFILLER_20_854 VPWR VGND sg13g2_decap_8
XFILLER_3_508 VPWR VGND sg13g2_decap_8
XFILLER_11_25 VPWR VGND sg13g2_decap_8
XFILLER_47_707 VPWR VGND sg13g2_decap_8
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_28_921 VPWR VGND sg13g2_decap_8
XFILLER_39_280 VPWR VGND sg13g2_decap_8
XFILLER_43_924 VPWR VGND sg13g2_decap_8
XFILLER_27_464 VPWR VGND sg13g2_decap_8
XFILLER_28_998 VPWR VGND sg13g2_decap_8
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_42_434 VPWR VGND sg13g2_decap_8
XFILLER_15_659 VPWR VGND sg13g2_decap_8
XFILLER_35_1001 VPWR VGND sg13g2_decap_8
XFILLER_10_331 VPWR VGND sg13g2_decap_8
XFILLER_7_803 VPWR VGND sg13g2_decap_8
XFILLER_11_854 VPWR VGND sg13g2_decap_8
XFILLER_22_191 VPWR VGND sg13g2_decap_8
XFILLER_6_313 VPWR VGND sg13g2_decap_8
XFILLER_2_574 VPWR VGND sg13g2_decap_8
X_31_ VPWR _08_ net44 VGND sg13g2_inv_1
XFILLER_38_707 VPWR VGND sg13g2_decap_8
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_19_965 VPWR VGND sg13g2_decap_8
XFILLER_46_784 VPWR VGND sg13g2_decap_8
XFILLER_18_486 VPWR VGND sg13g2_decap_8
XFILLER_34_924 VPWR VGND sg13g2_decap_8
XFILLER_45_294 VPWR VGND sg13g2_decap_8
XFILLER_33_434 VPWR VGND sg13g2_decap_8
XFILLER_14_681 VPWR VGND sg13g2_decap_8
XFILLER_9_195 VPWR VGND sg13g2_decap_8
XFILLER_6_880 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_29_718 VPWR VGND sg13g2_decap_8
XFILLER_28_228 VPWR VGND sg13g2_decap_8
XFILLER_25_935 VPWR VGND sg13g2_decap_8
XFILLER_37_784 VPWR VGND sg13g2_decap_8
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_24_445 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
XFILLER_12_618 VPWR VGND sg13g2_decap_8
XFILLER_40_938 VPWR VGND sg13g2_decap_8
XFILLER_20_651 VPWR VGND sg13g2_decap_8
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_4_806 VPWR VGND sg13g2_decap_8
XFILLER_3_305 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
XFILLER_16_902 VPWR VGND sg13g2_decap_8
XFILLER_27_261 VPWR VGND sg13g2_decap_8
XFILLER_28_795 VPWR VGND sg13g2_decap_8
XFILLER_43_721 VPWR VGND sg13g2_decap_8
XFILLER_42_231 VPWR VGND sg13g2_decap_8
XFILLER_15_456 VPWR VGND sg13g2_decap_8
XFILLER_16_979 VPWR VGND sg13g2_decap_8
XFILLER_43_798 VPWR VGND sg13g2_decap_8
XFILLER_31_938 VPWR VGND sg13g2_decap_8
XFILLER_7_600 VPWR VGND sg13g2_decap_8
XFILLER_11_651 VPWR VGND sg13g2_decap_8
XFILLER_30_448 VPWR VGND sg13g2_decap_8
XFILLER_6_110 VPWR VGND sg13g2_decap_8
XFILLER_7_677 VPWR VGND sg13g2_decap_8
XFILLER_6_187 VPWR VGND sg13g2_decap_8
XFILLER_3_872 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
XFILLER_2_371 VPWR VGND sg13g2_decap_8
XFILLER_38_504 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_19_762 VPWR VGND sg13g2_decap_8
XFILLER_46_581 VPWR VGND sg13g2_decap_8
XFILLER_18_283 VPWR VGND sg13g2_decap_8
XFILLER_34_721 VPWR VGND sg13g2_decap_8
XFILLER_22_905 VPWR VGND sg13g2_decap_8
XFILLER_33_231 VPWR VGND sg13g2_decap_8
XFILLER_21_437 VPWR VGND sg13g2_decap_8
XFILLER_34_798 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_29_515 VPWR VGND sg13g2_decap_8
XFILLER_44_518 VPWR VGND sg13g2_decap_8
XFILLER_16_209 VPWR VGND sg13g2_decap_8
XFILLER_25_732 VPWR VGND sg13g2_decap_8
XFILLER_37_581 VPWR VGND sg13g2_decap_8
XFILLER_13_916 VPWR VGND sg13g2_decap_8
XFILLER_24_242 VPWR VGND sg13g2_decap_8
XFILLER_9_909 VPWR VGND sg13g2_decap_8
XFILLER_12_415 VPWR VGND sg13g2_decap_8
XFILLER_40_735 VPWR VGND sg13g2_decap_8
XFILLER_8_408 VPWR VGND sg13g2_decap_8
XFILLER_33_56 VPWR VGND sg13g2_decap_8
XFILLER_32_1015 VPWR VGND sg13g2_decap_8
XFILLER_4_603 VPWR VGND sg13g2_decap_8
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_48_868 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_35_518 VPWR VGND sg13g2_decap_8
XFILLER_28_592 VPWR VGND sg13g2_decap_8
XFILLER_15_253 VPWR VGND sg13g2_decap_8
XFILLER_16_776 VPWR VGND sg13g2_decap_8
XFILLER_43_595 VPWR VGND sg13g2_decap_8
XFILLER_31_735 VPWR VGND sg13g2_decap_8
XFILLER_30_245 VPWR VGND sg13g2_decap_8
XFILLER_12_982 VPWR VGND sg13g2_decap_8
XFILLER_8_975 VPWR VGND sg13g2_decap_8
XFILLER_7_474 VPWR VGND sg13g2_decap_8
XFILLER_48_1022 VPWR VGND sg13g2_decap_8
XFILLER_38_301 VPWR VGND sg13g2_decap_8
XFILLER_39_868 VPWR VGND sg13g2_decap_8
XFILLER_26_529 VPWR VGND sg13g2_decap_8
XFILLER_38_378 VPWR VGND sg13g2_decap_8
XFILLER_22_702 VPWR VGND sg13g2_decap_8
XFILLER_34_595 VPWR VGND sg13g2_decap_8
XFILLER_10_919 VPWR VGND sg13g2_decap_8
XFILLER_21_234 VPWR VGND sg13g2_decap_8
XFILLER_22_779 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_29_312 VPWR VGND sg13g2_decap_8
XFILLER_45_805 VPWR VGND sg13g2_decap_8
XFILLER_17_507 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_8
XFILLER_44_315 VPWR VGND sg13g2_decap_8
XFILLER_29_389 VPWR VGND sg13g2_decap_8
XFILLER_44_77 VPWR VGND sg13g2_decap_8
XFILLER_12_212 VPWR VGND sg13g2_decap_8
XFILLER_13_713 VPWR VGND sg13g2_decap_8
XFILLER_9_706 VPWR VGND sg13g2_decap_8
XFILLER_40_532 VPWR VGND sg13g2_decap_8
XFILLER_8_205 VPWR VGND sg13g2_decap_8
XFILLER_12_289 VPWR VGND sg13g2_decap_8
XFILLER_4_400 VPWR VGND sg13g2_decap_8
XFILLER_5_934 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_4_477 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_48_665 VPWR VGND sg13g2_decap_8
XFILLER_36_805 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
XFILLER_35_315 VPWR VGND sg13g2_decap_8
XFILLER_44_882 VPWR VGND sg13g2_decap_8
XFILLER_16_573 VPWR VGND sg13g2_decap_8
XFILLER_43_392 VPWR VGND sg13g2_decap_8
XFILLER_31_532 VPWR VGND sg13g2_decap_8
XFILLER_8_772 VPWR VGND sg13g2_decap_8
XFILLER_7_271 VPWR VGND sg13g2_decap_8
XFILLER_22_1003 VPWR VGND sg13g2_decap_8
XFILLER_39_665 VPWR VGND sg13g2_decap_8
XFILLER_26_326 VPWR VGND sg13g2_decap_8
XFILLER_27_849 VPWR VGND sg13g2_decap_8
XFILLER_38_175 VPWR VGND sg13g2_decap_8
XFILLER_42_819 VPWR VGND sg13g2_decap_8
XFILLER_35_882 VPWR VGND sg13g2_decap_8
XFILLER_41_329 VPWR VGND sg13g2_decap_8
XFILLER_34_392 VPWR VGND sg13g2_decap_8
XFILLER_10_716 VPWR VGND sg13g2_decap_8
XFILLER_22_576 VPWR VGND sg13g2_decap_8
XFILLER_30_35 VPWR VGND sg13g2_decap_8
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_77 VPWR VGND sg13g2_decap_8
XFILLER_45_602 VPWR VGND sg13g2_decap_8
XFILLER_17_304 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_29_186 VPWR VGND sg13g2_decap_8
XFILLER_45_679 VPWR VGND sg13g2_decap_8
XFILLER_33_819 VPWR VGND sg13g2_decap_8
XFILLER_44_189 VPWR VGND sg13g2_decap_8
XFILLER_13_510 VPWR VGND sg13g2_decap_8
XFILLER_26_893 VPWR VGND sg13g2_decap_8
XFILLER_32_329 VPWR VGND sg13g2_decap_8
XFILLER_9_503 VPWR VGND sg13g2_decap_8
XFILLER_41_896 VPWR VGND sg13g2_decap_8
XFILLER_13_587 VPWR VGND sg13g2_decap_8
XFILLER_5_731 VPWR VGND sg13g2_decap_8
XFILLER_4_274 VPWR VGND sg13g2_decap_8
XFILLER_49_963 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
XFILLER_36_602 VPWR VGND sg13g2_decap_8
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_36_679 VPWR VGND sg13g2_decap_8
XFILLER_17_871 VPWR VGND sg13g2_decap_8
XFILLER_35_189 VPWR VGND sg13g2_decap_8
XFILLER_16_370 VPWR VGND sg13g2_decap_8
XFILLER_32_896 VPWR VGND sg13g2_decap_8
XFILLER_39_462 VPWR VGND sg13g2_decap_8
XFILLER_26_123 VPWR VGND sg13g2_decap_8
XFILLER_27_646 VPWR VGND sg13g2_decap_8
XFILLER_42_616 VPWR VGND sg13g2_decap_8
XFILLER_23_830 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_10_513 VPWR VGND sg13g2_decap_8
XFILLER_22_373 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_2_756 VPWR VGND sg13g2_decap_8
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_46_966 VPWR VGND sg13g2_decap_8
XFILLER_18_668 VPWR VGND sg13g2_decap_8
XFILLER_45_476 VPWR VGND sg13g2_decap_8
XFILLER_17_178 VPWR VGND sg13g2_decap_8
XFILLER_33_616 VPWR VGND sg13g2_decap_8
XFILLER_26_690 VPWR VGND sg13g2_decap_8
XFILLER_32_126 VPWR VGND sg13g2_decap_8
XFILLER_9_300 VPWR VGND sg13g2_decap_8
XFILLER_14_863 VPWR VGND sg13g2_decap_8
XFILLER_41_693 VPWR VGND sg13g2_decap_8
XFILLER_13_384 VPWR VGND sg13g2_decap_8
XFILLER_9_377 VPWR VGND sg13g2_decap_8
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
XFILLER_49_4 VPWR VGND sg13g2_decap_8
XFILLER_49_760 VPWR VGND sg13g2_decap_8
XFILLER_37_966 VPWR VGND sg13g2_decap_8
XFILLER_24_627 VPWR VGND sg13g2_decap_8
XFILLER_36_476 VPWR VGND sg13g2_decap_8
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_20_833 VPWR VGND sg13g2_decap_8
XFILLER_32_693 VPWR VGND sg13g2_decap_8
XFILLER_28_900 VPWR VGND sg13g2_decap_8
XFILLER_43_903 VPWR VGND sg13g2_decap_8
XFILLER_27_443 VPWR VGND sg13g2_decap_8
XFILLER_28_977 VPWR VGND sg13g2_decap_8
XFILLER_42_413 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_14_115 VPWR VGND sg13g2_decap_4
XFILLER_15_638 VPWR VGND sg13g2_decap_8
XFILLER_10_310 VPWR VGND sg13g2_decap_8
XFILLER_11_833 VPWR VGND sg13g2_decap_8
XFILLER_22_170 VPWR VGND sg13g2_decap_8
XFILLER_7_859 VPWR VGND sg13g2_decap_8
XFILLER_10_387 VPWR VGND sg13g2_decap_8
XFILLER_6_369 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_553 VPWR VGND sg13g2_decap_8
XFILLER_19_944 VPWR VGND sg13g2_decap_8
XFILLER_46_763 VPWR VGND sg13g2_decap_8
XFILLER_18_465 VPWR VGND sg13g2_decap_8
XFILLER_34_903 VPWR VGND sg13g2_decap_8
XFILLER_45_273 VPWR VGND sg13g2_decap_8
XFILLER_33_413 VPWR VGND sg13g2_decap_8
XFILLER_21_619 VPWR VGND sg13g2_decap_8
XFILLER_42_980 VPWR VGND sg13g2_decap_8
XFILLER_14_660 VPWR VGND sg13g2_decap_8
XFILLER_41_490 VPWR VGND sg13g2_decap_8
XFILLER_13_181 VPWR VGND sg13g2_decap_8
XFILLER_9_174 VPWR VGND sg13g2_decap_8
XFILLER_3_82 VPWR VGND sg13g2_decap_8
XFILLER_28_207 VPWR VGND sg13g2_decap_8
XFILLER_25_914 VPWR VGND sg13g2_decap_8
XFILLER_37_763 VPWR VGND sg13g2_decap_8
XFILLER_24_424 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_decap_8
XFILLER_40_917 VPWR VGND sg13g2_decap_8
XFILLER_33_980 VPWR VGND sg13g2_decap_8
XFILLER_20_630 VPWR VGND sg13g2_decap_8
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_32_490 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_43_700 VPWR VGND sg13g2_decap_8
XFILLER_27_240 VPWR VGND sg13g2_decap_8
XFILLER_28_774 VPWR VGND sg13g2_decap_8
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_15_435 VPWR VGND sg13g2_decap_8
XFILLER_16_958 VPWR VGND sg13g2_decap_8
XFILLER_43_777 VPWR VGND sg13g2_decap_8
XFILLER_31_917 VPWR VGND sg13g2_decap_8
XFILLER_42_287 VPWR VGND sg13g2_decap_8
XFILLER_24_991 VPWR VGND sg13g2_decap_8
XFILLER_30_427 VPWR VGND sg13g2_decap_8
XFILLER_11_630 VPWR VGND sg13g2_decap_8
XFILLER_10_184 VPWR VGND sg13g2_decap_8
XFILLER_7_656 VPWR VGND sg13g2_decap_8
XFILLER_6_166 VPWR VGND sg13g2_decap_8
XFILLER_3_851 VPWR VGND sg13g2_decap_8
XFILLER_2_350 VPWR VGND sg13g2_decap_8
XFILLER_33_7 VPWR VGND sg13g2_decap_8
XFILLER_19_741 VPWR VGND sg13g2_decap_8
XFILLER_46_560 VPWR VGND sg13g2_decap_8
XFILLER_34_700 VPWR VGND sg13g2_decap_8
XFILLER_18_262 VPWR VGND sg13g2_decap_8
XFILLER_33_210 VPWR VGND sg13g2_decap_8
XFILLER_34_777 VPWR VGND sg13g2_decap_8
XFILLER_21_416 VPWR VGND sg13g2_decap_8
XFILLER_33_287 VPWR VGND sg13g2_decap_8
XFILLER_30_994 VPWR VGND sg13g2_decap_8
XFILLER_25_1012 VPWR VGND sg13g2_decap_8
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_37_560 VPWR VGND sg13g2_decap_8
XFILLER_25_711 VPWR VGND sg13g2_decap_8
XFILLER_24_221 VPWR VGND sg13g2_decap_8
XFILLER_25_788 VPWR VGND sg13g2_decap_8
XFILLER_40_714 VPWR VGND sg13g2_decap_8
XFILLER_24_298 VPWR VGND sg13g2_decap_8
XFILLER_33_35 VPWR VGND sg13g2_decap_8
XFILLER_21_983 VPWR VGND sg13g2_decap_8
XFILLER_4_659 VPWR VGND sg13g2_decap_8
XFILLER_3_158 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_48_847 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_28_571 VPWR VGND sg13g2_decap_8
XFILLER_15_232 VPWR VGND sg13g2_decap_8
XFILLER_16_755 VPWR VGND sg13g2_decap_8
XFILLER_43_574 VPWR VGND sg13g2_decap_8
XFILLER_31_714 VPWR VGND sg13g2_decap_8
XFILLER_30_224 VPWR VGND sg13g2_decap_8
XFILLER_12_961 VPWR VGND sg13g2_decap_8
XFILLER_8_954 VPWR VGND sg13g2_decap_8
XFILLER_7_453 VPWR VGND sg13g2_decap_8
XFILLER_48_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_847 VPWR VGND sg13g2_decap_8
XFILLER_26_508 VPWR VGND sg13g2_decap_8
XFILLER_38_357 VPWR VGND sg13g2_decap_8
XFILLER_34_574 VPWR VGND sg13g2_decap_8
XFILLER_21_213 VPWR VGND sg13g2_decap_8
XFILLER_22_758 VPWR VGND sg13g2_decap_8
XFILLER_9_92 VPWR VGND sg13g2_decap_8
XFILLER_30_791 VPWR VGND sg13g2_decap_8
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_29_368 VPWR VGND sg13g2_decap_8
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_25_585 VPWR VGND sg13g2_decap_8
XFILLER_40_511 VPWR VGND sg13g2_decap_8
XFILLER_13_769 VPWR VGND sg13g2_decap_8
XFILLER_12_268 VPWR VGND sg13g2_decap_8
XFILLER_40_588 VPWR VGND sg13g2_decap_8
XFILLER_21_780 VPWR VGND sg13g2_decap_8
XFILLER_5_913 VPWR VGND sg13g2_decap_8
XFILLER_4_456 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_644 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_44_861 VPWR VGND sg13g2_decap_8
XFILLER_16_552 VPWR VGND sg13g2_decap_8
XFILLER_43_371 VPWR VGND sg13g2_decap_8
XFILLER_31_511 VPWR VGND sg13g2_decap_8
XFILLER_31_588 VPWR VGND sg13g2_decap_8
XFILLER_8_751 VPWR VGND sg13g2_decap_8
XFILLER_7_250 VPWR VGND sg13g2_decap_8
XFILLER_39_644 VPWR VGND sg13g2_decap_8
XFILLER_27_828 VPWR VGND sg13g2_decap_8
XFILLER_38_154 VPWR VGND sg13g2_decap_8
XFILLER_26_305 VPWR VGND sg13g2_decap_8
XFILLER_35_861 VPWR VGND sg13g2_decap_8
XFILLER_41_308 VPWR VGND sg13g2_decap_8
XFILLER_14_15 VPWR VGND sg13g2_fill_2
XFILLER_34_371 VPWR VGND sg13g2_decap_8
XFILLER_22_555 VPWR VGND sg13g2_decap_8
XFILLER_30_14 VPWR VGND sg13g2_decap_8
XFILLER_2_938 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_39_56 VPWR VGND sg13g2_decap_8
XFILLER_29_165 VPWR VGND sg13g2_decap_8
XFILLER_45_658 VPWR VGND sg13g2_decap_8
XFILLER_44_168 VPWR VGND sg13g2_decap_8
XFILLER_26_872 VPWR VGND sg13g2_decap_8
XFILLER_32_308 VPWR VGND sg13g2_decap_8
XFILLER_38_1022 VPWR VGND sg13g2_decap_8
XFILLER_25_382 VPWR VGND sg13g2_decap_8
XFILLER_41_875 VPWR VGND sg13g2_decap_8
XFILLER_13_566 VPWR VGND sg13g2_decap_8
XFILLER_9_559 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_5_710 VPWR VGND sg13g2_decap_8
XFILLER_5_787 VPWR VGND sg13g2_decap_8
XFILLER_4_253 VPWR VGND sg13g2_decap_8
XFILLER_45_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_91 VPWR VGND sg13g2_decap_8
XFILLER_49_942 VPWR VGND sg13g2_decap_8
XFILLER_48_441 VPWR VGND sg13g2_decap_8
XFILLER_17_850 VPWR VGND sg13g2_decap_8
XFILLER_24_809 VPWR VGND sg13g2_decap_8
XFILLER_36_658 VPWR VGND sg13g2_decap_8
XFILLER_23_319 VPWR VGND sg13g2_decap_8
XFILLER_35_168 VPWR VGND sg13g2_decap_8
XFILLER_32_875 VPWR VGND sg13g2_decap_8
XFILLER_31_385 VPWR VGND sg13g2_decap_8
XFILLER_6_82 VPWR VGND sg13g2_decap_8
XFILLER_6_1020 VPWR VGND sg13g2_decap_8
XFILLER_39_441 VPWR VGND sg13g2_decap_8
XFILLER_26_102 VPWR VGND sg13g2_decap_8
XFILLER_27_625 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_26_179 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
XFILLER_22_352 VPWR VGND sg13g2_decap_8
XFILLER_23_886 VPWR VGND sg13g2_decap_8
XFILLER_10_569 VPWR VGND sg13g2_decap_8
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_735 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_fill_2
XFILLER_2_29 VPWR VGND sg13g2_fill_2
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_46_945 VPWR VGND sg13g2_decap_8
XFILLER_45_455 VPWR VGND sg13g2_decap_8
XFILLER_18_647 VPWR VGND sg13g2_decap_8
XFILLER_17_157 VPWR VGND sg13g2_decap_8
XFILLER_32_105 VPWR VGND sg13g2_decap_8
XFILLER_14_842 VPWR VGND sg13g2_decap_8
XFILLER_41_672 VPWR VGND sg13g2_decap_8
XFILLER_13_363 VPWR VGND sg13g2_decap_8
XFILLER_9_356 VPWR VGND sg13g2_decap_8
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
XFILLER_5_584 VPWR VGND sg13g2_decap_8
XFILLER_37_945 VPWR VGND sg13g2_decap_8
XFILLER_24_606 VPWR VGND sg13g2_decap_8
XFILLER_36_455 VPWR VGND sg13g2_decap_8
XFILLER_23_116 VPWR VGND sg13g2_decap_8
XFILLER_20_812 VPWR VGND sg13g2_decap_8
XFILLER_32_672 VPWR VGND sg13g2_decap_8
XFILLER_31_182 VPWR VGND sg13g2_decap_8
XFILLER_20_889 VPWR VGND sg13g2_decap_8
XFILLER_27_422 VPWR VGND sg13g2_decap_8
XFILLER_28_956 VPWR VGND sg13g2_decap_8
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_15_617 VPWR VGND sg13g2_decap_8
XFILLER_43_959 VPWR VGND sg13g2_decap_8
XFILLER_27_499 VPWR VGND sg13g2_decap_8
XFILLER_42_469 VPWR VGND sg13g2_decap_8
XFILLER_14_149 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_decap_8
XFILLER_11_812 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_decap_8
XFILLER_10_366 VPWR VGND sg13g2_decap_8
XFILLER_7_838 VPWR VGND sg13g2_decap_8
XFILLER_11_889 VPWR VGND sg13g2_decap_8
XFILLER_6_348 VPWR VGND sg13g2_decap_8
XFILLER_2_532 VPWR VGND sg13g2_decap_8
XFILLER_19_923 VPWR VGND sg13g2_decap_8
XFILLER_46_742 VPWR VGND sg13g2_decap_8
XFILLER_18_444 VPWR VGND sg13g2_decap_8
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_34_959 VPWR VGND sg13g2_decap_8
XFILLER_33_469 VPWR VGND sg13g2_decap_8
XFILLER_20_119 VPWR VGND sg13g2_decap_8
XFILLER_9_153 VPWR VGND sg13g2_decap_8
XFILLER_5_381 VPWR VGND sg13g2_decap_8
XFILLER_3_61 VPWR VGND sg13g2_decap_8
XFILLER_3_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_742 VPWR VGND sg13g2_decap_8
XFILLER_24_403 VPWR VGND sg13g2_decap_8
XFILLER_36_252 VPWR VGND sg13g2_decap_8
XFILLER_20_686 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_28_753 VPWR VGND sg13g2_decap_8
XFILLER_15_414 VPWR VGND sg13g2_decap_8
XFILLER_16_937 VPWR VGND sg13g2_decap_8
XFILLER_27_296 VPWR VGND sg13g2_decap_8
XFILLER_43_756 VPWR VGND sg13g2_decap_8
XFILLER_42_266 VPWR VGND sg13g2_decap_8
XFILLER_24_970 VPWR VGND sg13g2_decap_8
XFILLER_30_406 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
XFILLER_23_480 VPWR VGND sg13g2_decap_8
XFILLER_10_163 VPWR VGND sg13g2_decap_8
XFILLER_7_635 VPWR VGND sg13g2_decap_8
XFILLER_11_686 VPWR VGND sg13g2_decap_8
XFILLER_6_145 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
XFILLER_3_830 VPWR VGND sg13g2_decap_8
XFILLER_19_720 VPWR VGND sg13g2_decap_8
XFILLER_38_539 VPWR VGND sg13g2_decap_8
XFILLER_18_241 VPWR VGND sg13g2_decap_8
XFILLER_19_797 VPWR VGND sg13g2_decap_8
XFILLER_34_756 VPWR VGND sg13g2_decap_8
XFILLER_15_981 VPWR VGND sg13g2_decap_8
XFILLER_33_266 VPWR VGND sg13g2_decap_8
XFILLER_30_973 VPWR VGND sg13g2_decap_8
XFILLER_24_200 VPWR VGND sg13g2_decap_8
XFILLER_25_767 VPWR VGND sg13g2_decap_8
XFILLER_24_277 VPWR VGND sg13g2_decap_8
XFILLER_33_14 VPWR VGND sg13g2_decap_8
XFILLER_21_962 VPWR VGND sg13g2_decap_8
XFILLER_20_483 VPWR VGND sg13g2_decap_8
XFILLER_4_638 VPWR VGND sg13g2_decap_8
XFILLER_3_137 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_48_826 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_28_550 VPWR VGND sg13g2_decap_8
XFILLER_15_211 VPWR VGND sg13g2_decap_8
XFILLER_16_734 VPWR VGND sg13g2_decap_8
XFILLER_43_553 VPWR VGND sg13g2_decap_8
XFILLER_30_203 VPWR VGND sg13g2_decap_8
XFILLER_12_940 VPWR VGND sg13g2_decap_8
XFILLER_15_288 VPWR VGND sg13g2_decap_8
XFILLER_8_933 VPWR VGND sg13g2_decap_8
XFILLER_7_432 VPWR VGND sg13g2_decap_8
XFILLER_11_483 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_39_826 VPWR VGND sg13g2_decap_8
XFILLER_38_336 VPWR VGND sg13g2_decap_8
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_19_594 VPWR VGND sg13g2_decap_8
XFILLER_34_553 VPWR VGND sg13g2_decap_8
XFILLER_22_737 VPWR VGND sg13g2_decap_8
XFILLER_9_60 VPWR VGND sg13g2_decap_8
XFILLER_21_269 VPWR VGND sg13g2_decap_8
XFILLER_30_770 VPWR VGND sg13g2_decap_8
XFILLER_28_25 VPWR VGND sg13g2_decap_8
XFILLER_29_347 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_25_564 VPWR VGND sg13g2_decap_8
XFILLER_13_748 VPWR VGND sg13g2_decap_8
XFILLER_12_247 VPWR VGND sg13g2_decap_8
XFILLER_40_567 VPWR VGND sg13g2_decap_8
XFILLER_20_280 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_fill_2
XFILLER_5_969 VPWR VGND sg13g2_decap_8
XFILLER_4_435 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_623 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_44_840 VPWR VGND sg13g2_decap_8
XFILLER_16_531 VPWR VGND sg13g2_decap_8
XFILLER_43_350 VPWR VGND sg13g2_decap_8
XFILLER_31_567 VPWR VGND sg13g2_decap_8
XFILLER_8_730 VPWR VGND sg13g2_decap_8
XFILLER_15_1023 VPWR VGND sg13g2_decap_4
XFILLER_11_280 VPWR VGND sg13g2_decap_8
XFILLER_39_623 VPWR VGND sg13g2_decap_8
XFILLER_27_807 VPWR VGND sg13g2_decap_8
XFILLER_38_133 VPWR VGND sg13g2_decap_8
XFILLER_19_391 VPWR VGND sg13g2_decap_8
XFILLER_35_840 VPWR VGND sg13g2_decap_8
XFILLER_34_350 VPWR VGND sg13g2_decap_8
XFILLER_22_534 VPWR VGND sg13g2_decap_8
XFILLER_2_917 VPWR VGND sg13g2_decap_8
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_39_35 VPWR VGND sg13g2_decap_8
XFILLER_29_144 VPWR VGND sg13g2_decap_8
XFILLER_45_637 VPWR VGND sg13g2_decap_8
XFILLER_18_829 VPWR VGND sg13g2_decap_8
XFILLER_44_147 VPWR VGND sg13g2_decap_8
XFILLER_17_339 VPWR VGND sg13g2_decap_8
XFILLER_26_851 VPWR VGND sg13g2_decap_8
XFILLER_25_361 VPWR VGND sg13g2_decap_8
XFILLER_38_1001 VPWR VGND sg13g2_decap_8
XFILLER_41_854 VPWR VGND sg13g2_decap_8
XFILLER_13_545 VPWR VGND sg13g2_decap_8
XFILLER_9_538 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_5_766 VPWR VGND sg13g2_decap_8
XFILLER_4_232 VPWR VGND sg13g2_decap_8
XFILLER_49_921 VPWR VGND sg13g2_decap_8
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_1_994 VPWR VGND sg13g2_decap_8
XFILLER_49_998 VPWR VGND sg13g2_decap_8
XFILLER_36_637 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_35_147 VPWR VGND sg13g2_decap_8
XFILLER_32_854 VPWR VGND sg13g2_decap_8
XFILLER_31_364 VPWR VGND sg13g2_decap_8
XFILLER_6_61 VPWR VGND sg13g2_decap_8
XFILLER_39_420 VPWR VGND sg13g2_decap_8
XFILLER_27_604 VPWR VGND sg13g2_decap_8
XFILLER_39_497 VPWR VGND sg13g2_decap_8
XFILLER_26_158 VPWR VGND sg13g2_decap_8
XFILLER_22_331 VPWR VGND sg13g2_decap_8
XFILLER_23_865 VPWR VGND sg13g2_decap_8
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_10_548 VPWR VGND sg13g2_decap_8
XFILLER_2_714 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_46_924 VPWR VGND sg13g2_decap_8
XFILLER_18_626 VPWR VGND sg13g2_decap_8
XFILLER_45_434 VPWR VGND sg13g2_decap_8
XFILLER_17_114 VPWR VGND sg13g2_decap_8
XFILLER_14_821 VPWR VGND sg13g2_decap_8
XFILLER_41_651 VPWR VGND sg13g2_decap_8
XFILLER_13_342 VPWR VGND sg13g2_decap_8
XFILLER_14_898 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_decap_8
XFILLER_40_161 VPWR VGND sg13g2_decap_8
XFILLER_9_335 VPWR VGND sg13g2_decap_8
XFILLER_5_563 VPWR VGND sg13g2_decap_8
XFILLER_31_91 VPWR VGND sg13g2_decap_8
XFILLER_1_791 VPWR VGND sg13g2_decap_8
XFILLER_49_795 VPWR VGND sg13g2_decap_8
XFILLER_37_924 VPWR VGND sg13g2_decap_8
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_36_434 VPWR VGND sg13g2_decap_8
XFILLER_32_651 VPWR VGND sg13g2_decap_8
XFILLER_31_161 VPWR VGND sg13g2_decap_8
XFILLER_20_868 VPWR VGND sg13g2_decap_8
XFILLER_11_39 VPWR VGND sg13g2_decap_8
XFILLER_27_401 VPWR VGND sg13g2_decap_8
XFILLER_28_935 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_27_478 VPWR VGND sg13g2_decap_8
XFILLER_43_938 VPWR VGND sg13g2_decap_8
XFILLER_14_128 VPWR VGND sg13g2_decap_4
XFILLER_42_448 VPWR VGND sg13g2_decap_8
XFILLER_23_662 VPWR VGND sg13g2_decap_8
XFILLER_35_1015 VPWR VGND sg13g2_decap_8
XFILLER_10_345 VPWR VGND sg13g2_decap_8
XFILLER_7_817 VPWR VGND sg13g2_decap_8
XFILLER_11_868 VPWR VGND sg13g2_decap_8
XFILLER_6_327 VPWR VGND sg13g2_decap_8
XFILLER_2_511 VPWR VGND sg13g2_decap_8
XFILLER_42_1008 VPWR VGND sg13g2_decap_8
XFILLER_2_588 VPWR VGND sg13g2_decap_8
XFILLER_19_902 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_decap_8
XFILLER_18_423 VPWR VGND sg13g2_decap_8
XFILLER_45_231 VPWR VGND sg13g2_decap_8
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_46_798 VPWR VGND sg13g2_decap_8
XFILLER_34_938 VPWR VGND sg13g2_decap_8
XFILLER_33_448 VPWR VGND sg13g2_decap_8
XFILLER_9_132 VPWR VGND sg13g2_decap_8
XFILLER_14_695 VPWR VGND sg13g2_decap_8
X_58__19 VPWR VGND net sg13g2_tiehi
XFILLER_6_894 VPWR VGND sg13g2_decap_8
XFILLER_5_360 VPWR VGND sg13g2_decap_8
XFILLER_3_40 VPWR VGND sg13g2_decap_8
XFILLER_49_592 VPWR VGND sg13g2_decap_8
XFILLER_37_721 VPWR VGND sg13g2_decap_8
XFILLER_36_231 VPWR VGND sg13g2_decap_8
XFILLER_18_990 VPWR VGND sg13g2_decap_8
XFILLER_25_949 VPWR VGND sg13g2_decap_8
XFILLER_37_798 VPWR VGND sg13g2_decap_8
XFILLER_24_459 VPWR VGND sg13g2_decap_8
XFILLER_20_665 VPWR VGND sg13g2_decap_8
XFILLER_3_319 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_19_209 VPWR VGND sg13g2_decap_8
XFILLER_28_732 VPWR VGND sg13g2_decap_8
XFILLER_16_916 VPWR VGND sg13g2_decap_8
XFILLER_43_735 VPWR VGND sg13g2_decap_8
XFILLER_27_275 VPWR VGND sg13g2_decap_8
XFILLER_42_245 VPWR VGND sg13g2_decap_8
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_10_142 VPWR VGND sg13g2_decap_8
XFILLER_7_614 VPWR VGND sg13g2_decap_8
XFILLER_11_665 VPWR VGND sg13g2_decap_8
XFILLER_6_124 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_decap_8
XFILLER_3_886 VPWR VGND sg13g2_decap_8
XFILLER_2_385 VPWR VGND sg13g2_decap_8
XFILLER_38_518 VPWR VGND sg13g2_decap_8
XFILLER_18_220 VPWR VGND sg13g2_decap_8
XFILLER_19_776 VPWR VGND sg13g2_decap_8
XFILLER_46_595 VPWR VGND sg13g2_decap_8
XFILLER_34_735 VPWR VGND sg13g2_decap_8
XFILLER_18_297 VPWR VGND sg13g2_decap_8
XFILLER_33_245 VPWR VGND sg13g2_decap_8
XFILLER_15_960 VPWR VGND sg13g2_decap_8
XFILLER_22_919 VPWR VGND sg13g2_decap_8
XFILLER_14_492 VPWR VGND sg13g2_decap_8
XFILLER_30_952 VPWR VGND sg13g2_decap_8
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_6_691 VPWR VGND sg13g2_decap_8
XFILLER_29_529 VPWR VGND sg13g2_decap_8
XFILLER_17_49 VPWR VGND sg13g2_decap_8
XFILLER_25_746 VPWR VGND sg13g2_decap_8
XFILLER_37_595 VPWR VGND sg13g2_decap_8
XFILLER_24_256 VPWR VGND sg13g2_decap_8
XFILLER_12_429 VPWR VGND sg13g2_decap_8
XFILLER_21_941 VPWR VGND sg13g2_decap_8
XFILLER_40_749 VPWR VGND sg13g2_decap_8
XFILLER_20_462 VPWR VGND sg13g2_decap_8
XFILLER_4_617 VPWR VGND sg13g2_decap_8
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_48_805 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_16_713 VPWR VGND sg13g2_decap_8
XFILLER_43_532 VPWR VGND sg13g2_decap_8
XFILLER_15_267 VPWR VGND sg13g2_decap_8
XFILLER_31_749 VPWR VGND sg13g2_decap_8
XFILLER_8_912 VPWR VGND sg13g2_decap_8
XFILLER_30_259 VPWR VGND sg13g2_decap_8
XFILLER_7_411 VPWR VGND sg13g2_decap_8
XFILLER_11_462 VPWR VGND sg13g2_decap_8
XFILLER_12_996 VPWR VGND sg13g2_decap_8
XFILLER_23_81 VPWR VGND sg13g2_decap_8
XFILLER_8_989 VPWR VGND sg13g2_decap_8
XFILLER_7_488 VPWR VGND sg13g2_decap_8
XFILLER_3_683 VPWR VGND sg13g2_decap_8
XFILLER_2_182 VPWR VGND sg13g2_decap_8
XFILLER_39_805 VPWR VGND sg13g2_decap_8
XFILLER_38_315 VPWR VGND sg13g2_decap_8
XFILLER_47_882 VPWR VGND sg13g2_decap_8
XFILLER_19_573 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_34_532 VPWR VGND sg13g2_decap_8
XFILLER_22_716 VPWR VGND sg13g2_decap_8
XFILLER_21_248 VPWR VGND sg13g2_decap_8
XFILLER_1_609 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_29_326 VPWR VGND sg13g2_decap_8
XFILLER_45_819 VPWR VGND sg13g2_decap_8
XFILLER_44_329 VPWR VGND sg13g2_decap_8
XFILLER_38_882 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_25_543 VPWR VGND sg13g2_decap_8
XFILLER_37_392 VPWR VGND sg13g2_decap_8
XFILLER_12_226 VPWR VGND sg13g2_decap_8
XFILLER_13_727 VPWR VGND sg13g2_decap_8
XFILLER_40_546 VPWR VGND sg13g2_decap_8
XFILLER_8_219 VPWR VGND sg13g2_decap_8
XFILLER_5_948 VPWR VGND sg13g2_decap_8
XFILLER_4_414 VPWR VGND sg13g2_decap_8
XFILLER_48_602 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_48_679 VPWR VGND sg13g2_decap_8
XFILLER_36_819 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_35_329 VPWR VGND sg13g2_decap_8
XFILLER_16_510 VPWR VGND sg13g2_decap_8
XFILLER_18_81 VPWR VGND sg13g2_decap_8
XFILLER_29_893 VPWR VGND sg13g2_decap_8
XFILLER_44_896 VPWR VGND sg13g2_decap_8
XFILLER_16_587 VPWR VGND sg13g2_decap_8
XFILLER_15_1002 VPWR VGND sg13g2_decap_8
XFILLER_31_546 VPWR VGND sg13g2_decap_8
XFILLER_34_91 VPWR VGND sg13g2_decap_8
XFILLER_12_793 VPWR VGND sg13g2_decap_8
XFILLER_8_786 VPWR VGND sg13g2_decap_8
XFILLER_7_285 VPWR VGND sg13g2_decap_8
XFILLER_4_981 VPWR VGND sg13g2_decap_8
XFILLER_3_480 VPWR VGND sg13g2_decap_8
XFILLER_39_602 VPWR VGND sg13g2_decap_8
XFILLER_38_112 VPWR VGND sg13g2_decap_8
XFILLER_22_1017 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_679 VPWR VGND sg13g2_decap_8
XFILLER_19_370 VPWR VGND sg13g2_decap_8
XFILLER_38_189 VPWR VGND sg13g2_decap_8
XFILLER_22_513 VPWR VGND sg13g2_decap_8
XFILLER_35_896 VPWR VGND sg13g2_decap_8
XFILLER_30_49 VPWR VGND sg13g2_decap_8
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_18_808 VPWR VGND sg13g2_decap_8
XFILLER_29_123 VPWR VGND sg13g2_decap_8
XFILLER_45_616 VPWR VGND sg13g2_decap_8
XFILLER_17_318 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_26_830 VPWR VGND sg13g2_decap_8
XFILLER_25_340 VPWR VGND sg13g2_decap_8
XFILLER_41_833 VPWR VGND sg13g2_decap_8
XFILLER_13_524 VPWR VGND sg13g2_decap_8
XFILLER_9_517 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_5_745 VPWR VGND sg13g2_decap_8
XFILLER_4_211 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_4_288 VPWR VGND sg13g2_decap_8
XFILLER_49_900 VPWR VGND sg13g2_decap_8
XFILLER_1_973 VPWR VGND sg13g2_decap_8
XFILLER_49_977 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_36_616 VPWR VGND sg13g2_decap_8
XFILLER_29_690 VPWR VGND sg13g2_decap_8
XFILLER_35_126 VPWR VGND sg13g2_decap_8
XFILLER_44_693 VPWR VGND sg13g2_decap_8
XFILLER_16_384 VPWR VGND sg13g2_decap_8
XFILLER_17_885 VPWR VGND sg13g2_decap_8
XFILLER_32_833 VPWR VGND sg13g2_decap_8
XFILLER_31_343 VPWR VGND sg13g2_decap_8
XFILLER_12_590 VPWR VGND sg13g2_decap_8
XFILLER_8_583 VPWR VGND sg13g2_decap_8
XFILLER_39_476 VPWR VGND sg13g2_decap_8
XFILLER_26_137 VPWR VGND sg13g2_decap_8
XFILLER_22_310 VPWR VGND sg13g2_decap_8
XFILLER_35_693 VPWR VGND sg13g2_decap_8
XFILLER_23_844 VPWR VGND sg13g2_decap_8
XFILLER_10_527 VPWR VGND sg13g2_decap_8
XFILLER_6_509 VPWR VGND sg13g2_decap_8
XFILLER_22_387 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_46_903 VPWR VGND sg13g2_decap_8
XFILLER_18_605 VPWR VGND sg13g2_decap_8
XFILLER_45_413 VPWR VGND sg13g2_decap_8
XFILLER_14_800 VPWR VGND sg13g2_decap_8
XFILLER_41_630 VPWR VGND sg13g2_decap_8
XFILLER_13_321 VPWR VGND sg13g2_decap_8
XFILLER_9_314 VPWR VGND sg13g2_decap_8
XFILLER_14_877 VPWR VGND sg13g2_decap_8
XFILLER_15_60 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_13_398 VPWR VGND sg13g2_decap_8
XFILLER_31_70 VPWR VGND sg13g2_decap_8
XFILLER_5_542 VPWR VGND sg13g2_decap_8
XFILLER_1_770 VPWR VGND sg13g2_decap_8
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_49_774 VPWR VGND sg13g2_decap_8
XFILLER_37_903 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_36_413 VPWR VGND sg13g2_decap_8
XFILLER_45_980 VPWR VGND sg13g2_decap_8
XFILLER_17_682 VPWR VGND sg13g2_decap_8
XFILLER_44_490 VPWR VGND sg13g2_decap_8
XFILLER_16_181 VPWR VGND sg13g2_decap_8
XFILLER_32_630 VPWR VGND sg13g2_decap_8
XFILLER_31_140 VPWR VGND sg13g2_decap_8
XFILLER_20_847 VPWR VGND sg13g2_decap_8
XFILLER_9_881 VPWR VGND sg13g2_decap_8
XFILLER_8_380 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_fill_2
XFILLER_28_1012 VPWR VGND sg13g2_decap_8
XFILLER_28_914 VPWR VGND sg13g2_decap_8
XFILLER_39_273 VPWR VGND sg13g2_decap_8
XFILLER_43_917 VPWR VGND sg13g2_decap_8
XFILLER_27_457 VPWR VGND sg13g2_decap_8
XFILLER_42_427 VPWR VGND sg13g2_decap_8
XFILLER_36_980 VPWR VGND sg13g2_decap_8
XFILLER_23_641 VPWR VGND sg13g2_decap_8
XFILLER_35_490 VPWR VGND sg13g2_decap_8
XFILLER_10_324 VPWR VGND sg13g2_decap_8
XFILLER_11_847 VPWR VGND sg13g2_decap_8
XFILLER_22_184 VPWR VGND sg13g2_decap_8
XFILLER_6_306 VPWR VGND sg13g2_decap_8
XFILLER_2_567 VPWR VGND sg13g2_decap_8
XFILLER_46_700 VPWR VGND sg13g2_decap_8
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_18_402 VPWR VGND sg13g2_decap_8
XFILLER_19_958 VPWR VGND sg13g2_decap_8
XFILLER_46_777 VPWR VGND sg13g2_decap_8
XFILLER_34_917 VPWR VGND sg13g2_decap_8
XFILLER_45_287 VPWR VGND sg13g2_decap_8
XFILLER_18_479 VPWR VGND sg13g2_decap_8
XFILLER_33_427 VPWR VGND sg13g2_decap_8
XFILLER_26_81 VPWR VGND sg13g2_decap_8
XFILLER_14_674 VPWR VGND sg13g2_decap_8
XFILLER_42_994 VPWR VGND sg13g2_decap_8
XFILLER_9_111 VPWR VGND sg13g2_fill_1
XFILLER_13_195 VPWR VGND sg13g2_decap_8
XFILLER_42_91 VPWR VGND sg13g2_decap_8
XFILLER_9_188 VPWR VGND sg13g2_decap_8
XFILLER_6_873 VPWR VGND sg13g2_decap_8
XFILLER_10_891 VPWR VGND sg13g2_decap_8
XFILLER_37_700 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_decap_8
XFILLER_36_210 VPWR VGND sg13g2_decap_8
XFILLER_37_777 VPWR VGND sg13g2_decap_8
XFILLER_25_928 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_8
XFILLER_24_438 VPWR VGND sg13g2_decap_8
XFILLER_33_994 VPWR VGND sg13g2_decap_8
XFILLER_20_644 VPWR VGND sg13g2_decap_8
XFILLER_22_39 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_711 VPWR VGND sg13g2_decap_8
XFILLER_43_714 VPWR VGND sg13g2_decap_8
XFILLER_27_254 VPWR VGND sg13g2_decap_8
XFILLER_28_788 VPWR VGND sg13g2_decap_8
XFILLER_42_224 VPWR VGND sg13g2_decap_8
XFILLER_15_449 VPWR VGND sg13g2_decap_8
XFILLER_10_121 VPWR VGND sg13g2_decap_8
XFILLER_11_644 VPWR VGND sg13g2_decap_8
XFILLER_6_103 VPWR VGND sg13g2_decap_8
XFILLER_10_198 VPWR VGND sg13g2_decap_8
XFILLER_3_865 VPWR VGND sg13g2_decap_8
XFILLER_2_364 VPWR VGND sg13g2_decap_8
XFILLER_19_755 VPWR VGND sg13g2_decap_8
XFILLER_46_574 VPWR VGND sg13g2_decap_8
XFILLER_18_276 VPWR VGND sg13g2_decap_8
XFILLER_34_714 VPWR VGND sg13g2_decap_8
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_33_224 VPWR VGND sg13g2_decap_8
XFILLER_18_1011 VPWR VGND sg13g2_decap_8
XFILLER_42_791 VPWR VGND sg13g2_decap_8
XFILLER_14_471 VPWR VGND sg13g2_decap_8
XFILLER_30_931 VPWR VGND sg13g2_decap_8
XFILLER_6_670 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_8
XFILLER_25_1026 VPWR VGND sg13g2_fill_2
XFILLER_29_508 VPWR VGND sg13g2_decap_8
XFILLER_25_725 VPWR VGND sg13g2_decap_8
XFILLER_37_574 VPWR VGND sg13g2_decap_8
XFILLER_13_909 VPWR VGND sg13g2_decap_8
XFILLER_24_235 VPWR VGND sg13g2_decap_8
XFILLER_12_408 VPWR VGND sg13g2_decap_8
XFILLER_40_728 VPWR VGND sg13g2_decap_8
XFILLER_21_920 VPWR VGND sg13g2_decap_8
XFILLER_33_49 VPWR VGND sg13g2_decap_8
XFILLER_33_791 VPWR VGND sg13g2_decap_8
XFILLER_20_441 VPWR VGND sg13g2_decap_8
XFILLER_32_1008 VPWR VGND sg13g2_decap_8
XFILLER_21_997 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_43_511 VPWR VGND sg13g2_decap_8
XFILLER_28_585 VPWR VGND sg13g2_decap_8
XFILLER_15_246 VPWR VGND sg13g2_decap_8
XFILLER_16_769 VPWR VGND sg13g2_decap_8
XFILLER_43_588 VPWR VGND sg13g2_decap_8
XFILLER_31_728 VPWR VGND sg13g2_decap_8
XFILLER_11_441 VPWR VGND sg13g2_decap_8
XFILLER_30_238 VPWR VGND sg13g2_decap_8
XFILLER_12_975 VPWR VGND sg13g2_decap_8
XFILLER_23_60 VPWR VGND sg13g2_decap_8
XFILLER_8_968 VPWR VGND sg13g2_decap_8
XFILLER_7_467 VPWR VGND sg13g2_decap_8
XFILLER_48_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_662 VPWR VGND sg13g2_decap_8
XFILLER_2_161 VPWR VGND sg13g2_decap_8
XFILLER_31_7 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_552 VPWR VGND sg13g2_decap_8
XFILLER_46_371 VPWR VGND sg13g2_decap_8
XFILLER_34_511 VPWR VGND sg13g2_decap_8
XFILLER_21_227 VPWR VGND sg13g2_decap_8
XFILLER_34_588 VPWR VGND sg13g2_decap_8
XFILLER_29_305 VPWR VGND sg13g2_decap_8
XFILLER_44_308 VPWR VGND sg13g2_decap_8
XFILLER_38_861 VPWR VGND sg13g2_decap_8
XFILLER_25_522 VPWR VGND sg13g2_decap_8
XFILLER_37_371 VPWR VGND sg13g2_decap_8
XFILLER_13_706 VPWR VGND sg13g2_decap_8
XFILLER_12_205 VPWR VGND sg13g2_decap_8
XFILLER_25_599 VPWR VGND sg13g2_decap_8
XFILLER_40_525 VPWR VGND sg13g2_decap_8
XFILLER_21_794 VPWR VGND sg13g2_decap_8
XFILLER_5_927 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_48_658 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_29_872 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_decap_8
XFILLER_28_382 VPWR VGND sg13g2_decap_8
XFILLER_44_875 VPWR VGND sg13g2_decap_8
XFILLER_16_566 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_31_525 VPWR VGND sg13g2_decap_8
XFILLER_34_70 VPWR VGND sg13g2_decap_8
XFILLER_12_772 VPWR VGND sg13g2_decap_8
XFILLER_8_765 VPWR VGND sg13g2_decap_8
XFILLER_7_264 VPWR VGND sg13g2_decap_8
XFILLER_4_960 VPWR VGND sg13g2_decap_8
XFILLER_39_658 VPWR VGND sg13g2_decap_8
XFILLER_26_319 VPWR VGND sg13g2_decap_8
XFILLER_38_168 VPWR VGND sg13g2_decap_8
XFILLER_35_875 VPWR VGND sg13g2_decap_8
XFILLER_34_385 VPWR VGND sg13g2_decap_8
XFILLER_10_709 VPWR VGND sg13g2_decap_8
XFILLER_22_569 VPWR VGND sg13g2_decap_8
XFILLER_30_28 VPWR VGND sg13g2_decap_8
XFILLER_29_102 VPWR VGND sg13g2_decap_8
XFILLER_29_179 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_41_812 VPWR VGND sg13g2_decap_8
XFILLER_13_503 VPWR VGND sg13g2_decap_8
XFILLER_26_886 VPWR VGND sg13g2_decap_8
XFILLER_25_396 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_decap_8
XFILLER_41_889 VPWR VGND sg13g2_decap_8
XFILLER_21_591 VPWR VGND sg13g2_decap_8
XFILLER_40_399 VPWR VGND sg13g2_decap_8
XFILLER_5_724 VPWR VGND sg13g2_decap_8
XFILLER_4_267 VPWR VGND sg13g2_decap_8
XFILLER_1_952 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_49_956 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_29_81 VPWR VGND sg13g2_decap_8
XFILLER_35_105 VPWR VGND sg13g2_decap_8
XFILLER_17_864 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XFILLER_44_672 VPWR VGND sg13g2_decap_8
XFILLER_16_363 VPWR VGND sg13g2_decap_8
XFILLER_32_812 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_decap_8
XFILLER_31_322 VPWR VGND sg13g2_decap_8
XFILLER_32_889 VPWR VGND sg13g2_decap_8
XFILLER_31_399 VPWR VGND sg13g2_decap_8
XFILLER_8_562 VPWR VGND sg13g2_decap_8
XFILLER_6_96 VPWR VGND sg13g2_decap_8
XFILLER_39_455 VPWR VGND sg13g2_decap_8
XFILLER_26_116 VPWR VGND sg13g2_decap_8
XFILLER_27_639 VPWR VGND sg13g2_decap_8
XFILLER_42_609 VPWR VGND sg13g2_decap_8
XFILLER_23_823 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_35_672 VPWR VGND sg13g2_decap_8
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_34_182 VPWR VGND sg13g2_decap_8
XFILLER_10_506 VPWR VGND sg13g2_decap_8
XFILLER_22_366 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_2_749 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_46_959 VPWR VGND sg13g2_decap_8
XFILLER_17_105 VPWR VGND sg13g2_decap_4
XFILLER_45_469 VPWR VGND sg13g2_decap_8
XFILLER_33_609 VPWR VGND sg13g2_decap_8
XFILLER_13_300 VPWR VGND sg13g2_decap_8
XFILLER_26_683 VPWR VGND sg13g2_decap_8
XFILLER_32_119 VPWR VGND sg13g2_decap_8
XFILLER_14_856 VPWR VGND sg13g2_decap_8
XFILLER_25_193 VPWR VGND sg13g2_decap_8
XFILLER_41_686 VPWR VGND sg13g2_decap_8
XFILLER_13_377 VPWR VGND sg13g2_decap_8
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_5_521 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_598 VPWR VGND sg13g2_decap_8
Xoutput3 net3 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_49_753 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_37_959 VPWR VGND sg13g2_decap_8
XFILLER_36_469 VPWR VGND sg13g2_decap_8
XFILLER_16_160 VPWR VGND sg13g2_decap_8
XFILLER_17_661 VPWR VGND sg13g2_decap_8
XFILLER_20_826 VPWR VGND sg13g2_decap_8
XFILLER_32_686 VPWR VGND sg13g2_decap_8
XFILLER_9_860 VPWR VGND sg13g2_decap_8
XFILLER_31_196 VPWR VGND sg13g2_decap_8
XFILLER_39_252 VPWR VGND sg13g2_decap_8
XFILLER_27_436 VPWR VGND sg13g2_decap_8
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_decap_8
XFILLER_14_108 VPWR VGND sg13g2_decap_8
XFILLER_23_620 VPWR VGND sg13g2_decap_8
XFILLER_10_303 VPWR VGND sg13g2_decap_8
XFILLER_11_826 VPWR VGND sg13g2_decap_8
XFILLER_22_163 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_decap_8
XFILLER_2_546 VPWR VGND sg13g2_decap_8
XFILLER_19_937 VPWR VGND sg13g2_decap_8
XFILLER_46_756 VPWR VGND sg13g2_decap_8
XFILLER_18_458 VPWR VGND sg13g2_decap_8
XFILLER_45_266 VPWR VGND sg13g2_decap_8
XFILLER_26_60 VPWR VGND sg13g2_decap_8
XFILLER_33_406 VPWR VGND sg13g2_decap_8
XFILLER_26_480 VPWR VGND sg13g2_decap_8
XFILLER_42_973 VPWR VGND sg13g2_decap_8
XFILLER_14_653 VPWR VGND sg13g2_decap_8
XFILLER_41_483 VPWR VGND sg13g2_decap_8
XFILLER_9_101 VPWR VGND sg13g2_fill_1
XFILLER_13_174 VPWR VGND sg13g2_decap_8
XFILLER_42_70 VPWR VGND sg13g2_decap_8
XFILLER_9_167 VPWR VGND sg13g2_decap_8
XFILLER_10_870 VPWR VGND sg13g2_decap_8
XFILLER_6_852 VPWR VGND sg13g2_decap_8
XFILLER_5_395 VPWR VGND sg13g2_decap_8
XFILLER_49_550 VPWR VGND sg13g2_decap_8
XFILLER_3_75 VPWR VGND sg13g2_decap_8
XFILLER_3_1026 VPWR VGND sg13g2_fill_2
XFILLER_25_907 VPWR VGND sg13g2_decap_8
XFILLER_37_756 VPWR VGND sg13g2_decap_8
XFILLER_24_417 VPWR VGND sg13g2_decap_8
XFILLER_36_266 VPWR VGND sg13g2_decap_8
XFILLER_33_973 VPWR VGND sg13g2_decap_8
XFILLER_20_623 VPWR VGND sg13g2_decap_8
XFILLER_32_483 VPWR VGND sg13g2_decap_8
XFILLER_22_18 VPWR VGND sg13g2_decap_8
X_57__21 VPWR VGND net20 sg13g2_tiehi
XFILLER_27_233 VPWR VGND sg13g2_decap_8
XFILLER_28_767 VPWR VGND sg13g2_decap_8
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_15_428 VPWR VGND sg13g2_decap_8
XFILLER_10_100 VPWR VGND sg13g2_decap_8
XFILLER_11_623 VPWR VGND sg13g2_decap_8
XFILLER_24_984 VPWR VGND sg13g2_decap_8
XFILLER_23_494 VPWR VGND sg13g2_decap_8
XFILLER_10_177 VPWR VGND sg13g2_decap_8
XFILLER_7_649 VPWR VGND sg13g2_decap_8
XFILLER_6_159 VPWR VGND sg13g2_decap_8
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_3_844 VPWR VGND sg13g2_decap_8
XFILLER_2_343 VPWR VGND sg13g2_decap_8
XFILLER_19_734 VPWR VGND sg13g2_decap_8
XFILLER_46_553 VPWR VGND sg13g2_decap_8
XFILLER_18_255 VPWR VGND sg13g2_decap_8
XFILLER_33_203 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_14_450 VPWR VGND sg13g2_decap_8
XFILLER_21_409 VPWR VGND sg13g2_decap_8
XFILLER_42_770 VPWR VGND sg13g2_decap_8
XFILLER_15_995 VPWR VGND sg13g2_decap_8
XFILLER_30_910 VPWR VGND sg13g2_decap_8
XFILLER_41_280 VPWR VGND sg13g2_decap_8
XFILLER_30_987 VPWR VGND sg13g2_decap_8
XFILLER_5_192 VPWR VGND sg13g2_decap_8
XFILLER_25_1005 VPWR VGND sg13g2_decap_8
XFILLER_25_704 VPWR VGND sg13g2_decap_8
XFILLER_37_553 VPWR VGND sg13g2_decap_8
XFILLER_24_214 VPWR VGND sg13g2_decap_8
XFILLER_40_707 VPWR VGND sg13g2_decap_8
XFILLER_33_28 VPWR VGND sg13g2_decap_8
XFILLER_33_770 VPWR VGND sg13g2_decap_8
XFILLER_20_420 VPWR VGND sg13g2_decap_8
XFILLER_32_280 VPWR VGND sg13g2_decap_8
XFILLER_21_976 VPWR VGND sg13g2_decap_8
XFILLER_20_497 VPWR VGND sg13g2_decap_8
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_28_564 VPWR VGND sg13g2_decap_8
XFILLER_15_225 VPWR VGND sg13g2_decap_8
XFILLER_16_748 VPWR VGND sg13g2_decap_8
XFILLER_43_567 VPWR VGND sg13g2_decap_8
XFILLER_31_707 VPWR VGND sg13g2_decap_8
XFILLER_24_781 VPWR VGND sg13g2_decap_8
XFILLER_30_217 VPWR VGND sg13g2_decap_8
XFILLER_11_420 VPWR VGND sg13g2_decap_8
XFILLER_12_954 VPWR VGND sg13g2_decap_8
XFILLER_23_291 VPWR VGND sg13g2_decap_8
XFILLER_8_947 VPWR VGND sg13g2_decap_8
XFILLER_7_446 VPWR VGND sg13g2_decap_8
XFILLER_11_497 VPWR VGND sg13g2_decap_8
XFILLER_3_641 VPWR VGND sg13g2_decap_8
XFILLER_2_140 VPWR VGND sg13g2_decap_8
XFILLER_47_840 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_19_531 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_34_567 VPWR VGND sg13g2_decap_8
XFILLER_21_206 VPWR VGND sg13g2_decap_8
XFILLER_15_792 VPWR VGND sg13g2_decap_8
XFILLER_9_74 VPWR VGND sg13g2_decap_8
XFILLER_30_784 VPWR VGND sg13g2_decap_8
XFILLER_9_1021 VPWR VGND sg13g2_decap_8
XFILLER_28_39 VPWR VGND sg13g2_decap_8
XFILLER_38_840 VPWR VGND sg13g2_decap_8
XFILLER_25_501 VPWR VGND sg13g2_decap_8
XFILLER_37_350 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_25_578 VPWR VGND sg13g2_decap_8
XFILLER_40_504 VPWR VGND sg13g2_decap_8
XFILLER_21_773 VPWR VGND sg13g2_decap_8
XFILLER_5_906 VPWR VGND sg13g2_decap_8
XFILLER_20_294 VPWR VGND sg13g2_decap_8
XFILLER_4_449 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_48_637 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_29_851 VPWR VGND sg13g2_decap_8
XFILLER_28_361 VPWR VGND sg13g2_decap_8
XFILLER_44_854 VPWR VGND sg13g2_decap_8
XFILLER_16_545 VPWR VGND sg13g2_decap_8
XFILLER_43_364 VPWR VGND sg13g2_decap_8
XFILLER_31_504 VPWR VGND sg13g2_decap_8
XFILLER_12_751 VPWR VGND sg13g2_decap_8
XFILLER_8_744 VPWR VGND sg13g2_decap_8
XFILLER_7_243 VPWR VGND sg13g2_decap_8
XFILLER_11_294 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_39_637 VPWR VGND sg13g2_decap_8
XFILLER_38_147 VPWR VGND sg13g2_decap_8
XFILLER_35_854 VPWR VGND sg13g2_decap_8
XFILLER_34_364 VPWR VGND sg13g2_decap_8
XFILLER_22_548 VPWR VGND sg13g2_decap_8
XFILLER_30_581 VPWR VGND sg13g2_decap_8
XFILLER_39_49 VPWR VGND sg13g2_decap_8
XFILLER_29_158 VPWR VGND sg13g2_decap_8
XFILLER_26_865 VPWR VGND sg13g2_decap_8
XFILLER_25_375 VPWR VGND sg13g2_decap_8
XFILLER_38_1015 VPWR VGND sg13g2_decap_8
XFILLER_40_301 VPWR VGND sg13g2_decap_8
XFILLER_41_868 VPWR VGND sg13g2_decap_8
XFILLER_13_559 VPWR VGND sg13g2_decap_8
XFILLER_40_378 VPWR VGND sg13g2_decap_8
XFILLER_21_570 VPWR VGND sg13g2_decap_8
XFILLER_5_703 VPWR VGND sg13g2_decap_8
XFILLER_4_246 VPWR VGND sg13g2_decap_8
XFILLER_45_1008 VPWR VGND sg13g2_decap_8
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_49_935 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_29_60 VPWR VGND sg13g2_decap_8
XFILLER_44_651 VPWR VGND sg13g2_decap_8
XFILLER_16_342 VPWR VGND sg13g2_decap_8
XFILLER_17_843 VPWR VGND sg13g2_decap_8
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_31_301 VPWR VGND sg13g2_decap_8
XFILLER_32_868 VPWR VGND sg13g2_decap_8
XFILLER_31_378 VPWR VGND sg13g2_decap_8
XFILLER_8_541 VPWR VGND sg13g2_decap_8
XFILLER_6_75 VPWR VGND sg13g2_decap_8
XFILLER_6_1013 VPWR VGND sg13g2_decap_8
XFILLER_39_434 VPWR VGND sg13g2_decap_8
XFILLER_27_618 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_35_651 VPWR VGND sg13g2_decap_8
XFILLER_23_802 VPWR VGND sg13g2_decap_8
XFILLER_34_161 VPWR VGND sg13g2_decap_8
XFILLER_22_345 VPWR VGND sg13g2_decap_8
XFILLER_23_879 VPWR VGND sg13g2_decap_8
XFILLER_41_28 VPWR VGND sg13g2_decap_8
XFILLER_2_728 VPWR VGND sg13g2_decap_8
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_46_938 VPWR VGND sg13g2_decap_8
XFILLER_45_448 VPWR VGND sg13g2_decap_8
XFILLER_17_128 VPWR VGND sg13g2_decap_4
XFILLER_26_662 VPWR VGND sg13g2_decap_8
XFILLER_14_835 VPWR VGND sg13g2_decap_8
XFILLER_25_172 VPWR VGND sg13g2_decap_8
XFILLER_41_665 VPWR VGND sg13g2_decap_8
XFILLER_13_356 VPWR VGND sg13g2_decap_8
XFILLER_9_349 VPWR VGND sg13g2_decap_8
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_5_500 VPWR VGND sg13g2_decap_8
XFILLER_5_577 VPWR VGND sg13g2_decap_8
Xoutput4 net4 uio_out[1] VPWR VGND sg13g2_buf_1
XFILLER_49_732 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_37_938 VPWR VGND sg13g2_decap_8
XFILLER_17_640 VPWR VGND sg13g2_decap_8
XFILLER_36_448 VPWR VGND sg13g2_decap_8
XFILLER_23_109 VPWR VGND sg13g2_decap_8
XFILLER_20_805 VPWR VGND sg13g2_decap_8
XFILLER_32_665 VPWR VGND sg13g2_decap_8
XFILLER_31_175 VPWR VGND sg13g2_decap_8
XFILLER_39_231 VPWR VGND sg13g2_decap_8
XFILLER_27_415 VPWR VGND sg13g2_decap_8
XFILLER_28_949 VPWR VGND sg13g2_decap_8
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_11_805 VPWR VGND sg13g2_decap_8
XFILLER_22_142 VPWR VGND sg13g2_decap_8
XFILLER_23_676 VPWR VGND sg13g2_decap_8
XFILLER_10_359 VPWR VGND sg13g2_decap_8
XFILLER_2_525 VPWR VGND sg13g2_decap_8
XFILLER_19_916 VPWR VGND sg13g2_decap_8
XFILLER_46_735 VPWR VGND sg13g2_decap_8
XFILLER_45_245 VPWR VGND sg13g2_decap_8
XFILLER_18_437 VPWR VGND sg13g2_decap_8
XFILLER_27_982 VPWR VGND sg13g2_decap_8
XFILLER_14_632 VPWR VGND sg13g2_decap_8
XFILLER_42_952 VPWR VGND sg13g2_decap_8
XFILLER_13_120 VPWR VGND sg13g2_decap_8
XFILLER_41_462 VPWR VGND sg13g2_decap_8
XFILLER_9_146 VPWR VGND sg13g2_decap_8
XFILLER_6_831 VPWR VGND sg13g2_decap_8
XFILLER_5_374 VPWR VGND sg13g2_decap_8
XFILLER_3_54 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_4
XFILLER_3_1005 VPWR VGND sg13g2_decap_8
X_85_ net10 net18 VPWR VGND sg13g2_buf_1
XFILLER_37_735 VPWR VGND sg13g2_decap_8
XFILLER_36_245 VPWR VGND sg13g2_decap_8
XFILLER_33_952 VPWR VGND sg13g2_decap_8
XFILLER_20_602 VPWR VGND sg13g2_decap_8
XFILLER_32_462 VPWR VGND sg13g2_decap_8
XFILLER_20_679 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_41_1022 VPWR VGND sg13g2_decap_8
XFILLER_27_212 VPWR VGND sg13g2_decap_8
XFILLER_28_746 VPWR VGND sg13g2_decap_8
XFILLER_15_407 VPWR VGND sg13g2_decap_8
XFILLER_43_749 VPWR VGND sg13g2_decap_8
XFILLER_27_289 VPWR VGND sg13g2_decap_8
XFILLER_42_259 VPWR VGND sg13g2_decap_8
XFILLER_24_963 VPWR VGND sg13g2_decap_8
XFILLER_11_602 VPWR VGND sg13g2_decap_8
XFILLER_23_473 VPWR VGND sg13g2_decap_8
XFILLER_10_156 VPWR VGND sg13g2_decap_8
XFILLER_7_628 VPWR VGND sg13g2_decap_8
XFILLER_11_679 VPWR VGND sg13g2_decap_8
XFILLER_6_138 VPWR VGND sg13g2_decap_8
XFILLER_12_74 VPWR VGND sg13g2_decap_8
XFILLER_3_823 VPWR VGND sg13g2_decap_8
XFILLER_2_322 VPWR VGND sg13g2_decap_8
XFILLER_2_399 VPWR VGND sg13g2_decap_8
XFILLER_19_713 VPWR VGND sg13g2_decap_8
XFILLER_46_532 VPWR VGND sg13g2_decap_8
XFILLER_18_234 VPWR VGND sg13g2_decap_8
XFILLER_34_749 VPWR VGND sg13g2_decap_8
XFILLER_33_259 VPWR VGND sg13g2_decap_8
XFILLER_15_974 VPWR VGND sg13g2_decap_8
XFILLER_30_966 VPWR VGND sg13g2_decap_8
XFILLER_5_171 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_532 VPWR VGND sg13g2_decap_8
XFILLER_21_955 VPWR VGND sg13g2_decap_8
XFILLER_20_476 VPWR VGND sg13g2_decap_8
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_48_819 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_28_543 VPWR VGND sg13g2_decap_8
XFILLER_15_204 VPWR VGND sg13g2_decap_8
XFILLER_16_727 VPWR VGND sg13g2_decap_8
XFILLER_43_546 VPWR VGND sg13g2_decap_8
XFILLER_24_760 VPWR VGND sg13g2_decap_8
XFILLER_12_933 VPWR VGND sg13g2_decap_8
XFILLER_23_270 VPWR VGND sg13g2_decap_8
XFILLER_8_926 VPWR VGND sg13g2_decap_8
XFILLER_7_425 VPWR VGND sg13g2_decap_8
XFILLER_11_476 VPWR VGND sg13g2_decap_8
XFILLER_23_95 VPWR VGND sg13g2_decap_8
XFILLER_3_620 VPWR VGND sg13g2_decap_8
XFILLER_3_697 VPWR VGND sg13g2_decap_8
XFILLER_2_196 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_39_819 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_19_510 VPWR VGND sg13g2_decap_8
XFILLER_38_329 VPWR VGND sg13g2_decap_8
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_896 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_19_587 VPWR VGND sg13g2_decap_8
XFILLER_34_546 VPWR VGND sg13g2_decap_8
XFILLER_9_20 VPWR VGND sg13g2_fill_1
XFILLER_15_771 VPWR VGND sg13g2_decap_8
XFILLER_9_53 VPWR VGND sg13g2_decap_8
XFILLER_30_763 VPWR VGND sg13g2_decap_8
XFILLER_7_992 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_9_1000 VPWR VGND sg13g2_decap_8
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_38_896 VPWR VGND sg13g2_decap_8
XFILLER_44_28 VPWR VGND sg13g2_decap_8
XFILLER_25_557 VPWR VGND sg13g2_decap_8
XFILLER_21_752 VPWR VGND sg13g2_decap_8
XFILLER_20_273 VPWR VGND sg13g2_decap_8
XFILLER_4_428 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_48_616 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_29_830 VPWR VGND sg13g2_decap_8
XFILLER_28_340 VPWR VGND sg13g2_decap_8
XFILLER_44_833 VPWR VGND sg13g2_decap_8
XFILLER_16_524 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_12_730 VPWR VGND sg13g2_decap_8
XFILLER_15_1016 VPWR VGND sg13g2_decap_8
XFILLER_15_1027 VPWR VGND sg13g2_fill_2
XFILLER_8_723 VPWR VGND sg13g2_decap_8
XFILLER_7_222 VPWR VGND sg13g2_decap_8
XFILLER_11_273 VPWR VGND sg13g2_decap_8
XFILLER_7_299 VPWR VGND sg13g2_decap_8
XFILLER_4_995 VPWR VGND sg13g2_decap_8
XFILLER_3_494 VPWR VGND sg13g2_decap_8
XFILLER_39_616 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_38_126 VPWR VGND sg13g2_decap_8
XFILLER_47_693 VPWR VGND sg13g2_decap_8
XFILLER_19_384 VPWR VGND sg13g2_decap_8
XFILLER_35_833 VPWR VGND sg13g2_decap_8
XFILLER_34_343 VPWR VGND sg13g2_decap_8
XFILLER_22_527 VPWR VGND sg13g2_decap_8
XFILLER_30_560 VPWR VGND sg13g2_decap_8
XFILLER_39_28 VPWR VGND sg13g2_decap_8
XFILLER_29_137 VPWR VGND sg13g2_decap_8
XFILLER_26_844 VPWR VGND sg13g2_decap_8
XFILLER_38_693 VPWR VGND sg13g2_decap_8
XFILLER_25_354 VPWR VGND sg13g2_decap_8
XFILLER_41_847 VPWR VGND sg13g2_decap_8
XFILLER_13_538 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_5_759 VPWR VGND sg13g2_decap_8
XFILLER_4_225 VPWR VGND sg13g2_decap_8
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_49_914 VPWR VGND sg13g2_decap_8
XFILLER_1_987 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_17_822 VPWR VGND sg13g2_decap_8
XFILLER_44_630 VPWR VGND sg13g2_decap_8
XFILLER_16_321 VPWR VGND sg13g2_decap_8
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_17_899 VPWR VGND sg13g2_decap_8
XFILLER_16_398 VPWR VGND sg13g2_decap_8
XFILLER_32_847 VPWR VGND sg13g2_decap_8
XFILLER_31_357 VPWR VGND sg13g2_decap_8
XFILLER_8_520 VPWR VGND sg13g2_decap_8
XFILLER_8_597 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_decap_4
XFILLER_6_54 VPWR VGND sg13g2_decap_8
XFILLER_4_792 VPWR VGND sg13g2_decap_8
XFILLER_3_291 VPWR VGND sg13g2_decap_8
XFILLER_39_413 VPWR VGND sg13g2_decap_8
XFILLER_48_980 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
XFILLER_19_181 VPWR VGND sg13g2_decap_8
XFILLER_35_630 VPWR VGND sg13g2_decap_8
XFILLER_34_140 VPWR VGND sg13g2_decap_8
XFILLER_22_324 VPWR VGND sg13g2_decap_8
XFILLER_23_858 VPWR VGND sg13g2_decap_8
XFILLER_2_707 VPWR VGND sg13g2_decap_8
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_46_917 VPWR VGND sg13g2_decap_8
Xheichips25_template_30 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_45_427 VPWR VGND sg13g2_decap_8
XFILLER_18_619 VPWR VGND sg13g2_decap_8
XFILLER_39_980 VPWR VGND sg13g2_decap_8
XFILLER_26_641 VPWR VGND sg13g2_decap_8
XFILLER_38_490 VPWR VGND sg13g2_decap_8
XFILLER_14_814 VPWR VGND sg13g2_decap_8
XFILLER_25_151 VPWR VGND sg13g2_decap_8
XFILLER_41_644 VPWR VGND sg13g2_decap_8
XFILLER_13_335 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_9_328 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_8
XFILLER_22_891 VPWR VGND sg13g2_decap_8
XFILLER_5_556 VPWR VGND sg13g2_decap_8
XFILLER_31_84 VPWR VGND sg13g2_decap_8
Xoutput5 net5 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_49_711 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_decap_8
XFILLER_49_788 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_36_427 VPWR VGND sg13g2_decap_8
XFILLER_45_994 VPWR VGND sg13g2_decap_8
XFILLER_17_696 VPWR VGND sg13g2_decap_8
XFILLER_16_195 VPWR VGND sg13g2_decap_8
XFILLER_32_644 VPWR VGND sg13g2_decap_8
XFILLER_31_154 VPWR VGND sg13g2_decap_8
XFILLER_9_895 VPWR VGND sg13g2_decap_8
XFILLER_8_394 VPWR VGND sg13g2_decap_8
XFILLER_28_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_210 VPWR VGND sg13g2_decap_8
XFILLER_28_928 VPWR VGND sg13g2_decap_8
XFILLER_39_287 VPWR VGND sg13g2_decap_8
XFILLER_36_994 VPWR VGND sg13g2_decap_8
XFILLER_22_121 VPWR VGND sg13g2_decap_8
XFILLER_23_655 VPWR VGND sg13g2_decap_8
XFILLER_35_1008 VPWR VGND sg13g2_decap_8
XFILLER_10_338 VPWR VGND sg13g2_decap_8
XFILLER_22_198 VPWR VGND sg13g2_decap_8
XFILLER_2_504 VPWR VGND sg13g2_decap_8
XFILLER_46_714 VPWR VGND sg13g2_decap_8
XFILLER_18_416 VPWR VGND sg13g2_decap_8
XFILLER_45_224 VPWR VGND sg13g2_decap_8
XFILLER_27_961 VPWR VGND sg13g2_decap_8
XFILLER_42_931 VPWR VGND sg13g2_decap_8
XFILLER_14_611 VPWR VGND sg13g2_decap_8
XFILLER_41_441 VPWR VGND sg13g2_decap_8
XFILLER_26_95 VPWR VGND sg13g2_decap_8
XFILLER_9_125 VPWR VGND sg13g2_decap_8
XFILLER_14_688 VPWR VGND sg13g2_decap_8
XFILLER_6_810 VPWR VGND sg13g2_decap_8
XFILLER_6_887 VPWR VGND sg13g2_decap_8
XFILLER_5_353 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_49_585 VPWR VGND sg13g2_decap_8
X_84_ net9 net17 VPWR VGND sg13g2_buf_1
XFILLER_37_714 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_36_224 VPWR VGND sg13g2_decap_8
XFILLER_45_791 VPWR VGND sg13g2_decap_8
XFILLER_18_983 VPWR VGND sg13g2_decap_8
XFILLER_33_931 VPWR VGND sg13g2_decap_8
XFILLER_17_493 VPWR VGND sg13g2_decap_8
XFILLER_32_441 VPWR VGND sg13g2_decap_8
XFILLER_20_658 VPWR VGND sg13g2_decap_8
XFILLER_9_692 VPWR VGND sg13g2_decap_8
XFILLER_8_191 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_41_1001 VPWR VGND sg13g2_decap_8
XFILLER_28_725 VPWR VGND sg13g2_decap_8
XFILLER_16_909 VPWR VGND sg13g2_decap_8
XFILLER_27_268 VPWR VGND sg13g2_decap_8
XFILLER_43_728 VPWR VGND sg13g2_decap_8
XFILLER_36_791 VPWR VGND sg13g2_decap_8
XFILLER_42_238 VPWR VGND sg13g2_decap_8
XFILLER_24_942 VPWR VGND sg13g2_decap_8
XFILLER_23_452 VPWR VGND sg13g2_decap_8
XFILLER_7_607 VPWR VGND sg13g2_decap_8
XFILLER_11_658 VPWR VGND sg13g2_decap_8
XFILLER_10_135 VPWR VGND sg13g2_decap_8
XFILLER_6_117 VPWR VGND sg13g2_decap_8
XFILLER_12_53 VPWR VGND sg13g2_decap_8
XFILLER_3_802 VPWR VGND sg13g2_decap_8
XFILLER_2_301 VPWR VGND sg13g2_decap_8
XFILLER_3_879 VPWR VGND sg13g2_decap_8
XFILLER_2_378 VPWR VGND sg13g2_decap_8
XFILLER_46_511 VPWR VGND sg13g2_decap_8
XFILLER_18_213 VPWR VGND sg13g2_decap_8
XFILLER_19_769 VPWR VGND sg13g2_decap_8
XFILLER_46_588 VPWR VGND sg13g2_decap_8
XFILLER_34_728 VPWR VGND sg13g2_decap_8
XFILLER_15_953 VPWR VGND sg13g2_decap_8
XFILLER_33_238 VPWR VGND sg13g2_decap_8
XFILLER_18_1025 VPWR VGND sg13g2_decap_4
XFILLER_14_485 VPWR VGND sg13g2_decap_8
XFILLER_30_945 VPWR VGND sg13g2_decap_8
X_54__26 VPWR VGND net25 sg13g2_tiehi
XFILLER_6_684 VPWR VGND sg13g2_decap_8
XFILLER_5_150 VPWR VGND sg13g2_decap_8
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_37_511 VPWR VGND sg13g2_decap_8
XFILLER_18_780 VPWR VGND sg13g2_decap_8
XFILLER_25_739 VPWR VGND sg13g2_decap_8
XFILLER_37_588 VPWR VGND sg13g2_decap_8
XFILLER_17_290 VPWR VGND sg13g2_decap_8
XFILLER_24_249 VPWR VGND sg13g2_decap_8
XFILLER_21_934 VPWR VGND sg13g2_decap_8
XFILLER_20_455 VPWR VGND sg13g2_decap_8
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_28_522 VPWR VGND sg13g2_decap_8
XFILLER_16_706 VPWR VGND sg13g2_decap_8
XFILLER_43_525 VPWR VGND sg13g2_decap_8
XFILLER_28_599 VPWR VGND sg13g2_decap_8
XFILLER_12_912 VPWR VGND sg13g2_decap_8
XFILLER_8_905 VPWR VGND sg13g2_decap_8
XFILLER_7_404 VPWR VGND sg13g2_decap_8
XFILLER_11_455 VPWR VGND sg13g2_decap_8
XFILLER_12_989 VPWR VGND sg13g2_decap_8
XFILLER_23_74 VPWR VGND sg13g2_decap_8
XFILLER_3_676 VPWR VGND sg13g2_decap_8
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_38_308 VPWR VGND sg13g2_decap_8
XFILLER_47_875 VPWR VGND sg13g2_decap_8
XFILLER_19_566 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_34_525 VPWR VGND sg13g2_decap_8
XFILLER_22_709 VPWR VGND sg13g2_decap_8
XFILLER_15_750 VPWR VGND sg13g2_decap_8
XFILLER_9_32 VPWR VGND sg13g2_decap_8
XFILLER_14_282 VPWR VGND sg13g2_decap_8
XFILLER_30_742 VPWR VGND sg13g2_decap_8
XFILLER_31_1022 VPWR VGND sg13g2_decap_8
XFILLER_7_971 VPWR VGND sg13g2_decap_8
XFILLER_6_481 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_29_319 VPWR VGND sg13g2_decap_8
XFILLER_38_875 VPWR VGND sg13g2_decap_8
XFILLER_37_385 VPWR VGND sg13g2_decap_8
XFILLER_25_536 VPWR VGND sg13g2_decap_8
XFILLER_12_219 VPWR VGND sg13g2_decap_8
XFILLER_21_731 VPWR VGND sg13g2_decap_8
XFILLER_40_539 VPWR VGND sg13g2_decap_8
XFILLER_20_252 VPWR VGND sg13g2_decap_8
XFILLER_4_407 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_44_812 VPWR VGND sg13g2_decap_8
XFILLER_16_503 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_29_886 VPWR VGND sg13g2_decap_8
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_28_396 VPWR VGND sg13g2_decap_8
XFILLER_44_889 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_31_539 VPWR VGND sg13g2_decap_8
XFILLER_8_702 VPWR VGND sg13g2_decap_8
XFILLER_34_84 VPWR VGND sg13g2_decap_8
XFILLER_7_201 VPWR VGND sg13g2_decap_8
XFILLER_11_252 VPWR VGND sg13g2_decap_8
XFILLER_12_786 VPWR VGND sg13g2_decap_8
XFILLER_8_779 VPWR VGND sg13g2_decap_8
XFILLER_7_278 VPWR VGND sg13g2_decap_8
XFILLER_4_974 VPWR VGND sg13g2_decap_8
XFILLER_3_473 VPWR VGND sg13g2_decap_8
XFILLER_38_105 VPWR VGND sg13g2_decap_8
XFILLER_47_672 VPWR VGND sg13g2_decap_8
XFILLER_19_363 VPWR VGND sg13g2_decap_8
XFILLER_35_812 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
XFILLER_34_322 VPWR VGND sg13g2_decap_8
XFILLER_22_506 VPWR VGND sg13g2_decap_8
XFILLER_35_889 VPWR VGND sg13g2_decap_8
XFILLER_34_399 VPWR VGND sg13g2_decap_8
XFILLER_29_116 VPWR VGND sg13g2_decap_8
XFILLER_45_609 VPWR VGND sg13g2_decap_8
XFILLER_44_119 VPWR VGND sg13g2_decap_8
XFILLER_26_823 VPWR VGND sg13g2_decap_8
XFILLER_38_672 VPWR VGND sg13g2_decap_8
XFILLER_25_333 VPWR VGND sg13g2_decap_8
XFILLER_37_182 VPWR VGND sg13g2_decap_8
XFILLER_13_517 VPWR VGND sg13g2_decap_8
XFILLER_41_826 VPWR VGND sg13g2_decap_8
XFILLER_40_336 VPWR VGND sg13g2_decap_8
XFILLER_5_738 VPWR VGND sg13g2_decap_8
XFILLER_4_204 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_1_966 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
Xhold40 _01_ VPWR VGND net40 sg13g2_dlygate4sd3_1
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_29_95 VPWR VGND sg13g2_decap_8
XFILLER_36_609 VPWR VGND sg13g2_decap_8
XFILLER_17_801 VPWR VGND sg13g2_decap_8
XFILLER_29_683 VPWR VGND sg13g2_decap_8
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_16_300 VPWR VGND sg13g2_decap_8
XFILLER_28_193 VPWR VGND sg13g2_decap_8
XFILLER_17_878 VPWR VGND sg13g2_decap_8
XFILLER_44_686 VPWR VGND sg13g2_decap_8
XFILLER_16_377 VPWR VGND sg13g2_decap_8
XFILLER_32_826 VPWR VGND sg13g2_decap_8
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_31_336 VPWR VGND sg13g2_decap_8
XFILLER_12_583 VPWR VGND sg13g2_decap_8
XFILLER_8_576 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_4_771 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_decap_8
XFILLER_39_469 VPWR VGND sg13g2_decap_8
XFILLER_19_160 VPWR VGND sg13g2_decap_8
XFILLER_22_303 VPWR VGND sg13g2_decap_8
XFILLER_23_837 VPWR VGND sg13g2_decap_8
XFILLER_35_686 VPWR VGND sg13g2_decap_8
XFILLER_34_196 VPWR VGND sg13g2_decap_8
XFILLER_45_406 VPWR VGND sg13g2_decap_8
Xheichips25_template_31 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_26_620 VPWR VGND sg13g2_decap_8
XFILLER_25_130 VPWR VGND sg13g2_decap_8
XFILLER_41_623 VPWR VGND sg13g2_decap_8
XFILLER_13_314 VPWR VGND sg13g2_decap_8
XFILLER_26_697 VPWR VGND sg13g2_decap_8
XFILLER_9_307 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_22_870 VPWR VGND sg13g2_decap_8
XFILLER_5_535 VPWR VGND sg13g2_decap_8
XFILLER_31_63 VPWR VGND sg13g2_decap_8
Xoutput6 net6 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_763 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_49_767 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_36_406 VPWR VGND sg13g2_decap_8
XFILLER_29_480 VPWR VGND sg13g2_decap_8
XFILLER_45_973 VPWR VGND sg13g2_decap_8
XFILLER_44_483 VPWR VGND sg13g2_decap_8
XFILLER_16_174 VPWR VGND sg13g2_decap_8
XFILLER_17_675 VPWR VGND sg13g2_decap_8
XFILLER_32_623 VPWR VGND sg13g2_decap_8
XFILLER_31_133 VPWR VGND sg13g2_decap_8
XFILLER_13_881 VPWR VGND sg13g2_decap_8
XFILLER_12_380 VPWR VGND sg13g2_decap_8
XFILLER_8_373 VPWR VGND sg13g2_decap_8
XFILLER_9_874 VPWR VGND sg13g2_decap_8
XFILLER_28_1005 VPWR VGND sg13g2_decap_8
.ends

