module heichips25_template (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net1;
 wire net2;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;

 sg13g2_inv_1 _31_ (.Y(_08_),
    .A(net44));
 sg13g2_inv_1 _32_ (.Y(_09_),
    .A(net1));
 sg13g2_and3_1 _33_ (.X(_10_),
    .A(net2),
    .B(net34),
    .C(net3));
 sg13g2_and3_1 _34_ (.X(_11_),
    .A(net44),
    .B(net41),
    .C(net5));
 sg13g2_and2_1 _35_ (.A(_10_),
    .B(_11_),
    .X(_12_));
 sg13g2_o21ai_1 _36_ (.B1(net1),
    .Y(_13_),
    .A1(net46),
    .A2(_12_));
 sg13g2_a21oi_1 _37_ (.A1(net46),
    .A2(_12_),
    .Y(_00_),
    .B1(_13_));
 sg13g2_a21oi_1 _38_ (.A1(net8),
    .A2(_12_),
    .Y(_14_),
    .B1(net38));
 sg13g2_and4_1 _39_ (.A(net38),
    .B(net8),
    .C(_10_),
    .D(_11_),
    .X(_15_));
 sg13g2_nor3_1 _40_ (.A(_09_),
    .B(net39),
    .C(_15_),
    .Y(_01_));
 sg13g2_o21ai_1 _41_ (.B1(net1),
    .Y(_16_),
    .A1(net36),
    .A2(_15_));
 sg13g2_a21oi_1 _42_ (.A1(net36),
    .A2(_15_),
    .Y(_02_),
    .B1(_16_));
 sg13g2_o21ai_1 _43_ (.B1(net1),
    .Y(_17_),
    .A1(net2),
    .A2(net47));
 sg13g2_a21oi_1 _44_ (.A1(net2),
    .A2(net47),
    .Y(_03_),
    .B1(_17_));
 sg13g2_a21oi_1 _45_ (.A1(net2),
    .A2(net3),
    .Y(_18_),
    .B1(net34));
 sg13g2_nor3_1 _46_ (.A(_09_),
    .B(_10_),
    .C(net35),
    .Y(_04_));
 sg13g2_o21ai_1 _47_ (.B1(net1),
    .Y(_19_),
    .A1(net48),
    .A2(_10_));
 sg13g2_a21oi_1 _48_ (.A1(net48),
    .A2(_10_),
    .Y(_05_),
    .B1(_19_));
 sg13g2_a21oi_1 _49_ (.A1(net5),
    .A2(_10_),
    .Y(_20_),
    .B1(net41));
 sg13g2_nand3_1 _50_ (.B(net5),
    .C(_10_),
    .A(net41),
    .Y(_21_));
 sg13g2_nand2_1 _51_ (.Y(_22_),
    .A(net1),
    .B(_21_));
 sg13g2_nor2_1 _52_ (.A(net42),
    .B(_22_),
    .Y(_06_));
 sg13g2_a221oi_1 _53_ (.B2(_08_),
    .C1(_09_),
    .B1(_21_),
    .A1(_10_),
    .Y(_07_),
    .A2(_11_));
 sg13g2_dfrbpq_1 _54_ (.RESET_B(net25),
    .D(_00_),
    .Q(net8),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _55_ (.RESET_B(net24),
    .D(net40),
    .Q(net9),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _56_ (.RESET_B(net22),
    .D(net37),
    .Q(net10),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _57_ (.RESET_B(net20),
    .D(_03_),
    .Q(net3),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _58_ (.RESET_B(net),
    .D(_04_),
    .Q(net4),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _59_ (.RESET_B(net23),
    .D(_05_),
    .Q(net5),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _60_ (.RESET_B(net19),
    .D(net43),
    .Q(net6),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _61_ (.RESET_B(net21),
    .D(net45),
    .Q(net7),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_tiehi _60__20 (.L_HI(net19));
 sg13g2_tiehi _57__21 (.L_HI(net20));
 sg13g2_tiehi _61__22 (.L_HI(net21));
 sg13g2_tiehi _56__23 (.L_HI(net22));
 sg13g2_tiehi _59__24 (.L_HI(net23));
 sg13g2_tiehi _55__25 (.L_HI(net24));
 sg13g2_tiehi _54__26 (.L_HI(net25));
 sg13g2_tiehi heichips25_template (.L_HI(net26));
 sg13g2_tiehi heichips25_template_27 (.L_HI(net27));
 sg13g2_tiehi heichips25_template_28 (.L_HI(net28));
 sg13g2_tiehi heichips25_template_29 (.L_HI(net29));
 sg13g2_tiehi heichips25_template_30 (.L_HI(net30));
 sg13g2_tiehi heichips25_template_31 (.L_HI(net31));
 sg13g2_tiehi heichips25_template_32 (.L_HI(net32));
 sg13g2_tiehi heichips25_template_33 (.L_HI(net33));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_1 _78_ (.A(net3),
    .X(net11));
 sg13g2_buf_1 _79_ (.A(net4),
    .X(net12));
 sg13g2_buf_1 _80_ (.A(net5),
    .X(net13));
 sg13g2_buf_1 _81_ (.A(net6),
    .X(net14));
 sg13g2_buf_1 _82_ (.A(net7),
    .X(net15));
 sg13g2_buf_1 _83_ (.A(net8),
    .X(net16));
 sg13g2_buf_1 _84_ (.A(net9),
    .X(net17));
 sg13g2_buf_1 _85_ (.A(net10),
    .X(net18));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_tiehi _58__19 (.L_HI(net));
 sg13g2_buf_16 clkbuf_1_0__f_clk (.X(clknet_1_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_1_1__f_clk (.X(clknet_1_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold34 (.A(net4),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold35 (.A(_18_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold36 (.A(net10),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold37 (.A(_02_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold38 (.A(net9),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold39 (.A(_14_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold40 (.A(_01_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold41 (.A(net6),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold42 (.A(_20_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold43 (.A(_06_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold44 (.A(net7),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold45 (.A(_07_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold46 (.A(net8),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold47 (.A(net3),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold48 (.A(net5),
    .X(net48));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_fill_2 FILLER_2_18 ();
 sg13g2_fill_1 FILLER_2_20 ();
 sg13g2_decap_4 FILLER_2_25 ();
 sg13g2_fill_2 FILLER_2_29 ();
 sg13g2_decap_8 FILLER_2_58 ();
 sg13g2_decap_8 FILLER_2_65 ();
 sg13g2_decap_8 FILLER_2_72 ();
 sg13g2_decap_8 FILLER_2_79 ();
 sg13g2_decap_8 FILLER_2_86 ();
 sg13g2_fill_1 FILLER_2_93 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_4 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_40 ();
 sg13g2_decap_8 FILLER_3_47 ();
 sg13g2_decap_8 FILLER_3_54 ();
 sg13g2_decap_8 FILLER_3_61 ();
 sg13g2_decap_8 FILLER_3_68 ();
 sg13g2_decap_8 FILLER_3_75 ();
 sg13g2_decap_8 FILLER_3_82 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_424 ();
 sg13g2_decap_8 FILLER_3_431 ();
 sg13g2_decap_8 FILLER_3_438 ();
 sg13g2_decap_8 FILLER_3_445 ();
 sg13g2_decap_8 FILLER_3_452 ();
 sg13g2_decap_8 FILLER_3_459 ();
 sg13g2_decap_8 FILLER_3_466 ();
 sg13g2_decap_8 FILLER_3_473 ();
 sg13g2_decap_8 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_decap_8 FILLER_3_494 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_522 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_557 ();
 sg13g2_decap_8 FILLER_3_564 ();
 sg13g2_decap_8 FILLER_3_571 ();
 sg13g2_decap_8 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_585 ();
 sg13g2_decap_8 FILLER_3_592 ();
 sg13g2_decap_8 FILLER_3_599 ();
 sg13g2_decap_8 FILLER_3_606 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_decap_8 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_648 ();
 sg13g2_decap_8 FILLER_3_655 ();
 sg13g2_decap_8 FILLER_3_662 ();
 sg13g2_decap_8 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_676 ();
 sg13g2_decap_8 FILLER_3_683 ();
 sg13g2_decap_8 FILLER_3_690 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_8 FILLER_3_704 ();
 sg13g2_decap_8 FILLER_3_711 ();
 sg13g2_decap_8 FILLER_3_718 ();
 sg13g2_decap_8 FILLER_3_725 ();
 sg13g2_decap_8 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_8 FILLER_3_746 ();
 sg13g2_decap_8 FILLER_3_753 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_decap_8 FILLER_3_767 ();
 sg13g2_decap_8 FILLER_3_774 ();
 sg13g2_decap_8 FILLER_3_781 ();
 sg13g2_decap_8 FILLER_3_788 ();
 sg13g2_decap_8 FILLER_3_795 ();
 sg13g2_decap_8 FILLER_3_802 ();
 sg13g2_decap_8 FILLER_3_809 ();
 sg13g2_decap_8 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_3_823 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_837 ();
 sg13g2_decap_8 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_decap_8 FILLER_3_858 ();
 sg13g2_decap_8 FILLER_3_865 ();
 sg13g2_decap_8 FILLER_3_872 ();
 sg13g2_decap_8 FILLER_3_879 ();
 sg13g2_decap_8 FILLER_3_886 ();
 sg13g2_decap_8 FILLER_3_893 ();
 sg13g2_decap_8 FILLER_3_900 ();
 sg13g2_decap_8 FILLER_3_907 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_8 FILLER_3_921 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_decap_8 FILLER_3_935 ();
 sg13g2_decap_8 FILLER_3_942 ();
 sg13g2_decap_8 FILLER_3_949 ();
 sg13g2_decap_8 FILLER_3_956 ();
 sg13g2_decap_8 FILLER_3_963 ();
 sg13g2_decap_8 FILLER_3_970 ();
 sg13g2_decap_8 FILLER_3_977 ();
 sg13g2_decap_8 FILLER_3_984 ();
 sg13g2_decap_8 FILLER_3_991 ();
 sg13g2_decap_8 FILLER_3_998 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_fill_2 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_fill_2 FILLER_4_18 ();
 sg13g2_fill_1 FILLER_4_20 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_4 FILLER_4_32 ();
 sg13g2_fill_2 FILLER_4_45 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_4 FILLER_4_84 ();
 sg13g2_fill_2 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_fill_2 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_113 ();
 sg13g2_decap_8 FILLER_4_120 ();
 sg13g2_decap_8 FILLER_4_127 ();
 sg13g2_decap_8 FILLER_4_134 ();
 sg13g2_decap_8 FILLER_4_141 ();
 sg13g2_decap_8 FILLER_4_148 ();
 sg13g2_decap_8 FILLER_4_155 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_decap_8 FILLER_4_169 ();
 sg13g2_decap_8 FILLER_4_176 ();
 sg13g2_decap_8 FILLER_4_183 ();
 sg13g2_decap_8 FILLER_4_190 ();
 sg13g2_decap_8 FILLER_4_197 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_decap_8 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_246 ();
 sg13g2_decap_8 FILLER_4_253 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_decap_8 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_4_414 ();
 sg13g2_decap_8 FILLER_4_421 ();
 sg13g2_decap_8 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_4_435 ();
 sg13g2_decap_8 FILLER_4_442 ();
 sg13g2_decap_8 FILLER_4_449 ();
 sg13g2_decap_8 FILLER_4_456 ();
 sg13g2_decap_8 FILLER_4_463 ();
 sg13g2_decap_8 FILLER_4_470 ();
 sg13g2_decap_8 FILLER_4_477 ();
 sg13g2_decap_8 FILLER_4_484 ();
 sg13g2_decap_8 FILLER_4_491 ();
 sg13g2_decap_8 FILLER_4_498 ();
 sg13g2_decap_8 FILLER_4_505 ();
 sg13g2_decap_8 FILLER_4_512 ();
 sg13g2_decap_8 FILLER_4_519 ();
 sg13g2_decap_8 FILLER_4_526 ();
 sg13g2_decap_8 FILLER_4_533 ();
 sg13g2_decap_8 FILLER_4_540 ();
 sg13g2_decap_8 FILLER_4_547 ();
 sg13g2_decap_8 FILLER_4_554 ();
 sg13g2_decap_8 FILLER_4_561 ();
 sg13g2_decap_8 FILLER_4_568 ();
 sg13g2_decap_8 FILLER_4_575 ();
 sg13g2_decap_8 FILLER_4_582 ();
 sg13g2_decap_8 FILLER_4_589 ();
 sg13g2_decap_8 FILLER_4_596 ();
 sg13g2_decap_8 FILLER_4_603 ();
 sg13g2_decap_8 FILLER_4_610 ();
 sg13g2_decap_8 FILLER_4_617 ();
 sg13g2_decap_8 FILLER_4_624 ();
 sg13g2_decap_8 FILLER_4_631 ();
 sg13g2_decap_8 FILLER_4_638 ();
 sg13g2_decap_8 FILLER_4_645 ();
 sg13g2_decap_8 FILLER_4_652 ();
 sg13g2_decap_8 FILLER_4_659 ();
 sg13g2_decap_8 FILLER_4_666 ();
 sg13g2_decap_8 FILLER_4_673 ();
 sg13g2_decap_8 FILLER_4_680 ();
 sg13g2_decap_8 FILLER_4_687 ();
 sg13g2_decap_8 FILLER_4_694 ();
 sg13g2_decap_8 FILLER_4_701 ();
 sg13g2_decap_8 FILLER_4_708 ();
 sg13g2_decap_8 FILLER_4_715 ();
 sg13g2_decap_8 FILLER_4_722 ();
 sg13g2_decap_8 FILLER_4_729 ();
 sg13g2_decap_8 FILLER_4_736 ();
 sg13g2_decap_8 FILLER_4_743 ();
 sg13g2_decap_8 FILLER_4_750 ();
 sg13g2_decap_8 FILLER_4_757 ();
 sg13g2_decap_8 FILLER_4_764 ();
 sg13g2_decap_8 FILLER_4_771 ();
 sg13g2_decap_8 FILLER_4_778 ();
 sg13g2_decap_8 FILLER_4_785 ();
 sg13g2_decap_8 FILLER_4_792 ();
 sg13g2_decap_8 FILLER_4_799 ();
 sg13g2_decap_8 FILLER_4_806 ();
 sg13g2_decap_8 FILLER_4_813 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_decap_8 FILLER_4_827 ();
 sg13g2_decap_8 FILLER_4_834 ();
 sg13g2_decap_8 FILLER_4_841 ();
 sg13g2_decap_8 FILLER_4_848 ();
 sg13g2_decap_8 FILLER_4_855 ();
 sg13g2_decap_8 FILLER_4_862 ();
 sg13g2_decap_8 FILLER_4_869 ();
 sg13g2_decap_8 FILLER_4_876 ();
 sg13g2_decap_8 FILLER_4_883 ();
 sg13g2_decap_8 FILLER_4_890 ();
 sg13g2_decap_8 FILLER_4_897 ();
 sg13g2_decap_8 FILLER_4_904 ();
 sg13g2_decap_8 FILLER_4_911 ();
 sg13g2_decap_8 FILLER_4_918 ();
 sg13g2_decap_8 FILLER_4_925 ();
 sg13g2_decap_8 FILLER_4_932 ();
 sg13g2_decap_8 FILLER_4_939 ();
 sg13g2_decap_8 FILLER_4_946 ();
 sg13g2_decap_8 FILLER_4_953 ();
 sg13g2_decap_8 FILLER_4_960 ();
 sg13g2_decap_8 FILLER_4_967 ();
 sg13g2_decap_8 FILLER_4_974 ();
 sg13g2_decap_8 FILLER_4_981 ();
 sg13g2_decap_8 FILLER_4_988 ();
 sg13g2_decap_8 FILLER_4_995 ();
 sg13g2_decap_8 FILLER_4_1002 ();
 sg13g2_decap_8 FILLER_4_1009 ();
 sg13g2_decap_8 FILLER_4_1016 ();
 sg13g2_decap_4 FILLER_4_1023 ();
 sg13g2_fill_2 FILLER_4_1027 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_fill_2 FILLER_5_18 ();
 sg13g2_fill_1 FILLER_5_20 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_fill_1 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_4 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_94 ();
 sg13g2_decap_8 FILLER_5_101 ();
 sg13g2_decap_8 FILLER_5_108 ();
 sg13g2_decap_8 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_122 ();
 sg13g2_decap_8 FILLER_5_129 ();
 sg13g2_decap_8 FILLER_5_136 ();
 sg13g2_decap_8 FILLER_5_143 ();
 sg13g2_decap_8 FILLER_5_150 ();
 sg13g2_decap_8 FILLER_5_157 ();
 sg13g2_decap_8 FILLER_5_164 ();
 sg13g2_decap_8 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_decap_8 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_206 ();
 sg13g2_decap_8 FILLER_5_213 ();
 sg13g2_decap_8 FILLER_5_220 ();
 sg13g2_decap_8 FILLER_5_227 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_decap_8 FILLER_5_262 ();
 sg13g2_decap_8 FILLER_5_269 ();
 sg13g2_decap_8 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_5_430 ();
 sg13g2_decap_8 FILLER_5_437 ();
 sg13g2_decap_8 FILLER_5_444 ();
 sg13g2_decap_8 FILLER_5_451 ();
 sg13g2_decap_8 FILLER_5_458 ();
 sg13g2_decap_8 FILLER_5_465 ();
 sg13g2_decap_8 FILLER_5_472 ();
 sg13g2_decap_8 FILLER_5_479 ();
 sg13g2_decap_8 FILLER_5_486 ();
 sg13g2_decap_8 FILLER_5_493 ();
 sg13g2_decap_8 FILLER_5_500 ();
 sg13g2_decap_8 FILLER_5_507 ();
 sg13g2_decap_8 FILLER_5_514 ();
 sg13g2_decap_8 FILLER_5_521 ();
 sg13g2_decap_8 FILLER_5_528 ();
 sg13g2_decap_8 FILLER_5_535 ();
 sg13g2_decap_8 FILLER_5_542 ();
 sg13g2_decap_8 FILLER_5_549 ();
 sg13g2_decap_8 FILLER_5_556 ();
 sg13g2_decap_8 FILLER_5_563 ();
 sg13g2_decap_8 FILLER_5_570 ();
 sg13g2_decap_8 FILLER_5_577 ();
 sg13g2_decap_8 FILLER_5_584 ();
 sg13g2_decap_8 FILLER_5_591 ();
 sg13g2_decap_8 FILLER_5_598 ();
 sg13g2_decap_8 FILLER_5_605 ();
 sg13g2_decap_8 FILLER_5_612 ();
 sg13g2_decap_8 FILLER_5_619 ();
 sg13g2_decap_8 FILLER_5_626 ();
 sg13g2_decap_8 FILLER_5_633 ();
 sg13g2_decap_8 FILLER_5_640 ();
 sg13g2_decap_8 FILLER_5_647 ();
 sg13g2_decap_8 FILLER_5_654 ();
 sg13g2_decap_8 FILLER_5_661 ();
 sg13g2_decap_8 FILLER_5_668 ();
 sg13g2_decap_8 FILLER_5_675 ();
 sg13g2_decap_8 FILLER_5_682 ();
 sg13g2_decap_8 FILLER_5_689 ();
 sg13g2_decap_8 FILLER_5_696 ();
 sg13g2_decap_8 FILLER_5_703 ();
 sg13g2_decap_8 FILLER_5_710 ();
 sg13g2_decap_8 FILLER_5_717 ();
 sg13g2_decap_8 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_731 ();
 sg13g2_decap_8 FILLER_5_738 ();
 sg13g2_decap_8 FILLER_5_745 ();
 sg13g2_decap_8 FILLER_5_752 ();
 sg13g2_decap_8 FILLER_5_759 ();
 sg13g2_decap_8 FILLER_5_766 ();
 sg13g2_decap_8 FILLER_5_773 ();
 sg13g2_decap_8 FILLER_5_780 ();
 sg13g2_decap_8 FILLER_5_787 ();
 sg13g2_decap_8 FILLER_5_794 ();
 sg13g2_decap_8 FILLER_5_801 ();
 sg13g2_decap_8 FILLER_5_808 ();
 sg13g2_decap_8 FILLER_5_815 ();
 sg13g2_decap_8 FILLER_5_822 ();
 sg13g2_decap_8 FILLER_5_829 ();
 sg13g2_decap_8 FILLER_5_836 ();
 sg13g2_decap_8 FILLER_5_843 ();
 sg13g2_decap_8 FILLER_5_850 ();
 sg13g2_decap_8 FILLER_5_857 ();
 sg13g2_decap_8 FILLER_5_864 ();
 sg13g2_decap_8 FILLER_5_871 ();
 sg13g2_decap_8 FILLER_5_878 ();
 sg13g2_decap_8 FILLER_5_885 ();
 sg13g2_decap_8 FILLER_5_892 ();
 sg13g2_decap_8 FILLER_5_899 ();
 sg13g2_decap_8 FILLER_5_906 ();
 sg13g2_decap_8 FILLER_5_913 ();
 sg13g2_decap_8 FILLER_5_920 ();
 sg13g2_decap_8 FILLER_5_927 ();
 sg13g2_decap_8 FILLER_5_934 ();
 sg13g2_decap_8 FILLER_5_941 ();
 sg13g2_decap_8 FILLER_5_948 ();
 sg13g2_decap_8 FILLER_5_955 ();
 sg13g2_decap_8 FILLER_5_962 ();
 sg13g2_decap_8 FILLER_5_969 ();
 sg13g2_decap_8 FILLER_5_976 ();
 sg13g2_decap_8 FILLER_5_983 ();
 sg13g2_decap_8 FILLER_5_990 ();
 sg13g2_decap_8 FILLER_5_997 ();
 sg13g2_decap_8 FILLER_5_1004 ();
 sg13g2_decap_8 FILLER_5_1011 ();
 sg13g2_decap_8 FILLER_5_1018 ();
 sg13g2_decap_4 FILLER_5_1025 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_4 FILLER_6_32 ();
 sg13g2_fill_2 FILLER_6_36 ();
 sg13g2_decap_8 FILLER_6_47 ();
 sg13g2_decap_8 FILLER_6_54 ();
 sg13g2_decap_8 FILLER_6_61 ();
 sg13g2_decap_8 FILLER_6_68 ();
 sg13g2_decap_8 FILLER_6_75 ();
 sg13g2_decap_8 FILLER_6_82 ();
 sg13g2_decap_8 FILLER_6_89 ();
 sg13g2_decap_8 FILLER_6_96 ();
 sg13g2_decap_8 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_124 ();
 sg13g2_decap_8 FILLER_6_131 ();
 sg13g2_decap_8 FILLER_6_138 ();
 sg13g2_decap_8 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_152 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_166 ();
 sg13g2_decap_8 FILLER_6_173 ();
 sg13g2_decap_8 FILLER_6_180 ();
 sg13g2_decap_8 FILLER_6_187 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_decap_8 FILLER_6_201 ();
 sg13g2_decap_8 FILLER_6_208 ();
 sg13g2_decap_8 FILLER_6_215 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_236 ();
 sg13g2_decap_8 FILLER_6_243 ();
 sg13g2_decap_8 FILLER_6_250 ();
 sg13g2_decap_8 FILLER_6_257 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_8 FILLER_6_425 ();
 sg13g2_decap_8 FILLER_6_432 ();
 sg13g2_decap_8 FILLER_6_439 ();
 sg13g2_decap_8 FILLER_6_446 ();
 sg13g2_decap_8 FILLER_6_453 ();
 sg13g2_decap_8 FILLER_6_460 ();
 sg13g2_decap_8 FILLER_6_467 ();
 sg13g2_decap_8 FILLER_6_474 ();
 sg13g2_decap_8 FILLER_6_481 ();
 sg13g2_decap_8 FILLER_6_488 ();
 sg13g2_decap_8 FILLER_6_495 ();
 sg13g2_decap_8 FILLER_6_502 ();
 sg13g2_decap_8 FILLER_6_509 ();
 sg13g2_decap_8 FILLER_6_516 ();
 sg13g2_decap_8 FILLER_6_523 ();
 sg13g2_decap_8 FILLER_6_530 ();
 sg13g2_decap_8 FILLER_6_537 ();
 sg13g2_decap_8 FILLER_6_544 ();
 sg13g2_decap_8 FILLER_6_551 ();
 sg13g2_decap_8 FILLER_6_558 ();
 sg13g2_decap_8 FILLER_6_565 ();
 sg13g2_decap_8 FILLER_6_572 ();
 sg13g2_decap_8 FILLER_6_579 ();
 sg13g2_decap_8 FILLER_6_586 ();
 sg13g2_decap_8 FILLER_6_593 ();
 sg13g2_decap_8 FILLER_6_600 ();
 sg13g2_decap_8 FILLER_6_607 ();
 sg13g2_decap_8 FILLER_6_614 ();
 sg13g2_decap_8 FILLER_6_621 ();
 sg13g2_decap_8 FILLER_6_628 ();
 sg13g2_decap_8 FILLER_6_635 ();
 sg13g2_decap_8 FILLER_6_642 ();
 sg13g2_decap_8 FILLER_6_649 ();
 sg13g2_decap_8 FILLER_6_656 ();
 sg13g2_decap_8 FILLER_6_663 ();
 sg13g2_decap_8 FILLER_6_670 ();
 sg13g2_decap_8 FILLER_6_677 ();
 sg13g2_decap_8 FILLER_6_684 ();
 sg13g2_decap_8 FILLER_6_691 ();
 sg13g2_decap_8 FILLER_6_698 ();
 sg13g2_decap_8 FILLER_6_705 ();
 sg13g2_decap_8 FILLER_6_712 ();
 sg13g2_decap_8 FILLER_6_719 ();
 sg13g2_decap_8 FILLER_6_726 ();
 sg13g2_decap_8 FILLER_6_733 ();
 sg13g2_decap_8 FILLER_6_740 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_8 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_768 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_8 FILLER_6_789 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_decap_8 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_831 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_decap_8 FILLER_6_859 ();
 sg13g2_decap_8 FILLER_6_866 ();
 sg13g2_decap_8 FILLER_6_873 ();
 sg13g2_decap_8 FILLER_6_880 ();
 sg13g2_decap_8 FILLER_6_887 ();
 sg13g2_decap_8 FILLER_6_894 ();
 sg13g2_decap_8 FILLER_6_901 ();
 sg13g2_decap_8 FILLER_6_908 ();
 sg13g2_decap_8 FILLER_6_915 ();
 sg13g2_decap_8 FILLER_6_922 ();
 sg13g2_decap_8 FILLER_6_929 ();
 sg13g2_decap_8 FILLER_6_936 ();
 sg13g2_decap_8 FILLER_6_943 ();
 sg13g2_decap_8 FILLER_6_950 ();
 sg13g2_decap_8 FILLER_6_957 ();
 sg13g2_decap_8 FILLER_6_964 ();
 sg13g2_decap_8 FILLER_6_971 ();
 sg13g2_decap_8 FILLER_6_978 ();
 sg13g2_decap_8 FILLER_6_985 ();
 sg13g2_decap_8 FILLER_6_992 ();
 sg13g2_decap_8 FILLER_6_999 ();
 sg13g2_decap_8 FILLER_6_1006 ();
 sg13g2_decap_8 FILLER_6_1013 ();
 sg13g2_decap_8 FILLER_6_1020 ();
 sg13g2_fill_2 FILLER_6_1027 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_25 ();
 sg13g2_decap_8 FILLER_7_32 ();
 sg13g2_decap_4 FILLER_7_39 ();
 sg13g2_decap_8 FILLER_7_47 ();
 sg13g2_decap_8 FILLER_7_54 ();
 sg13g2_decap_8 FILLER_7_61 ();
 sg13g2_decap_8 FILLER_7_68 ();
 sg13g2_decap_8 FILLER_7_75 ();
 sg13g2_decap_8 FILLER_7_82 ();
 sg13g2_decap_8 FILLER_7_89 ();
 sg13g2_decap_8 FILLER_7_96 ();
 sg13g2_decap_8 FILLER_7_103 ();
 sg13g2_decap_8 FILLER_7_110 ();
 sg13g2_decap_8 FILLER_7_117 ();
 sg13g2_decap_8 FILLER_7_124 ();
 sg13g2_decap_8 FILLER_7_131 ();
 sg13g2_decap_8 FILLER_7_138 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_152 ();
 sg13g2_decap_8 FILLER_7_159 ();
 sg13g2_decap_8 FILLER_7_166 ();
 sg13g2_decap_8 FILLER_7_173 ();
 sg13g2_decap_8 FILLER_7_180 ();
 sg13g2_decap_8 FILLER_7_187 ();
 sg13g2_decap_8 FILLER_7_194 ();
 sg13g2_decap_8 FILLER_7_201 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_decap_8 FILLER_7_215 ();
 sg13g2_decap_8 FILLER_7_222 ();
 sg13g2_decap_8 FILLER_7_229 ();
 sg13g2_decap_8 FILLER_7_236 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_8 FILLER_7_250 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_decap_8 FILLER_7_264 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_8 FILLER_7_404 ();
 sg13g2_decap_8 FILLER_7_411 ();
 sg13g2_decap_8 FILLER_7_418 ();
 sg13g2_decap_8 FILLER_7_425 ();
 sg13g2_decap_8 FILLER_7_432 ();
 sg13g2_decap_8 FILLER_7_439 ();
 sg13g2_decap_8 FILLER_7_446 ();
 sg13g2_decap_8 FILLER_7_453 ();
 sg13g2_decap_8 FILLER_7_460 ();
 sg13g2_decap_8 FILLER_7_467 ();
 sg13g2_decap_8 FILLER_7_474 ();
 sg13g2_decap_8 FILLER_7_481 ();
 sg13g2_decap_8 FILLER_7_488 ();
 sg13g2_decap_8 FILLER_7_495 ();
 sg13g2_decap_8 FILLER_7_502 ();
 sg13g2_decap_8 FILLER_7_509 ();
 sg13g2_decap_8 FILLER_7_516 ();
 sg13g2_decap_8 FILLER_7_523 ();
 sg13g2_decap_8 FILLER_7_530 ();
 sg13g2_decap_8 FILLER_7_537 ();
 sg13g2_decap_8 FILLER_7_544 ();
 sg13g2_decap_8 FILLER_7_551 ();
 sg13g2_decap_8 FILLER_7_558 ();
 sg13g2_decap_8 FILLER_7_565 ();
 sg13g2_decap_8 FILLER_7_572 ();
 sg13g2_decap_8 FILLER_7_579 ();
 sg13g2_decap_8 FILLER_7_586 ();
 sg13g2_decap_8 FILLER_7_593 ();
 sg13g2_decap_8 FILLER_7_600 ();
 sg13g2_decap_8 FILLER_7_607 ();
 sg13g2_decap_8 FILLER_7_614 ();
 sg13g2_decap_8 FILLER_7_621 ();
 sg13g2_decap_8 FILLER_7_628 ();
 sg13g2_decap_8 FILLER_7_635 ();
 sg13g2_decap_8 FILLER_7_642 ();
 sg13g2_decap_8 FILLER_7_649 ();
 sg13g2_decap_8 FILLER_7_656 ();
 sg13g2_decap_8 FILLER_7_663 ();
 sg13g2_decap_8 FILLER_7_670 ();
 sg13g2_decap_8 FILLER_7_677 ();
 sg13g2_decap_8 FILLER_7_684 ();
 sg13g2_decap_8 FILLER_7_691 ();
 sg13g2_decap_8 FILLER_7_698 ();
 sg13g2_decap_8 FILLER_7_705 ();
 sg13g2_decap_8 FILLER_7_712 ();
 sg13g2_decap_8 FILLER_7_719 ();
 sg13g2_decap_8 FILLER_7_726 ();
 sg13g2_decap_8 FILLER_7_733 ();
 sg13g2_decap_8 FILLER_7_740 ();
 sg13g2_decap_8 FILLER_7_747 ();
 sg13g2_decap_8 FILLER_7_754 ();
 sg13g2_decap_8 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_768 ();
 sg13g2_decap_8 FILLER_7_775 ();
 sg13g2_decap_8 FILLER_7_782 ();
 sg13g2_decap_8 FILLER_7_789 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_decap_8 FILLER_7_803 ();
 sg13g2_decap_8 FILLER_7_810 ();
 sg13g2_decap_8 FILLER_7_817 ();
 sg13g2_decap_8 FILLER_7_824 ();
 sg13g2_decap_8 FILLER_7_831 ();
 sg13g2_decap_8 FILLER_7_838 ();
 sg13g2_decap_8 FILLER_7_845 ();
 sg13g2_decap_8 FILLER_7_852 ();
 sg13g2_decap_8 FILLER_7_859 ();
 sg13g2_decap_8 FILLER_7_866 ();
 sg13g2_decap_8 FILLER_7_873 ();
 sg13g2_decap_8 FILLER_7_880 ();
 sg13g2_decap_8 FILLER_7_887 ();
 sg13g2_decap_8 FILLER_7_894 ();
 sg13g2_decap_8 FILLER_7_901 ();
 sg13g2_decap_8 FILLER_7_908 ();
 sg13g2_decap_8 FILLER_7_915 ();
 sg13g2_decap_8 FILLER_7_922 ();
 sg13g2_decap_8 FILLER_7_929 ();
 sg13g2_decap_8 FILLER_7_936 ();
 sg13g2_decap_8 FILLER_7_943 ();
 sg13g2_decap_8 FILLER_7_950 ();
 sg13g2_decap_8 FILLER_7_957 ();
 sg13g2_decap_8 FILLER_7_964 ();
 sg13g2_decap_8 FILLER_7_971 ();
 sg13g2_decap_8 FILLER_7_978 ();
 sg13g2_decap_8 FILLER_7_985 ();
 sg13g2_decap_8 FILLER_7_992 ();
 sg13g2_decap_8 FILLER_7_999 ();
 sg13g2_decap_8 FILLER_7_1006 ();
 sg13g2_decap_8 FILLER_7_1013 ();
 sg13g2_decap_8 FILLER_7_1020 ();
 sg13g2_fill_2 FILLER_7_1027 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_fill_2 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_4 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_113 ();
 sg13g2_decap_8 FILLER_8_142 ();
 sg13g2_decap_8 FILLER_8_149 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_decap_8 FILLER_8_163 ();
 sg13g2_decap_8 FILLER_8_170 ();
 sg13g2_decap_8 FILLER_8_177 ();
 sg13g2_decap_8 FILLER_8_184 ();
 sg13g2_decap_8 FILLER_8_191 ();
 sg13g2_decap_8 FILLER_8_198 ();
 sg13g2_decap_8 FILLER_8_205 ();
 sg13g2_decap_8 FILLER_8_212 ();
 sg13g2_decap_8 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_decap_8 FILLER_8_240 ();
 sg13g2_decap_8 FILLER_8_247 ();
 sg13g2_decap_8 FILLER_8_254 ();
 sg13g2_decap_8 FILLER_8_261 ();
 sg13g2_decap_8 FILLER_8_268 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_decap_8 FILLER_8_289 ();
 sg13g2_decap_8 FILLER_8_296 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_310 ();
 sg13g2_decap_8 FILLER_8_317 ();
 sg13g2_decap_8 FILLER_8_324 ();
 sg13g2_decap_8 FILLER_8_331 ();
 sg13g2_decap_8 FILLER_8_338 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_8 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_415 ();
 sg13g2_decap_8 FILLER_8_422 ();
 sg13g2_decap_8 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_8_436 ();
 sg13g2_decap_8 FILLER_8_443 ();
 sg13g2_decap_8 FILLER_8_450 ();
 sg13g2_decap_8 FILLER_8_457 ();
 sg13g2_decap_8 FILLER_8_464 ();
 sg13g2_decap_8 FILLER_8_471 ();
 sg13g2_decap_8 FILLER_8_478 ();
 sg13g2_decap_8 FILLER_8_485 ();
 sg13g2_decap_8 FILLER_8_492 ();
 sg13g2_decap_8 FILLER_8_499 ();
 sg13g2_decap_8 FILLER_8_506 ();
 sg13g2_decap_8 FILLER_8_513 ();
 sg13g2_decap_8 FILLER_8_520 ();
 sg13g2_decap_8 FILLER_8_527 ();
 sg13g2_decap_8 FILLER_8_534 ();
 sg13g2_decap_8 FILLER_8_541 ();
 sg13g2_decap_8 FILLER_8_548 ();
 sg13g2_decap_8 FILLER_8_555 ();
 sg13g2_decap_8 FILLER_8_562 ();
 sg13g2_decap_8 FILLER_8_569 ();
 sg13g2_decap_8 FILLER_8_576 ();
 sg13g2_decap_8 FILLER_8_583 ();
 sg13g2_decap_8 FILLER_8_590 ();
 sg13g2_decap_8 FILLER_8_597 ();
 sg13g2_decap_8 FILLER_8_604 ();
 sg13g2_decap_8 FILLER_8_611 ();
 sg13g2_decap_8 FILLER_8_618 ();
 sg13g2_decap_8 FILLER_8_625 ();
 sg13g2_decap_8 FILLER_8_632 ();
 sg13g2_decap_8 FILLER_8_639 ();
 sg13g2_decap_8 FILLER_8_646 ();
 sg13g2_decap_8 FILLER_8_653 ();
 sg13g2_decap_8 FILLER_8_660 ();
 sg13g2_decap_8 FILLER_8_667 ();
 sg13g2_decap_8 FILLER_8_674 ();
 sg13g2_decap_8 FILLER_8_681 ();
 sg13g2_decap_8 FILLER_8_688 ();
 sg13g2_decap_8 FILLER_8_695 ();
 sg13g2_decap_8 FILLER_8_702 ();
 sg13g2_decap_8 FILLER_8_709 ();
 sg13g2_decap_8 FILLER_8_716 ();
 sg13g2_decap_8 FILLER_8_723 ();
 sg13g2_decap_8 FILLER_8_730 ();
 sg13g2_decap_8 FILLER_8_737 ();
 sg13g2_decap_8 FILLER_8_744 ();
 sg13g2_decap_8 FILLER_8_751 ();
 sg13g2_decap_8 FILLER_8_758 ();
 sg13g2_decap_8 FILLER_8_765 ();
 sg13g2_decap_8 FILLER_8_772 ();
 sg13g2_decap_8 FILLER_8_779 ();
 sg13g2_decap_8 FILLER_8_786 ();
 sg13g2_decap_8 FILLER_8_793 ();
 sg13g2_decap_8 FILLER_8_800 ();
 sg13g2_decap_8 FILLER_8_807 ();
 sg13g2_decap_8 FILLER_8_814 ();
 sg13g2_decap_8 FILLER_8_821 ();
 sg13g2_decap_8 FILLER_8_828 ();
 sg13g2_decap_8 FILLER_8_835 ();
 sg13g2_decap_8 FILLER_8_842 ();
 sg13g2_decap_8 FILLER_8_849 ();
 sg13g2_decap_8 FILLER_8_856 ();
 sg13g2_decap_8 FILLER_8_863 ();
 sg13g2_decap_8 FILLER_8_870 ();
 sg13g2_decap_8 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_8_884 ();
 sg13g2_decap_8 FILLER_8_891 ();
 sg13g2_decap_8 FILLER_8_898 ();
 sg13g2_decap_8 FILLER_8_905 ();
 sg13g2_decap_8 FILLER_8_912 ();
 sg13g2_decap_8 FILLER_8_919 ();
 sg13g2_decap_8 FILLER_8_926 ();
 sg13g2_decap_8 FILLER_8_933 ();
 sg13g2_decap_8 FILLER_8_940 ();
 sg13g2_decap_8 FILLER_8_947 ();
 sg13g2_decap_8 FILLER_8_954 ();
 sg13g2_decap_8 FILLER_8_961 ();
 sg13g2_decap_8 FILLER_8_968 ();
 sg13g2_decap_8 FILLER_8_975 ();
 sg13g2_decap_8 FILLER_8_982 ();
 sg13g2_decap_8 FILLER_8_989 ();
 sg13g2_decap_8 FILLER_8_996 ();
 sg13g2_decap_8 FILLER_8_1003 ();
 sg13g2_decap_8 FILLER_8_1010 ();
 sg13g2_decap_8 FILLER_8_1017 ();
 sg13g2_decap_4 FILLER_8_1024 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_fill_2 FILLER_9_18 ();
 sg13g2_fill_1 FILLER_9_20 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_101 ();
 sg13g2_fill_1 FILLER_9_111 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_132 ();
 sg13g2_decap_8 FILLER_9_139 ();
 sg13g2_decap_8 FILLER_9_146 ();
 sg13g2_decap_8 FILLER_9_153 ();
 sg13g2_decap_8 FILLER_9_160 ();
 sg13g2_decap_8 FILLER_9_167 ();
 sg13g2_decap_8 FILLER_9_174 ();
 sg13g2_decap_8 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_188 ();
 sg13g2_decap_8 FILLER_9_195 ();
 sg13g2_decap_8 FILLER_9_202 ();
 sg13g2_decap_8 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_230 ();
 sg13g2_decap_8 FILLER_9_237 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_265 ();
 sg13g2_decap_8 FILLER_9_272 ();
 sg13g2_decap_8 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_8 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_8 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_9_433 ();
 sg13g2_decap_8 FILLER_9_440 ();
 sg13g2_decap_8 FILLER_9_447 ();
 sg13g2_decap_8 FILLER_9_454 ();
 sg13g2_decap_8 FILLER_9_461 ();
 sg13g2_decap_8 FILLER_9_468 ();
 sg13g2_decap_8 FILLER_9_475 ();
 sg13g2_decap_8 FILLER_9_482 ();
 sg13g2_decap_8 FILLER_9_489 ();
 sg13g2_decap_8 FILLER_9_496 ();
 sg13g2_decap_8 FILLER_9_503 ();
 sg13g2_decap_8 FILLER_9_510 ();
 sg13g2_decap_8 FILLER_9_517 ();
 sg13g2_decap_8 FILLER_9_524 ();
 sg13g2_decap_8 FILLER_9_531 ();
 sg13g2_decap_8 FILLER_9_538 ();
 sg13g2_decap_8 FILLER_9_545 ();
 sg13g2_decap_8 FILLER_9_552 ();
 sg13g2_decap_8 FILLER_9_559 ();
 sg13g2_decap_8 FILLER_9_566 ();
 sg13g2_decap_8 FILLER_9_573 ();
 sg13g2_decap_8 FILLER_9_580 ();
 sg13g2_decap_8 FILLER_9_587 ();
 sg13g2_decap_8 FILLER_9_594 ();
 sg13g2_decap_8 FILLER_9_601 ();
 sg13g2_decap_8 FILLER_9_608 ();
 sg13g2_decap_8 FILLER_9_615 ();
 sg13g2_decap_8 FILLER_9_622 ();
 sg13g2_decap_8 FILLER_9_629 ();
 sg13g2_decap_8 FILLER_9_636 ();
 sg13g2_decap_8 FILLER_9_643 ();
 sg13g2_decap_8 FILLER_9_650 ();
 sg13g2_decap_8 FILLER_9_657 ();
 sg13g2_decap_8 FILLER_9_664 ();
 sg13g2_decap_8 FILLER_9_671 ();
 sg13g2_decap_8 FILLER_9_678 ();
 sg13g2_decap_8 FILLER_9_685 ();
 sg13g2_decap_8 FILLER_9_692 ();
 sg13g2_decap_8 FILLER_9_699 ();
 sg13g2_decap_8 FILLER_9_706 ();
 sg13g2_decap_8 FILLER_9_713 ();
 sg13g2_decap_8 FILLER_9_720 ();
 sg13g2_decap_8 FILLER_9_727 ();
 sg13g2_decap_8 FILLER_9_734 ();
 sg13g2_decap_8 FILLER_9_741 ();
 sg13g2_decap_8 FILLER_9_748 ();
 sg13g2_decap_8 FILLER_9_755 ();
 sg13g2_decap_8 FILLER_9_762 ();
 sg13g2_decap_8 FILLER_9_769 ();
 sg13g2_decap_8 FILLER_9_776 ();
 sg13g2_decap_8 FILLER_9_783 ();
 sg13g2_decap_8 FILLER_9_790 ();
 sg13g2_decap_8 FILLER_9_797 ();
 sg13g2_decap_8 FILLER_9_804 ();
 sg13g2_decap_8 FILLER_9_811 ();
 sg13g2_decap_8 FILLER_9_818 ();
 sg13g2_decap_8 FILLER_9_825 ();
 sg13g2_decap_8 FILLER_9_832 ();
 sg13g2_decap_8 FILLER_9_839 ();
 sg13g2_decap_8 FILLER_9_846 ();
 sg13g2_decap_8 FILLER_9_853 ();
 sg13g2_decap_8 FILLER_9_860 ();
 sg13g2_decap_8 FILLER_9_867 ();
 sg13g2_decap_8 FILLER_9_874 ();
 sg13g2_decap_8 FILLER_9_881 ();
 sg13g2_decap_8 FILLER_9_888 ();
 sg13g2_decap_8 FILLER_9_895 ();
 sg13g2_decap_8 FILLER_9_902 ();
 sg13g2_decap_8 FILLER_9_909 ();
 sg13g2_decap_8 FILLER_9_916 ();
 sg13g2_decap_8 FILLER_9_923 ();
 sg13g2_decap_8 FILLER_9_930 ();
 sg13g2_decap_8 FILLER_9_937 ();
 sg13g2_decap_8 FILLER_9_944 ();
 sg13g2_decap_8 FILLER_9_951 ();
 sg13g2_decap_8 FILLER_9_958 ();
 sg13g2_decap_8 FILLER_9_965 ();
 sg13g2_decap_8 FILLER_9_972 ();
 sg13g2_decap_8 FILLER_9_979 ();
 sg13g2_decap_8 FILLER_9_986 ();
 sg13g2_decap_8 FILLER_9_993 ();
 sg13g2_decap_8 FILLER_9_1000 ();
 sg13g2_decap_8 FILLER_9_1007 ();
 sg13g2_decap_8 FILLER_9_1014 ();
 sg13g2_decap_8 FILLER_9_1021 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_4 FILLER_10_11 ();
 sg13g2_fill_2 FILLER_10_15 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_4 FILLER_10_60 ();
 sg13g2_fill_1 FILLER_10_64 ();
 sg13g2_decap_8 FILLER_10_72 ();
 sg13g2_decap_8 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_86 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_8 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_135 ();
 sg13g2_decap_8 FILLER_10_142 ();
 sg13g2_decap_8 FILLER_10_149 ();
 sg13g2_decap_8 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_decap_8 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_254 ();
 sg13g2_decap_8 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_268 ();
 sg13g2_decap_8 FILLER_10_275 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_decap_8 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_decap_8 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_10_436 ();
 sg13g2_decap_8 FILLER_10_443 ();
 sg13g2_decap_8 FILLER_10_450 ();
 sg13g2_decap_8 FILLER_10_457 ();
 sg13g2_decap_8 FILLER_10_464 ();
 sg13g2_decap_8 FILLER_10_471 ();
 sg13g2_decap_8 FILLER_10_478 ();
 sg13g2_decap_8 FILLER_10_485 ();
 sg13g2_decap_8 FILLER_10_492 ();
 sg13g2_decap_8 FILLER_10_499 ();
 sg13g2_decap_8 FILLER_10_506 ();
 sg13g2_decap_8 FILLER_10_513 ();
 sg13g2_decap_8 FILLER_10_520 ();
 sg13g2_decap_8 FILLER_10_527 ();
 sg13g2_decap_8 FILLER_10_534 ();
 sg13g2_decap_8 FILLER_10_541 ();
 sg13g2_decap_8 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_562 ();
 sg13g2_decap_8 FILLER_10_569 ();
 sg13g2_decap_8 FILLER_10_576 ();
 sg13g2_decap_8 FILLER_10_583 ();
 sg13g2_decap_8 FILLER_10_590 ();
 sg13g2_decap_8 FILLER_10_597 ();
 sg13g2_decap_8 FILLER_10_604 ();
 sg13g2_decap_8 FILLER_10_611 ();
 sg13g2_decap_8 FILLER_10_618 ();
 sg13g2_decap_8 FILLER_10_625 ();
 sg13g2_decap_8 FILLER_10_632 ();
 sg13g2_decap_8 FILLER_10_639 ();
 sg13g2_decap_8 FILLER_10_646 ();
 sg13g2_decap_8 FILLER_10_653 ();
 sg13g2_decap_8 FILLER_10_660 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_decap_8 FILLER_10_674 ();
 sg13g2_decap_8 FILLER_10_681 ();
 sg13g2_decap_8 FILLER_10_688 ();
 sg13g2_decap_8 FILLER_10_695 ();
 sg13g2_decap_8 FILLER_10_702 ();
 sg13g2_decap_8 FILLER_10_709 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_decap_8 FILLER_10_723 ();
 sg13g2_decap_8 FILLER_10_730 ();
 sg13g2_decap_8 FILLER_10_737 ();
 sg13g2_decap_8 FILLER_10_744 ();
 sg13g2_decap_8 FILLER_10_751 ();
 sg13g2_decap_8 FILLER_10_758 ();
 sg13g2_decap_8 FILLER_10_765 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_8 FILLER_10_842 ();
 sg13g2_decap_8 FILLER_10_849 ();
 sg13g2_decap_8 FILLER_10_856 ();
 sg13g2_decap_8 FILLER_10_863 ();
 sg13g2_decap_8 FILLER_10_870 ();
 sg13g2_decap_8 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_10_884 ();
 sg13g2_decap_8 FILLER_10_891 ();
 sg13g2_decap_8 FILLER_10_898 ();
 sg13g2_decap_8 FILLER_10_905 ();
 sg13g2_decap_8 FILLER_10_912 ();
 sg13g2_decap_8 FILLER_10_919 ();
 sg13g2_decap_8 FILLER_10_926 ();
 sg13g2_decap_8 FILLER_10_933 ();
 sg13g2_decap_8 FILLER_10_940 ();
 sg13g2_decap_8 FILLER_10_947 ();
 sg13g2_decap_8 FILLER_10_954 ();
 sg13g2_decap_8 FILLER_10_961 ();
 sg13g2_decap_8 FILLER_10_968 ();
 sg13g2_decap_8 FILLER_10_975 ();
 sg13g2_decap_8 FILLER_10_982 ();
 sg13g2_decap_8 FILLER_10_989 ();
 sg13g2_decap_8 FILLER_10_996 ();
 sg13g2_decap_8 FILLER_10_1003 ();
 sg13g2_decap_8 FILLER_10_1010 ();
 sg13g2_decap_8 FILLER_10_1017 ();
 sg13g2_decap_4 FILLER_10_1024 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_fill_2 FILLER_11_18 ();
 sg13g2_fill_1 FILLER_11_20 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_decap_4 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_decap_8 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_4 FILLER_11_95 ();
 sg13g2_fill_2 FILLER_11_99 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_8 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_decap_8 FILLER_11_875 ();
 sg13g2_decap_8 FILLER_11_882 ();
 sg13g2_decap_8 FILLER_11_889 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_decap_8 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_910 ();
 sg13g2_decap_8 FILLER_11_917 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_decap_8 FILLER_11_945 ();
 sg13g2_decap_8 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_8 FILLER_11_1001 ();
 sg13g2_decap_8 FILLER_11_1008 ();
 sg13g2_decap_8 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1022 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_149 ();
 sg13g2_decap_8 FILLER_12_156 ();
 sg13g2_decap_8 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_170 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_decap_8 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_decap_8 FILLER_12_205 ();
 sg13g2_decap_8 FILLER_12_212 ();
 sg13g2_decap_8 FILLER_12_219 ();
 sg13g2_decap_8 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_8 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_decap_8 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_12_436 ();
 sg13g2_decap_8 FILLER_12_443 ();
 sg13g2_decap_8 FILLER_12_450 ();
 sg13g2_decap_8 FILLER_12_457 ();
 sg13g2_decap_8 FILLER_12_464 ();
 sg13g2_decap_8 FILLER_12_471 ();
 sg13g2_decap_8 FILLER_12_478 ();
 sg13g2_decap_8 FILLER_12_485 ();
 sg13g2_decap_8 FILLER_12_492 ();
 sg13g2_decap_8 FILLER_12_499 ();
 sg13g2_decap_8 FILLER_12_506 ();
 sg13g2_decap_8 FILLER_12_513 ();
 sg13g2_decap_8 FILLER_12_520 ();
 sg13g2_decap_8 FILLER_12_527 ();
 sg13g2_decap_8 FILLER_12_534 ();
 sg13g2_decap_8 FILLER_12_541 ();
 sg13g2_decap_8 FILLER_12_548 ();
 sg13g2_decap_8 FILLER_12_555 ();
 sg13g2_decap_8 FILLER_12_562 ();
 sg13g2_decap_8 FILLER_12_569 ();
 sg13g2_decap_8 FILLER_12_576 ();
 sg13g2_decap_8 FILLER_12_583 ();
 sg13g2_decap_8 FILLER_12_590 ();
 sg13g2_decap_8 FILLER_12_597 ();
 sg13g2_decap_8 FILLER_12_604 ();
 sg13g2_decap_8 FILLER_12_611 ();
 sg13g2_decap_8 FILLER_12_618 ();
 sg13g2_decap_8 FILLER_12_625 ();
 sg13g2_decap_8 FILLER_12_632 ();
 sg13g2_decap_8 FILLER_12_639 ();
 sg13g2_decap_8 FILLER_12_646 ();
 sg13g2_decap_8 FILLER_12_653 ();
 sg13g2_decap_8 FILLER_12_660 ();
 sg13g2_decap_8 FILLER_12_667 ();
 sg13g2_decap_8 FILLER_12_674 ();
 sg13g2_decap_8 FILLER_12_681 ();
 sg13g2_decap_8 FILLER_12_688 ();
 sg13g2_decap_8 FILLER_12_695 ();
 sg13g2_decap_8 FILLER_12_702 ();
 sg13g2_decap_8 FILLER_12_709 ();
 sg13g2_decap_8 FILLER_12_716 ();
 sg13g2_decap_8 FILLER_12_723 ();
 sg13g2_decap_8 FILLER_12_730 ();
 sg13g2_decap_8 FILLER_12_737 ();
 sg13g2_decap_8 FILLER_12_744 ();
 sg13g2_decap_8 FILLER_12_751 ();
 sg13g2_decap_8 FILLER_12_758 ();
 sg13g2_decap_8 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_772 ();
 sg13g2_decap_8 FILLER_12_779 ();
 sg13g2_decap_8 FILLER_12_786 ();
 sg13g2_decap_8 FILLER_12_793 ();
 sg13g2_decap_8 FILLER_12_800 ();
 sg13g2_decap_8 FILLER_12_807 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_8 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_828 ();
 sg13g2_decap_8 FILLER_12_835 ();
 sg13g2_decap_8 FILLER_12_842 ();
 sg13g2_decap_8 FILLER_12_849 ();
 sg13g2_decap_8 FILLER_12_856 ();
 sg13g2_decap_8 FILLER_12_863 ();
 sg13g2_decap_8 FILLER_12_870 ();
 sg13g2_decap_8 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_12_884 ();
 sg13g2_decap_8 FILLER_12_891 ();
 sg13g2_decap_8 FILLER_12_898 ();
 sg13g2_decap_8 FILLER_12_905 ();
 sg13g2_decap_8 FILLER_12_912 ();
 sg13g2_decap_8 FILLER_12_919 ();
 sg13g2_decap_8 FILLER_12_926 ();
 sg13g2_decap_8 FILLER_12_933 ();
 sg13g2_decap_8 FILLER_12_940 ();
 sg13g2_decap_8 FILLER_12_947 ();
 sg13g2_decap_8 FILLER_12_954 ();
 sg13g2_decap_8 FILLER_12_961 ();
 sg13g2_decap_8 FILLER_12_968 ();
 sg13g2_decap_8 FILLER_12_975 ();
 sg13g2_decap_8 FILLER_12_982 ();
 sg13g2_decap_8 FILLER_12_989 ();
 sg13g2_decap_8 FILLER_12_996 ();
 sg13g2_decap_8 FILLER_12_1003 ();
 sg13g2_decap_8 FILLER_12_1010 ();
 sg13g2_decap_8 FILLER_12_1017 ();
 sg13g2_decap_4 FILLER_12_1024 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_99 ();
 sg13g2_decap_8 FILLER_13_106 ();
 sg13g2_decap_8 FILLER_13_113 ();
 sg13g2_decap_8 FILLER_13_120 ();
 sg13g2_decap_8 FILLER_13_127 ();
 sg13g2_decap_4 FILLER_13_134 ();
 sg13g2_fill_2 FILLER_13_138 ();
 sg13g2_decap_8 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_174 ();
 sg13g2_decap_8 FILLER_13_181 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_195 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_decap_8 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_216 ();
 sg13g2_decap_8 FILLER_13_223 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_244 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_decap_8 FILLER_13_279 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_314 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_8 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_8 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_13_433 ();
 sg13g2_decap_8 FILLER_13_440 ();
 sg13g2_decap_8 FILLER_13_447 ();
 sg13g2_decap_8 FILLER_13_454 ();
 sg13g2_decap_8 FILLER_13_461 ();
 sg13g2_decap_8 FILLER_13_468 ();
 sg13g2_decap_8 FILLER_13_475 ();
 sg13g2_decap_8 FILLER_13_482 ();
 sg13g2_decap_8 FILLER_13_489 ();
 sg13g2_decap_8 FILLER_13_496 ();
 sg13g2_decap_8 FILLER_13_503 ();
 sg13g2_decap_8 FILLER_13_510 ();
 sg13g2_decap_8 FILLER_13_517 ();
 sg13g2_decap_8 FILLER_13_524 ();
 sg13g2_decap_8 FILLER_13_531 ();
 sg13g2_decap_8 FILLER_13_538 ();
 sg13g2_decap_8 FILLER_13_545 ();
 sg13g2_decap_8 FILLER_13_552 ();
 sg13g2_decap_8 FILLER_13_559 ();
 sg13g2_decap_8 FILLER_13_566 ();
 sg13g2_decap_8 FILLER_13_573 ();
 sg13g2_decap_8 FILLER_13_580 ();
 sg13g2_decap_8 FILLER_13_587 ();
 sg13g2_decap_8 FILLER_13_594 ();
 sg13g2_decap_8 FILLER_13_601 ();
 sg13g2_decap_8 FILLER_13_608 ();
 sg13g2_decap_8 FILLER_13_615 ();
 sg13g2_decap_8 FILLER_13_622 ();
 sg13g2_decap_8 FILLER_13_629 ();
 sg13g2_decap_8 FILLER_13_636 ();
 sg13g2_decap_8 FILLER_13_643 ();
 sg13g2_decap_8 FILLER_13_650 ();
 sg13g2_decap_8 FILLER_13_657 ();
 sg13g2_decap_8 FILLER_13_664 ();
 sg13g2_decap_8 FILLER_13_671 ();
 sg13g2_decap_8 FILLER_13_678 ();
 sg13g2_decap_8 FILLER_13_685 ();
 sg13g2_decap_8 FILLER_13_692 ();
 sg13g2_decap_8 FILLER_13_699 ();
 sg13g2_decap_8 FILLER_13_706 ();
 sg13g2_decap_8 FILLER_13_713 ();
 sg13g2_decap_8 FILLER_13_720 ();
 sg13g2_decap_8 FILLER_13_727 ();
 sg13g2_decap_8 FILLER_13_734 ();
 sg13g2_decap_8 FILLER_13_741 ();
 sg13g2_decap_8 FILLER_13_748 ();
 sg13g2_decap_8 FILLER_13_755 ();
 sg13g2_decap_8 FILLER_13_762 ();
 sg13g2_decap_8 FILLER_13_769 ();
 sg13g2_decap_8 FILLER_13_776 ();
 sg13g2_decap_8 FILLER_13_783 ();
 sg13g2_decap_8 FILLER_13_790 ();
 sg13g2_decap_8 FILLER_13_797 ();
 sg13g2_decap_8 FILLER_13_804 ();
 sg13g2_decap_8 FILLER_13_811 ();
 sg13g2_decap_8 FILLER_13_818 ();
 sg13g2_decap_8 FILLER_13_825 ();
 sg13g2_decap_8 FILLER_13_832 ();
 sg13g2_decap_8 FILLER_13_839 ();
 sg13g2_decap_8 FILLER_13_846 ();
 sg13g2_decap_8 FILLER_13_853 ();
 sg13g2_decap_8 FILLER_13_860 ();
 sg13g2_decap_8 FILLER_13_867 ();
 sg13g2_decap_8 FILLER_13_874 ();
 sg13g2_decap_8 FILLER_13_881 ();
 sg13g2_decap_8 FILLER_13_888 ();
 sg13g2_decap_8 FILLER_13_895 ();
 sg13g2_decap_8 FILLER_13_902 ();
 sg13g2_decap_8 FILLER_13_909 ();
 sg13g2_decap_8 FILLER_13_916 ();
 sg13g2_decap_8 FILLER_13_923 ();
 sg13g2_decap_8 FILLER_13_930 ();
 sg13g2_decap_8 FILLER_13_937 ();
 sg13g2_decap_8 FILLER_13_944 ();
 sg13g2_decap_8 FILLER_13_951 ();
 sg13g2_decap_8 FILLER_13_958 ();
 sg13g2_decap_8 FILLER_13_965 ();
 sg13g2_decap_8 FILLER_13_972 ();
 sg13g2_decap_8 FILLER_13_979 ();
 sg13g2_decap_8 FILLER_13_986 ();
 sg13g2_decap_8 FILLER_13_993 ();
 sg13g2_decap_8 FILLER_13_1000 ();
 sg13g2_decap_8 FILLER_13_1007 ();
 sg13g2_decap_8 FILLER_13_1014 ();
 sg13g2_decap_8 FILLER_13_1021 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_4 FILLER_14_11 ();
 sg13g2_fill_2 FILLER_14_15 ();
 sg13g2_decap_8 FILLER_14_43 ();
 sg13g2_decap_8 FILLER_14_50 ();
 sg13g2_decap_8 FILLER_14_57 ();
 sg13g2_decap_8 FILLER_14_64 ();
 sg13g2_decap_8 FILLER_14_71 ();
 sg13g2_decap_4 FILLER_14_78 ();
 sg13g2_decap_4 FILLER_14_90 ();
 sg13g2_decap_8 FILLER_14_108 ();
 sg13g2_decap_4 FILLER_14_115 ();
 sg13g2_decap_4 FILLER_14_128 ();
 sg13g2_fill_1 FILLER_14_132 ();
 sg13g2_decap_8 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_decap_8 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_decap_8 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_14_436 ();
 sg13g2_decap_8 FILLER_14_443 ();
 sg13g2_decap_8 FILLER_14_450 ();
 sg13g2_decap_8 FILLER_14_457 ();
 sg13g2_decap_8 FILLER_14_464 ();
 sg13g2_decap_8 FILLER_14_471 ();
 sg13g2_decap_8 FILLER_14_478 ();
 sg13g2_decap_8 FILLER_14_485 ();
 sg13g2_decap_8 FILLER_14_492 ();
 sg13g2_decap_8 FILLER_14_499 ();
 sg13g2_decap_8 FILLER_14_506 ();
 sg13g2_decap_8 FILLER_14_513 ();
 sg13g2_decap_8 FILLER_14_520 ();
 sg13g2_decap_8 FILLER_14_527 ();
 sg13g2_decap_8 FILLER_14_534 ();
 sg13g2_decap_8 FILLER_14_541 ();
 sg13g2_decap_8 FILLER_14_548 ();
 sg13g2_decap_8 FILLER_14_555 ();
 sg13g2_decap_8 FILLER_14_562 ();
 sg13g2_decap_8 FILLER_14_569 ();
 sg13g2_decap_8 FILLER_14_576 ();
 sg13g2_decap_8 FILLER_14_583 ();
 sg13g2_decap_8 FILLER_14_590 ();
 sg13g2_decap_8 FILLER_14_597 ();
 sg13g2_decap_8 FILLER_14_604 ();
 sg13g2_decap_8 FILLER_14_611 ();
 sg13g2_decap_8 FILLER_14_618 ();
 sg13g2_decap_8 FILLER_14_625 ();
 sg13g2_decap_8 FILLER_14_632 ();
 sg13g2_decap_8 FILLER_14_639 ();
 sg13g2_decap_8 FILLER_14_646 ();
 sg13g2_decap_8 FILLER_14_653 ();
 sg13g2_decap_8 FILLER_14_660 ();
 sg13g2_decap_8 FILLER_14_667 ();
 sg13g2_decap_8 FILLER_14_674 ();
 sg13g2_decap_8 FILLER_14_681 ();
 sg13g2_decap_8 FILLER_14_688 ();
 sg13g2_decap_8 FILLER_14_695 ();
 sg13g2_decap_8 FILLER_14_702 ();
 sg13g2_decap_8 FILLER_14_709 ();
 sg13g2_decap_8 FILLER_14_716 ();
 sg13g2_decap_8 FILLER_14_723 ();
 sg13g2_decap_8 FILLER_14_730 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_decap_8 FILLER_14_744 ();
 sg13g2_decap_8 FILLER_14_751 ();
 sg13g2_decap_8 FILLER_14_758 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_835 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_8 FILLER_14_849 ();
 sg13g2_decap_8 FILLER_14_856 ();
 sg13g2_decap_8 FILLER_14_863 ();
 sg13g2_decap_8 FILLER_14_870 ();
 sg13g2_decap_8 FILLER_14_877 ();
 sg13g2_decap_8 FILLER_14_884 ();
 sg13g2_decap_8 FILLER_14_891 ();
 sg13g2_decap_8 FILLER_14_898 ();
 sg13g2_decap_8 FILLER_14_905 ();
 sg13g2_decap_8 FILLER_14_912 ();
 sg13g2_decap_8 FILLER_14_919 ();
 sg13g2_decap_8 FILLER_14_926 ();
 sg13g2_decap_8 FILLER_14_933 ();
 sg13g2_decap_8 FILLER_14_940 ();
 sg13g2_decap_8 FILLER_14_947 ();
 sg13g2_decap_8 FILLER_14_954 ();
 sg13g2_decap_8 FILLER_14_961 ();
 sg13g2_decap_8 FILLER_14_968 ();
 sg13g2_decap_8 FILLER_14_975 ();
 sg13g2_decap_8 FILLER_14_982 ();
 sg13g2_decap_8 FILLER_14_989 ();
 sg13g2_decap_8 FILLER_14_996 ();
 sg13g2_decap_8 FILLER_14_1003 ();
 sg13g2_decap_8 FILLER_14_1010 ();
 sg13g2_decap_8 FILLER_14_1017 ();
 sg13g2_decap_4 FILLER_14_1024 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_183 ();
 sg13g2_decap_8 FILLER_15_190 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_decap_8 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_15_414 ();
 sg13g2_decap_8 FILLER_15_421 ();
 sg13g2_decap_8 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_15_435 ();
 sg13g2_decap_8 FILLER_15_442 ();
 sg13g2_decap_8 FILLER_15_449 ();
 sg13g2_decap_8 FILLER_15_456 ();
 sg13g2_decap_8 FILLER_15_463 ();
 sg13g2_decap_8 FILLER_15_470 ();
 sg13g2_decap_8 FILLER_15_477 ();
 sg13g2_decap_8 FILLER_15_484 ();
 sg13g2_decap_8 FILLER_15_491 ();
 sg13g2_decap_8 FILLER_15_498 ();
 sg13g2_decap_8 FILLER_15_505 ();
 sg13g2_decap_8 FILLER_15_512 ();
 sg13g2_decap_8 FILLER_15_519 ();
 sg13g2_decap_8 FILLER_15_526 ();
 sg13g2_decap_8 FILLER_15_533 ();
 sg13g2_decap_8 FILLER_15_540 ();
 sg13g2_decap_8 FILLER_15_547 ();
 sg13g2_decap_8 FILLER_15_554 ();
 sg13g2_decap_8 FILLER_15_561 ();
 sg13g2_decap_8 FILLER_15_568 ();
 sg13g2_decap_8 FILLER_15_575 ();
 sg13g2_decap_8 FILLER_15_582 ();
 sg13g2_decap_8 FILLER_15_589 ();
 sg13g2_decap_8 FILLER_15_596 ();
 sg13g2_decap_8 FILLER_15_603 ();
 sg13g2_decap_8 FILLER_15_610 ();
 sg13g2_decap_8 FILLER_15_617 ();
 sg13g2_decap_8 FILLER_15_624 ();
 sg13g2_decap_8 FILLER_15_631 ();
 sg13g2_decap_8 FILLER_15_638 ();
 sg13g2_decap_8 FILLER_15_645 ();
 sg13g2_decap_8 FILLER_15_652 ();
 sg13g2_decap_8 FILLER_15_659 ();
 sg13g2_decap_8 FILLER_15_666 ();
 sg13g2_decap_8 FILLER_15_673 ();
 sg13g2_decap_8 FILLER_15_680 ();
 sg13g2_decap_8 FILLER_15_687 ();
 sg13g2_decap_8 FILLER_15_694 ();
 sg13g2_decap_8 FILLER_15_701 ();
 sg13g2_decap_8 FILLER_15_708 ();
 sg13g2_decap_8 FILLER_15_715 ();
 sg13g2_decap_8 FILLER_15_722 ();
 sg13g2_decap_8 FILLER_15_729 ();
 sg13g2_decap_8 FILLER_15_736 ();
 sg13g2_decap_8 FILLER_15_743 ();
 sg13g2_decap_8 FILLER_15_750 ();
 sg13g2_decap_8 FILLER_15_757 ();
 sg13g2_decap_8 FILLER_15_764 ();
 sg13g2_decap_8 FILLER_15_771 ();
 sg13g2_decap_8 FILLER_15_778 ();
 sg13g2_decap_8 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_792 ();
 sg13g2_decap_8 FILLER_15_799 ();
 sg13g2_decap_8 FILLER_15_806 ();
 sg13g2_decap_8 FILLER_15_813 ();
 sg13g2_decap_8 FILLER_15_820 ();
 sg13g2_decap_8 FILLER_15_827 ();
 sg13g2_decap_8 FILLER_15_834 ();
 sg13g2_decap_8 FILLER_15_841 ();
 sg13g2_decap_8 FILLER_15_848 ();
 sg13g2_decap_8 FILLER_15_855 ();
 sg13g2_decap_8 FILLER_15_862 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_decap_8 FILLER_15_876 ();
 sg13g2_decap_8 FILLER_15_883 ();
 sg13g2_decap_8 FILLER_15_890 ();
 sg13g2_decap_8 FILLER_15_897 ();
 sg13g2_decap_8 FILLER_15_904 ();
 sg13g2_decap_8 FILLER_15_911 ();
 sg13g2_decap_8 FILLER_15_918 ();
 sg13g2_decap_8 FILLER_15_925 ();
 sg13g2_decap_8 FILLER_15_932 ();
 sg13g2_decap_8 FILLER_15_939 ();
 sg13g2_decap_8 FILLER_15_946 ();
 sg13g2_decap_8 FILLER_15_953 ();
 sg13g2_decap_8 FILLER_15_960 ();
 sg13g2_decap_8 FILLER_15_967 ();
 sg13g2_decap_8 FILLER_15_974 ();
 sg13g2_decap_8 FILLER_15_981 ();
 sg13g2_decap_8 FILLER_15_988 ();
 sg13g2_decap_8 FILLER_15_995 ();
 sg13g2_decap_8 FILLER_15_1002 ();
 sg13g2_decap_8 FILLER_15_1009 ();
 sg13g2_decap_8 FILLER_15_1016 ();
 sg13g2_decap_4 FILLER_15_1023 ();
 sg13g2_fill_2 FILLER_15_1027 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_4 FILLER_16_18 ();
 sg13g2_fill_2 FILLER_16_22 ();
 sg13g2_decap_8 FILLER_16_37 ();
 sg13g2_decap_8 FILLER_16_44 ();
 sg13g2_decap_8 FILLER_16_51 ();
 sg13g2_decap_8 FILLER_16_58 ();
 sg13g2_decap_8 FILLER_16_65 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_decap_8 FILLER_16_86 ();
 sg13g2_decap_4 FILLER_16_93 ();
 sg13g2_fill_2 FILLER_16_97 ();
 sg13g2_decap_8 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_decap_8 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_188 ();
 sg13g2_decap_8 FILLER_16_195 ();
 sg13g2_decap_8 FILLER_16_202 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_8 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_16_433 ();
 sg13g2_decap_8 FILLER_16_440 ();
 sg13g2_decap_8 FILLER_16_447 ();
 sg13g2_decap_8 FILLER_16_454 ();
 sg13g2_decap_8 FILLER_16_461 ();
 sg13g2_decap_8 FILLER_16_468 ();
 sg13g2_decap_8 FILLER_16_475 ();
 sg13g2_decap_8 FILLER_16_482 ();
 sg13g2_decap_8 FILLER_16_489 ();
 sg13g2_decap_8 FILLER_16_496 ();
 sg13g2_decap_8 FILLER_16_503 ();
 sg13g2_decap_8 FILLER_16_510 ();
 sg13g2_decap_8 FILLER_16_517 ();
 sg13g2_decap_8 FILLER_16_524 ();
 sg13g2_decap_8 FILLER_16_531 ();
 sg13g2_decap_8 FILLER_16_538 ();
 sg13g2_decap_8 FILLER_16_545 ();
 sg13g2_decap_8 FILLER_16_552 ();
 sg13g2_decap_8 FILLER_16_559 ();
 sg13g2_decap_8 FILLER_16_566 ();
 sg13g2_decap_8 FILLER_16_573 ();
 sg13g2_decap_8 FILLER_16_580 ();
 sg13g2_decap_8 FILLER_16_587 ();
 sg13g2_decap_8 FILLER_16_594 ();
 sg13g2_decap_8 FILLER_16_601 ();
 sg13g2_decap_8 FILLER_16_608 ();
 sg13g2_decap_8 FILLER_16_615 ();
 sg13g2_decap_8 FILLER_16_622 ();
 sg13g2_decap_8 FILLER_16_629 ();
 sg13g2_decap_8 FILLER_16_636 ();
 sg13g2_decap_8 FILLER_16_643 ();
 sg13g2_decap_8 FILLER_16_650 ();
 sg13g2_decap_8 FILLER_16_657 ();
 sg13g2_decap_8 FILLER_16_664 ();
 sg13g2_decap_8 FILLER_16_671 ();
 sg13g2_decap_8 FILLER_16_678 ();
 sg13g2_decap_8 FILLER_16_685 ();
 sg13g2_decap_8 FILLER_16_692 ();
 sg13g2_decap_8 FILLER_16_699 ();
 sg13g2_decap_8 FILLER_16_706 ();
 sg13g2_decap_8 FILLER_16_713 ();
 sg13g2_decap_8 FILLER_16_720 ();
 sg13g2_decap_8 FILLER_16_727 ();
 sg13g2_decap_8 FILLER_16_734 ();
 sg13g2_decap_8 FILLER_16_741 ();
 sg13g2_decap_8 FILLER_16_748 ();
 sg13g2_decap_8 FILLER_16_755 ();
 sg13g2_decap_8 FILLER_16_762 ();
 sg13g2_decap_8 FILLER_16_769 ();
 sg13g2_decap_8 FILLER_16_776 ();
 sg13g2_decap_8 FILLER_16_783 ();
 sg13g2_decap_8 FILLER_16_790 ();
 sg13g2_decap_8 FILLER_16_797 ();
 sg13g2_decap_8 FILLER_16_804 ();
 sg13g2_decap_8 FILLER_16_811 ();
 sg13g2_decap_8 FILLER_16_818 ();
 sg13g2_decap_8 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_832 ();
 sg13g2_decap_8 FILLER_16_839 ();
 sg13g2_decap_8 FILLER_16_846 ();
 sg13g2_decap_8 FILLER_16_853 ();
 sg13g2_decap_8 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_16_867 ();
 sg13g2_decap_8 FILLER_16_874 ();
 sg13g2_decap_8 FILLER_16_881 ();
 sg13g2_decap_8 FILLER_16_888 ();
 sg13g2_decap_8 FILLER_16_895 ();
 sg13g2_decap_8 FILLER_16_902 ();
 sg13g2_decap_8 FILLER_16_909 ();
 sg13g2_decap_8 FILLER_16_916 ();
 sg13g2_decap_8 FILLER_16_923 ();
 sg13g2_decap_8 FILLER_16_930 ();
 sg13g2_decap_8 FILLER_16_937 ();
 sg13g2_decap_8 FILLER_16_944 ();
 sg13g2_decap_8 FILLER_16_951 ();
 sg13g2_decap_8 FILLER_16_958 ();
 sg13g2_decap_8 FILLER_16_965 ();
 sg13g2_decap_8 FILLER_16_972 ();
 sg13g2_decap_8 FILLER_16_979 ();
 sg13g2_decap_8 FILLER_16_986 ();
 sg13g2_decap_8 FILLER_16_993 ();
 sg13g2_decap_8 FILLER_16_1000 ();
 sg13g2_decap_8 FILLER_16_1007 ();
 sg13g2_decap_8 FILLER_16_1014 ();
 sg13g2_decap_8 FILLER_16_1021 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_4 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_114 ();
 sg13g2_decap_8 FILLER_17_121 ();
 sg13g2_decap_4 FILLER_17_128 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_decap_8 FILLER_17_143 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_decap_8 FILLER_17_157 ();
 sg13g2_decap_8 FILLER_17_164 ();
 sg13g2_decap_8 FILLER_17_171 ();
 sg13g2_decap_8 FILLER_17_178 ();
 sg13g2_decap_8 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_192 ();
 sg13g2_decap_8 FILLER_17_199 ();
 sg13g2_decap_8 FILLER_17_206 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_220 ();
 sg13g2_decap_8 FILLER_17_227 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_262 ();
 sg13g2_decap_8 FILLER_17_269 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_17_409 ();
 sg13g2_decap_8 FILLER_17_416 ();
 sg13g2_decap_8 FILLER_17_423 ();
 sg13g2_decap_8 FILLER_17_430 ();
 sg13g2_decap_8 FILLER_17_437 ();
 sg13g2_decap_8 FILLER_17_444 ();
 sg13g2_decap_8 FILLER_17_451 ();
 sg13g2_decap_8 FILLER_17_458 ();
 sg13g2_decap_8 FILLER_17_465 ();
 sg13g2_decap_8 FILLER_17_472 ();
 sg13g2_decap_8 FILLER_17_479 ();
 sg13g2_decap_8 FILLER_17_486 ();
 sg13g2_decap_8 FILLER_17_493 ();
 sg13g2_decap_8 FILLER_17_500 ();
 sg13g2_decap_8 FILLER_17_507 ();
 sg13g2_decap_8 FILLER_17_514 ();
 sg13g2_decap_8 FILLER_17_521 ();
 sg13g2_decap_8 FILLER_17_528 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_decap_8 FILLER_17_542 ();
 sg13g2_decap_8 FILLER_17_549 ();
 sg13g2_decap_8 FILLER_17_556 ();
 sg13g2_decap_8 FILLER_17_563 ();
 sg13g2_decap_8 FILLER_17_570 ();
 sg13g2_decap_8 FILLER_17_577 ();
 sg13g2_decap_8 FILLER_17_584 ();
 sg13g2_decap_8 FILLER_17_591 ();
 sg13g2_decap_8 FILLER_17_598 ();
 sg13g2_decap_8 FILLER_17_605 ();
 sg13g2_decap_8 FILLER_17_612 ();
 sg13g2_decap_8 FILLER_17_619 ();
 sg13g2_decap_8 FILLER_17_626 ();
 sg13g2_decap_8 FILLER_17_633 ();
 sg13g2_decap_8 FILLER_17_640 ();
 sg13g2_decap_8 FILLER_17_647 ();
 sg13g2_decap_8 FILLER_17_654 ();
 sg13g2_decap_8 FILLER_17_661 ();
 sg13g2_decap_8 FILLER_17_668 ();
 sg13g2_decap_8 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_682 ();
 sg13g2_decap_8 FILLER_17_689 ();
 sg13g2_decap_8 FILLER_17_696 ();
 sg13g2_decap_8 FILLER_17_703 ();
 sg13g2_decap_8 FILLER_17_710 ();
 sg13g2_decap_8 FILLER_17_717 ();
 sg13g2_decap_8 FILLER_17_724 ();
 sg13g2_decap_8 FILLER_17_731 ();
 sg13g2_decap_8 FILLER_17_738 ();
 sg13g2_decap_8 FILLER_17_745 ();
 sg13g2_decap_8 FILLER_17_752 ();
 sg13g2_decap_8 FILLER_17_759 ();
 sg13g2_decap_8 FILLER_17_766 ();
 sg13g2_decap_8 FILLER_17_773 ();
 sg13g2_decap_8 FILLER_17_780 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_decap_8 FILLER_17_794 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_decap_8 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_decap_8 FILLER_17_836 ();
 sg13g2_decap_8 FILLER_17_843 ();
 sg13g2_decap_8 FILLER_17_850 ();
 sg13g2_decap_8 FILLER_17_857 ();
 sg13g2_decap_8 FILLER_17_864 ();
 sg13g2_decap_8 FILLER_17_871 ();
 sg13g2_decap_8 FILLER_17_878 ();
 sg13g2_decap_8 FILLER_17_885 ();
 sg13g2_decap_8 FILLER_17_892 ();
 sg13g2_decap_8 FILLER_17_899 ();
 sg13g2_decap_8 FILLER_17_906 ();
 sg13g2_decap_8 FILLER_17_913 ();
 sg13g2_decap_8 FILLER_17_920 ();
 sg13g2_decap_8 FILLER_17_927 ();
 sg13g2_decap_8 FILLER_17_934 ();
 sg13g2_decap_8 FILLER_17_941 ();
 sg13g2_decap_8 FILLER_17_948 ();
 sg13g2_decap_8 FILLER_17_955 ();
 sg13g2_decap_8 FILLER_17_962 ();
 sg13g2_decap_8 FILLER_17_969 ();
 sg13g2_decap_8 FILLER_17_976 ();
 sg13g2_decap_8 FILLER_17_983 ();
 sg13g2_decap_8 FILLER_17_990 ();
 sg13g2_decap_8 FILLER_17_997 ();
 sg13g2_decap_8 FILLER_17_1004 ();
 sg13g2_decap_8 FILLER_17_1011 ();
 sg13g2_decap_8 FILLER_17_1018 ();
 sg13g2_decap_4 FILLER_17_1025 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_213 ();
 sg13g2_decap_8 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_227 ();
 sg13g2_decap_8 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_decap_8 FILLER_18_430 ();
 sg13g2_decap_8 FILLER_18_437 ();
 sg13g2_decap_8 FILLER_18_444 ();
 sg13g2_decap_8 FILLER_18_451 ();
 sg13g2_decap_8 FILLER_18_458 ();
 sg13g2_decap_8 FILLER_18_465 ();
 sg13g2_decap_8 FILLER_18_472 ();
 sg13g2_decap_8 FILLER_18_479 ();
 sg13g2_decap_8 FILLER_18_486 ();
 sg13g2_decap_8 FILLER_18_493 ();
 sg13g2_decap_8 FILLER_18_500 ();
 sg13g2_decap_8 FILLER_18_507 ();
 sg13g2_decap_8 FILLER_18_514 ();
 sg13g2_decap_8 FILLER_18_521 ();
 sg13g2_decap_8 FILLER_18_528 ();
 sg13g2_decap_8 FILLER_18_535 ();
 sg13g2_decap_8 FILLER_18_542 ();
 sg13g2_decap_8 FILLER_18_549 ();
 sg13g2_decap_8 FILLER_18_556 ();
 sg13g2_decap_8 FILLER_18_563 ();
 sg13g2_decap_8 FILLER_18_570 ();
 sg13g2_decap_8 FILLER_18_577 ();
 sg13g2_decap_8 FILLER_18_584 ();
 sg13g2_decap_8 FILLER_18_591 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_decap_8 FILLER_18_605 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_decap_8 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_8 FILLER_18_640 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_8 FILLER_18_654 ();
 sg13g2_decap_8 FILLER_18_661 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_decap_8 FILLER_18_675 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_decap_8 FILLER_18_689 ();
 sg13g2_decap_8 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_8 FILLER_18_857 ();
 sg13g2_decap_8 FILLER_18_864 ();
 sg13g2_decap_8 FILLER_18_871 ();
 sg13g2_decap_8 FILLER_18_878 ();
 sg13g2_decap_8 FILLER_18_885 ();
 sg13g2_decap_8 FILLER_18_892 ();
 sg13g2_decap_8 FILLER_18_899 ();
 sg13g2_decap_8 FILLER_18_906 ();
 sg13g2_decap_8 FILLER_18_913 ();
 sg13g2_decap_8 FILLER_18_920 ();
 sg13g2_decap_8 FILLER_18_927 ();
 sg13g2_decap_8 FILLER_18_934 ();
 sg13g2_decap_8 FILLER_18_941 ();
 sg13g2_decap_8 FILLER_18_948 ();
 sg13g2_decap_8 FILLER_18_955 ();
 sg13g2_decap_8 FILLER_18_962 ();
 sg13g2_decap_8 FILLER_18_969 ();
 sg13g2_decap_8 FILLER_18_976 ();
 sg13g2_decap_8 FILLER_18_983 ();
 sg13g2_decap_8 FILLER_18_990 ();
 sg13g2_decap_8 FILLER_18_997 ();
 sg13g2_decap_8 FILLER_18_1004 ();
 sg13g2_decap_8 FILLER_18_1011 ();
 sg13g2_decap_8 FILLER_18_1018 ();
 sg13g2_decap_4 FILLER_18_1025 ();
 sg13g2_decap_8 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_4 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_decap_8 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_decap_8 FILLER_19_139 ();
 sg13g2_decap_8 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_decap_8 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_19_412 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_8 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_19_433 ();
 sg13g2_decap_8 FILLER_19_440 ();
 sg13g2_decap_8 FILLER_19_447 ();
 sg13g2_decap_8 FILLER_19_454 ();
 sg13g2_decap_8 FILLER_19_461 ();
 sg13g2_decap_8 FILLER_19_468 ();
 sg13g2_decap_8 FILLER_19_475 ();
 sg13g2_decap_8 FILLER_19_482 ();
 sg13g2_decap_8 FILLER_19_489 ();
 sg13g2_decap_8 FILLER_19_496 ();
 sg13g2_decap_8 FILLER_19_503 ();
 sg13g2_decap_8 FILLER_19_510 ();
 sg13g2_decap_8 FILLER_19_517 ();
 sg13g2_decap_8 FILLER_19_524 ();
 sg13g2_decap_8 FILLER_19_531 ();
 sg13g2_decap_8 FILLER_19_538 ();
 sg13g2_decap_8 FILLER_19_545 ();
 sg13g2_decap_8 FILLER_19_552 ();
 sg13g2_decap_8 FILLER_19_559 ();
 sg13g2_decap_8 FILLER_19_566 ();
 sg13g2_decap_8 FILLER_19_573 ();
 sg13g2_decap_8 FILLER_19_580 ();
 sg13g2_decap_8 FILLER_19_587 ();
 sg13g2_decap_8 FILLER_19_594 ();
 sg13g2_decap_8 FILLER_19_601 ();
 sg13g2_decap_8 FILLER_19_608 ();
 sg13g2_decap_8 FILLER_19_615 ();
 sg13g2_decap_8 FILLER_19_622 ();
 sg13g2_decap_8 FILLER_19_629 ();
 sg13g2_decap_8 FILLER_19_636 ();
 sg13g2_decap_8 FILLER_19_643 ();
 sg13g2_decap_8 FILLER_19_650 ();
 sg13g2_decap_8 FILLER_19_657 ();
 sg13g2_decap_8 FILLER_19_664 ();
 sg13g2_decap_8 FILLER_19_671 ();
 sg13g2_decap_8 FILLER_19_678 ();
 sg13g2_decap_8 FILLER_19_685 ();
 sg13g2_decap_8 FILLER_19_692 ();
 sg13g2_decap_8 FILLER_19_699 ();
 sg13g2_decap_8 FILLER_19_706 ();
 sg13g2_decap_8 FILLER_19_713 ();
 sg13g2_decap_8 FILLER_19_720 ();
 sg13g2_decap_8 FILLER_19_727 ();
 sg13g2_decap_8 FILLER_19_734 ();
 sg13g2_decap_8 FILLER_19_741 ();
 sg13g2_decap_8 FILLER_19_748 ();
 sg13g2_decap_8 FILLER_19_755 ();
 sg13g2_decap_8 FILLER_19_762 ();
 sg13g2_decap_8 FILLER_19_769 ();
 sg13g2_decap_8 FILLER_19_776 ();
 sg13g2_decap_8 FILLER_19_783 ();
 sg13g2_decap_8 FILLER_19_790 ();
 sg13g2_decap_8 FILLER_19_797 ();
 sg13g2_decap_8 FILLER_19_804 ();
 sg13g2_decap_8 FILLER_19_811 ();
 sg13g2_decap_8 FILLER_19_818 ();
 sg13g2_decap_8 FILLER_19_825 ();
 sg13g2_decap_8 FILLER_19_832 ();
 sg13g2_decap_8 FILLER_19_839 ();
 sg13g2_decap_8 FILLER_19_846 ();
 sg13g2_decap_8 FILLER_19_853 ();
 sg13g2_decap_8 FILLER_19_860 ();
 sg13g2_decap_8 FILLER_19_867 ();
 sg13g2_decap_8 FILLER_19_874 ();
 sg13g2_decap_8 FILLER_19_881 ();
 sg13g2_decap_8 FILLER_19_888 ();
 sg13g2_decap_8 FILLER_19_895 ();
 sg13g2_decap_8 FILLER_19_902 ();
 sg13g2_decap_8 FILLER_19_909 ();
 sg13g2_decap_8 FILLER_19_916 ();
 sg13g2_decap_8 FILLER_19_923 ();
 sg13g2_decap_8 FILLER_19_930 ();
 sg13g2_decap_8 FILLER_19_937 ();
 sg13g2_decap_8 FILLER_19_944 ();
 sg13g2_decap_8 FILLER_19_951 ();
 sg13g2_decap_8 FILLER_19_958 ();
 sg13g2_decap_8 FILLER_19_965 ();
 sg13g2_decap_8 FILLER_19_972 ();
 sg13g2_decap_8 FILLER_19_979 ();
 sg13g2_decap_8 FILLER_19_986 ();
 sg13g2_decap_8 FILLER_19_993 ();
 sg13g2_decap_8 FILLER_19_1000 ();
 sg13g2_decap_8 FILLER_19_1007 ();
 sg13g2_decap_8 FILLER_19_1014 ();
 sg13g2_decap_8 FILLER_19_1021 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_decap_8 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_20_868 ();
 sg13g2_decap_8 FILLER_20_875 ();
 sg13g2_decap_8 FILLER_20_882 ();
 sg13g2_decap_8 FILLER_20_889 ();
 sg13g2_decap_8 FILLER_20_896 ();
 sg13g2_decap_8 FILLER_20_903 ();
 sg13g2_decap_8 FILLER_20_910 ();
 sg13g2_decap_8 FILLER_20_917 ();
 sg13g2_decap_8 FILLER_20_924 ();
 sg13g2_decap_8 FILLER_20_931 ();
 sg13g2_decap_8 FILLER_20_938 ();
 sg13g2_decap_8 FILLER_20_945 ();
 sg13g2_decap_8 FILLER_20_952 ();
 sg13g2_decap_8 FILLER_20_959 ();
 sg13g2_decap_8 FILLER_20_966 ();
 sg13g2_decap_8 FILLER_20_973 ();
 sg13g2_decap_8 FILLER_20_980 ();
 sg13g2_decap_8 FILLER_20_987 ();
 sg13g2_decap_8 FILLER_20_994 ();
 sg13g2_decap_8 FILLER_20_1001 ();
 sg13g2_decap_8 FILLER_20_1008 ();
 sg13g2_decap_8 FILLER_20_1015 ();
 sg13g2_decap_8 FILLER_20_1022 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_4 FILLER_21_87 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_101 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_decap_8 FILLER_21_115 ();
 sg13g2_decap_8 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_185 ();
 sg13g2_decap_8 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_decap_8 FILLER_21_227 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_decap_8 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_283 ();
 sg13g2_decap_8 FILLER_21_290 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_416 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_21_430 ();
 sg13g2_decap_8 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_444 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_decap_8 FILLER_21_458 ();
 sg13g2_decap_8 FILLER_21_465 ();
 sg13g2_decap_8 FILLER_21_472 ();
 sg13g2_decap_8 FILLER_21_479 ();
 sg13g2_decap_8 FILLER_21_486 ();
 sg13g2_decap_8 FILLER_21_493 ();
 sg13g2_decap_8 FILLER_21_500 ();
 sg13g2_decap_8 FILLER_21_507 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_decap_8 FILLER_21_521 ();
 sg13g2_decap_8 FILLER_21_528 ();
 sg13g2_decap_8 FILLER_21_535 ();
 sg13g2_decap_8 FILLER_21_542 ();
 sg13g2_decap_8 FILLER_21_549 ();
 sg13g2_decap_8 FILLER_21_556 ();
 sg13g2_decap_8 FILLER_21_563 ();
 sg13g2_decap_8 FILLER_21_570 ();
 sg13g2_decap_8 FILLER_21_577 ();
 sg13g2_decap_8 FILLER_21_584 ();
 sg13g2_decap_8 FILLER_21_591 ();
 sg13g2_decap_8 FILLER_21_598 ();
 sg13g2_decap_8 FILLER_21_605 ();
 sg13g2_decap_8 FILLER_21_612 ();
 sg13g2_decap_8 FILLER_21_619 ();
 sg13g2_decap_8 FILLER_21_626 ();
 sg13g2_decap_8 FILLER_21_633 ();
 sg13g2_decap_8 FILLER_21_640 ();
 sg13g2_decap_8 FILLER_21_647 ();
 sg13g2_decap_8 FILLER_21_654 ();
 sg13g2_decap_8 FILLER_21_661 ();
 sg13g2_decap_8 FILLER_21_668 ();
 sg13g2_decap_8 FILLER_21_675 ();
 sg13g2_decap_8 FILLER_21_682 ();
 sg13g2_decap_8 FILLER_21_689 ();
 sg13g2_decap_8 FILLER_21_696 ();
 sg13g2_decap_8 FILLER_21_703 ();
 sg13g2_decap_8 FILLER_21_710 ();
 sg13g2_decap_8 FILLER_21_717 ();
 sg13g2_decap_8 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_731 ();
 sg13g2_decap_8 FILLER_21_738 ();
 sg13g2_decap_8 FILLER_21_745 ();
 sg13g2_decap_8 FILLER_21_752 ();
 sg13g2_decap_8 FILLER_21_759 ();
 sg13g2_decap_8 FILLER_21_766 ();
 sg13g2_decap_8 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_780 ();
 sg13g2_decap_8 FILLER_21_787 ();
 sg13g2_decap_8 FILLER_21_794 ();
 sg13g2_decap_8 FILLER_21_801 ();
 sg13g2_decap_8 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_815 ();
 sg13g2_decap_8 FILLER_21_822 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_decap_8 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_850 ();
 sg13g2_decap_8 FILLER_21_857 ();
 sg13g2_decap_8 FILLER_21_864 ();
 sg13g2_decap_8 FILLER_21_871 ();
 sg13g2_decap_8 FILLER_21_878 ();
 sg13g2_decap_8 FILLER_21_885 ();
 sg13g2_decap_8 FILLER_21_892 ();
 sg13g2_decap_8 FILLER_21_899 ();
 sg13g2_decap_8 FILLER_21_906 ();
 sg13g2_decap_8 FILLER_21_913 ();
 sg13g2_decap_8 FILLER_21_920 ();
 sg13g2_decap_8 FILLER_21_927 ();
 sg13g2_decap_8 FILLER_21_934 ();
 sg13g2_decap_8 FILLER_21_941 ();
 sg13g2_decap_8 FILLER_21_948 ();
 sg13g2_decap_8 FILLER_21_955 ();
 sg13g2_decap_8 FILLER_21_962 ();
 sg13g2_decap_8 FILLER_21_969 ();
 sg13g2_decap_8 FILLER_21_976 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_decap_8 FILLER_21_990 ();
 sg13g2_decap_8 FILLER_21_997 ();
 sg13g2_decap_8 FILLER_21_1004 ();
 sg13g2_decap_8 FILLER_21_1011 ();
 sg13g2_decap_8 FILLER_21_1018 ();
 sg13g2_decap_4 FILLER_21_1025 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_decap_4 FILLER_22_67 ();
 sg13g2_fill_2 FILLER_22_71 ();
 sg13g2_decap_8 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_107 ();
 sg13g2_decap_8 FILLER_22_114 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_decap_8 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_149 ();
 sg13g2_decap_8 FILLER_22_156 ();
 sg13g2_decap_8 FILLER_22_163 ();
 sg13g2_decap_8 FILLER_22_170 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_decap_8 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_decap_8 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_decap_8 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_decap_8 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_22_436 ();
 sg13g2_decap_8 FILLER_22_443 ();
 sg13g2_decap_8 FILLER_22_450 ();
 sg13g2_decap_8 FILLER_22_457 ();
 sg13g2_decap_8 FILLER_22_464 ();
 sg13g2_decap_8 FILLER_22_471 ();
 sg13g2_decap_8 FILLER_22_478 ();
 sg13g2_decap_8 FILLER_22_485 ();
 sg13g2_decap_8 FILLER_22_492 ();
 sg13g2_decap_8 FILLER_22_499 ();
 sg13g2_decap_8 FILLER_22_506 ();
 sg13g2_decap_8 FILLER_22_513 ();
 sg13g2_decap_8 FILLER_22_520 ();
 sg13g2_decap_8 FILLER_22_527 ();
 sg13g2_decap_8 FILLER_22_534 ();
 sg13g2_decap_8 FILLER_22_541 ();
 sg13g2_decap_8 FILLER_22_548 ();
 sg13g2_decap_8 FILLER_22_555 ();
 sg13g2_decap_8 FILLER_22_562 ();
 sg13g2_decap_8 FILLER_22_569 ();
 sg13g2_decap_8 FILLER_22_576 ();
 sg13g2_decap_8 FILLER_22_583 ();
 sg13g2_decap_8 FILLER_22_590 ();
 sg13g2_decap_8 FILLER_22_597 ();
 sg13g2_decap_8 FILLER_22_604 ();
 sg13g2_decap_8 FILLER_22_611 ();
 sg13g2_decap_8 FILLER_22_618 ();
 sg13g2_decap_8 FILLER_22_625 ();
 sg13g2_decap_8 FILLER_22_632 ();
 sg13g2_decap_8 FILLER_22_639 ();
 sg13g2_decap_8 FILLER_22_646 ();
 sg13g2_decap_8 FILLER_22_653 ();
 sg13g2_decap_8 FILLER_22_660 ();
 sg13g2_decap_8 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_674 ();
 sg13g2_decap_8 FILLER_22_681 ();
 sg13g2_decap_8 FILLER_22_688 ();
 sg13g2_decap_8 FILLER_22_695 ();
 sg13g2_decap_8 FILLER_22_702 ();
 sg13g2_decap_8 FILLER_22_709 ();
 sg13g2_decap_8 FILLER_22_716 ();
 sg13g2_decap_8 FILLER_22_723 ();
 sg13g2_decap_8 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_744 ();
 sg13g2_decap_8 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_758 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_decap_8 FILLER_22_779 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_793 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_decap_8 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_842 ();
 sg13g2_decap_8 FILLER_22_849 ();
 sg13g2_decap_8 FILLER_22_856 ();
 sg13g2_decap_8 FILLER_22_863 ();
 sg13g2_decap_8 FILLER_22_870 ();
 sg13g2_decap_8 FILLER_22_877 ();
 sg13g2_decap_8 FILLER_22_884 ();
 sg13g2_decap_8 FILLER_22_891 ();
 sg13g2_decap_8 FILLER_22_898 ();
 sg13g2_decap_8 FILLER_22_905 ();
 sg13g2_decap_8 FILLER_22_912 ();
 sg13g2_decap_8 FILLER_22_919 ();
 sg13g2_decap_8 FILLER_22_926 ();
 sg13g2_decap_8 FILLER_22_933 ();
 sg13g2_decap_8 FILLER_22_940 ();
 sg13g2_decap_8 FILLER_22_947 ();
 sg13g2_decap_8 FILLER_22_954 ();
 sg13g2_decap_8 FILLER_22_961 ();
 sg13g2_decap_8 FILLER_22_968 ();
 sg13g2_decap_8 FILLER_22_975 ();
 sg13g2_decap_8 FILLER_22_982 ();
 sg13g2_decap_8 FILLER_22_989 ();
 sg13g2_decap_8 FILLER_22_996 ();
 sg13g2_decap_8 FILLER_22_1003 ();
 sg13g2_decap_8 FILLER_22_1010 ();
 sg13g2_decap_8 FILLER_22_1017 ();
 sg13g2_decap_4 FILLER_22_1024 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_81 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_decap_8 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_473 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_decap_8 FILLER_23_508 ();
 sg13g2_decap_8 FILLER_23_515 ();
 sg13g2_decap_8 FILLER_23_522 ();
 sg13g2_decap_8 FILLER_23_529 ();
 sg13g2_decap_8 FILLER_23_536 ();
 sg13g2_decap_8 FILLER_23_543 ();
 sg13g2_decap_8 FILLER_23_550 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_decap_8 FILLER_23_564 ();
 sg13g2_decap_8 FILLER_23_571 ();
 sg13g2_decap_8 FILLER_23_578 ();
 sg13g2_decap_8 FILLER_23_585 ();
 sg13g2_decap_8 FILLER_23_592 ();
 sg13g2_decap_8 FILLER_23_599 ();
 sg13g2_decap_8 FILLER_23_606 ();
 sg13g2_decap_8 FILLER_23_613 ();
 sg13g2_decap_8 FILLER_23_620 ();
 sg13g2_decap_8 FILLER_23_627 ();
 sg13g2_decap_8 FILLER_23_634 ();
 sg13g2_decap_8 FILLER_23_641 ();
 sg13g2_decap_8 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_655 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_decap_8 FILLER_23_718 ();
 sg13g2_decap_8 FILLER_23_725 ();
 sg13g2_decap_8 FILLER_23_732 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_decap_8 FILLER_23_753 ();
 sg13g2_decap_8 FILLER_23_760 ();
 sg13g2_decap_8 FILLER_23_767 ();
 sg13g2_decap_8 FILLER_23_774 ();
 sg13g2_decap_8 FILLER_23_781 ();
 sg13g2_decap_8 FILLER_23_788 ();
 sg13g2_decap_8 FILLER_23_795 ();
 sg13g2_decap_8 FILLER_23_802 ();
 sg13g2_decap_8 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_816 ();
 sg13g2_decap_8 FILLER_23_823 ();
 sg13g2_decap_8 FILLER_23_830 ();
 sg13g2_decap_8 FILLER_23_837 ();
 sg13g2_decap_8 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_851 ();
 sg13g2_decap_8 FILLER_23_858 ();
 sg13g2_decap_8 FILLER_23_865 ();
 sg13g2_decap_8 FILLER_23_872 ();
 sg13g2_decap_8 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_886 ();
 sg13g2_decap_8 FILLER_23_893 ();
 sg13g2_decap_8 FILLER_23_900 ();
 sg13g2_decap_8 FILLER_23_907 ();
 sg13g2_decap_8 FILLER_23_914 ();
 sg13g2_decap_8 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_23_928 ();
 sg13g2_decap_8 FILLER_23_935 ();
 sg13g2_decap_8 FILLER_23_942 ();
 sg13g2_decap_8 FILLER_23_949 ();
 sg13g2_decap_8 FILLER_23_956 ();
 sg13g2_decap_8 FILLER_23_963 ();
 sg13g2_decap_8 FILLER_23_970 ();
 sg13g2_decap_8 FILLER_23_977 ();
 sg13g2_decap_8 FILLER_23_984 ();
 sg13g2_decap_8 FILLER_23_991 ();
 sg13g2_decap_8 FILLER_23_998 ();
 sg13g2_decap_8 FILLER_23_1005 ();
 sg13g2_decap_8 FILLER_23_1012 ();
 sg13g2_decap_8 FILLER_23_1019 ();
 sg13g2_fill_2 FILLER_23_1026 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_424 ();
 sg13g2_decap_8 FILLER_24_431 ();
 sg13g2_decap_8 FILLER_24_438 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_473 ();
 sg13g2_decap_8 FILLER_24_480 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_decap_8 FILLER_24_508 ();
 sg13g2_decap_8 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_522 ();
 sg13g2_decap_8 FILLER_24_529 ();
 sg13g2_decap_8 FILLER_24_536 ();
 sg13g2_decap_8 FILLER_24_543 ();
 sg13g2_decap_8 FILLER_24_550 ();
 sg13g2_decap_8 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_8 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_decap_8 FILLER_24_599 ();
 sg13g2_decap_8 FILLER_24_606 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_decap_8 FILLER_24_620 ();
 sg13g2_decap_8 FILLER_24_627 ();
 sg13g2_decap_8 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_641 ();
 sg13g2_decap_8 FILLER_24_648 ();
 sg13g2_decap_8 FILLER_24_655 ();
 sg13g2_decap_8 FILLER_24_662 ();
 sg13g2_decap_8 FILLER_24_669 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_690 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_704 ();
 sg13g2_decap_8 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_718 ();
 sg13g2_decap_8 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_8 FILLER_24_746 ();
 sg13g2_decap_8 FILLER_24_753 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_decap_8 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_decap_8 FILLER_24_788 ();
 sg13g2_decap_8 FILLER_24_795 ();
 sg13g2_decap_8 FILLER_24_802 ();
 sg13g2_decap_8 FILLER_24_809 ();
 sg13g2_decap_8 FILLER_24_816 ();
 sg13g2_decap_8 FILLER_24_823 ();
 sg13g2_decap_8 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_837 ();
 sg13g2_decap_8 FILLER_24_844 ();
 sg13g2_decap_8 FILLER_24_851 ();
 sg13g2_decap_8 FILLER_24_858 ();
 sg13g2_decap_8 FILLER_24_865 ();
 sg13g2_decap_8 FILLER_24_872 ();
 sg13g2_decap_8 FILLER_24_879 ();
 sg13g2_decap_8 FILLER_24_886 ();
 sg13g2_decap_8 FILLER_24_893 ();
 sg13g2_decap_8 FILLER_24_900 ();
 sg13g2_decap_8 FILLER_24_907 ();
 sg13g2_decap_8 FILLER_24_914 ();
 sg13g2_decap_8 FILLER_24_921 ();
 sg13g2_decap_8 FILLER_24_928 ();
 sg13g2_decap_8 FILLER_24_935 ();
 sg13g2_decap_8 FILLER_24_942 ();
 sg13g2_decap_8 FILLER_24_949 ();
 sg13g2_decap_8 FILLER_24_956 ();
 sg13g2_decap_8 FILLER_24_963 ();
 sg13g2_decap_8 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_decap_8 FILLER_24_984 ();
 sg13g2_decap_8 FILLER_24_991 ();
 sg13g2_decap_8 FILLER_24_998 ();
 sg13g2_decap_8 FILLER_24_1005 ();
 sg13g2_decap_8 FILLER_24_1012 ();
 sg13g2_decap_8 FILLER_24_1019 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_74 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_179 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_424 ();
 sg13g2_decap_8 FILLER_25_431 ();
 sg13g2_decap_8 FILLER_25_438 ();
 sg13g2_decap_8 FILLER_25_445 ();
 sg13g2_decap_8 FILLER_25_452 ();
 sg13g2_decap_8 FILLER_25_459 ();
 sg13g2_decap_8 FILLER_25_466 ();
 sg13g2_decap_8 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_480 ();
 sg13g2_decap_8 FILLER_25_487 ();
 sg13g2_decap_8 FILLER_25_494 ();
 sg13g2_decap_8 FILLER_25_501 ();
 sg13g2_decap_8 FILLER_25_508 ();
 sg13g2_decap_8 FILLER_25_515 ();
 sg13g2_decap_8 FILLER_25_522 ();
 sg13g2_decap_8 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_decap_8 FILLER_25_564 ();
 sg13g2_decap_8 FILLER_25_571 ();
 sg13g2_decap_8 FILLER_25_578 ();
 sg13g2_decap_8 FILLER_25_585 ();
 sg13g2_decap_8 FILLER_25_592 ();
 sg13g2_decap_8 FILLER_25_599 ();
 sg13g2_decap_8 FILLER_25_606 ();
 sg13g2_decap_8 FILLER_25_613 ();
 sg13g2_decap_8 FILLER_25_620 ();
 sg13g2_decap_8 FILLER_25_627 ();
 sg13g2_decap_8 FILLER_25_634 ();
 sg13g2_decap_8 FILLER_25_641 ();
 sg13g2_decap_8 FILLER_25_648 ();
 sg13g2_decap_8 FILLER_25_655 ();
 sg13g2_decap_8 FILLER_25_662 ();
 sg13g2_decap_8 FILLER_25_669 ();
 sg13g2_decap_8 FILLER_25_676 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_8 FILLER_25_690 ();
 sg13g2_decap_8 FILLER_25_697 ();
 sg13g2_decap_8 FILLER_25_704 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_8 FILLER_25_718 ();
 sg13g2_decap_8 FILLER_25_725 ();
 sg13g2_decap_8 FILLER_25_732 ();
 sg13g2_decap_8 FILLER_25_739 ();
 sg13g2_decap_8 FILLER_25_746 ();
 sg13g2_decap_8 FILLER_25_753 ();
 sg13g2_decap_8 FILLER_25_760 ();
 sg13g2_decap_8 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_774 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_8 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_8 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_8 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_25_865 ();
 sg13g2_decap_8 FILLER_25_872 ();
 sg13g2_decap_8 FILLER_25_879 ();
 sg13g2_decap_8 FILLER_25_886 ();
 sg13g2_decap_8 FILLER_25_893 ();
 sg13g2_decap_8 FILLER_25_900 ();
 sg13g2_decap_8 FILLER_25_907 ();
 sg13g2_decap_8 FILLER_25_914 ();
 sg13g2_decap_8 FILLER_25_921 ();
 sg13g2_decap_8 FILLER_25_928 ();
 sg13g2_decap_8 FILLER_25_935 ();
 sg13g2_decap_8 FILLER_25_942 ();
 sg13g2_decap_8 FILLER_25_949 ();
 sg13g2_decap_8 FILLER_25_956 ();
 sg13g2_decap_8 FILLER_25_963 ();
 sg13g2_decap_8 FILLER_25_970 ();
 sg13g2_decap_8 FILLER_25_977 ();
 sg13g2_decap_8 FILLER_25_984 ();
 sg13g2_decap_8 FILLER_25_991 ();
 sg13g2_decap_8 FILLER_25_998 ();
 sg13g2_decap_8 FILLER_25_1005 ();
 sg13g2_decap_8 FILLER_25_1012 ();
 sg13g2_decap_8 FILLER_25_1019 ();
 sg13g2_fill_2 FILLER_25_1026 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_fill_2 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_8 FILLER_26_424 ();
 sg13g2_decap_8 FILLER_26_431 ();
 sg13g2_decap_8 FILLER_26_438 ();
 sg13g2_decap_8 FILLER_26_445 ();
 sg13g2_decap_8 FILLER_26_452 ();
 sg13g2_decap_8 FILLER_26_459 ();
 sg13g2_decap_8 FILLER_26_466 ();
 sg13g2_decap_8 FILLER_26_473 ();
 sg13g2_decap_8 FILLER_26_480 ();
 sg13g2_decap_8 FILLER_26_487 ();
 sg13g2_decap_8 FILLER_26_494 ();
 sg13g2_decap_8 FILLER_26_501 ();
 sg13g2_decap_8 FILLER_26_508 ();
 sg13g2_decap_8 FILLER_26_515 ();
 sg13g2_decap_8 FILLER_26_522 ();
 sg13g2_decap_8 FILLER_26_529 ();
 sg13g2_decap_8 FILLER_26_536 ();
 sg13g2_decap_8 FILLER_26_543 ();
 sg13g2_decap_8 FILLER_26_550 ();
 sg13g2_decap_8 FILLER_26_557 ();
 sg13g2_decap_8 FILLER_26_564 ();
 sg13g2_decap_8 FILLER_26_571 ();
 sg13g2_decap_8 FILLER_26_578 ();
 sg13g2_decap_8 FILLER_26_585 ();
 sg13g2_decap_8 FILLER_26_592 ();
 sg13g2_decap_8 FILLER_26_599 ();
 sg13g2_decap_8 FILLER_26_606 ();
 sg13g2_decap_8 FILLER_26_613 ();
 sg13g2_decap_8 FILLER_26_620 ();
 sg13g2_decap_8 FILLER_26_627 ();
 sg13g2_decap_8 FILLER_26_634 ();
 sg13g2_decap_8 FILLER_26_641 ();
 sg13g2_decap_8 FILLER_26_648 ();
 sg13g2_decap_8 FILLER_26_655 ();
 sg13g2_decap_8 FILLER_26_662 ();
 sg13g2_decap_8 FILLER_26_669 ();
 sg13g2_decap_8 FILLER_26_676 ();
 sg13g2_decap_8 FILLER_26_683 ();
 sg13g2_decap_8 FILLER_26_690 ();
 sg13g2_decap_8 FILLER_26_697 ();
 sg13g2_decap_8 FILLER_26_704 ();
 sg13g2_decap_8 FILLER_26_711 ();
 sg13g2_decap_8 FILLER_26_718 ();
 sg13g2_decap_8 FILLER_26_725 ();
 sg13g2_decap_8 FILLER_26_732 ();
 sg13g2_decap_8 FILLER_26_739 ();
 sg13g2_decap_8 FILLER_26_746 ();
 sg13g2_decap_8 FILLER_26_753 ();
 sg13g2_decap_8 FILLER_26_760 ();
 sg13g2_decap_8 FILLER_26_767 ();
 sg13g2_decap_8 FILLER_26_774 ();
 sg13g2_decap_8 FILLER_26_781 ();
 sg13g2_decap_8 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_795 ();
 sg13g2_decap_8 FILLER_26_802 ();
 sg13g2_decap_8 FILLER_26_809 ();
 sg13g2_decap_8 FILLER_26_816 ();
 sg13g2_decap_8 FILLER_26_823 ();
 sg13g2_decap_8 FILLER_26_830 ();
 sg13g2_decap_8 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_844 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_decap_8 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_26_865 ();
 sg13g2_decap_8 FILLER_26_872 ();
 sg13g2_decap_8 FILLER_26_879 ();
 sg13g2_decap_8 FILLER_26_886 ();
 sg13g2_decap_8 FILLER_26_893 ();
 sg13g2_decap_8 FILLER_26_900 ();
 sg13g2_decap_8 FILLER_26_907 ();
 sg13g2_decap_8 FILLER_26_914 ();
 sg13g2_decap_8 FILLER_26_921 ();
 sg13g2_decap_8 FILLER_26_928 ();
 sg13g2_decap_8 FILLER_26_935 ();
 sg13g2_decap_8 FILLER_26_942 ();
 sg13g2_decap_8 FILLER_26_949 ();
 sg13g2_decap_8 FILLER_26_956 ();
 sg13g2_decap_8 FILLER_26_963 ();
 sg13g2_decap_8 FILLER_26_970 ();
 sg13g2_decap_8 FILLER_26_977 ();
 sg13g2_decap_8 FILLER_26_984 ();
 sg13g2_decap_8 FILLER_26_991 ();
 sg13g2_decap_8 FILLER_26_998 ();
 sg13g2_decap_8 FILLER_26_1005 ();
 sg13g2_decap_8 FILLER_26_1012 ();
 sg13g2_decap_8 FILLER_26_1019 ();
 sg13g2_fill_2 FILLER_26_1026 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_44 ();
 sg13g2_decap_8 FILLER_27_72 ();
 sg13g2_decap_8 FILLER_27_79 ();
 sg13g2_decap_8 FILLER_27_86 ();
 sg13g2_decap_8 FILLER_27_93 ();
 sg13g2_decap_8 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_107 ();
 sg13g2_decap_8 FILLER_27_114 ();
 sg13g2_decap_8 FILLER_27_121 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_156 ();
 sg13g2_decap_8 FILLER_27_163 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_177 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_decap_8 FILLER_27_226 ();
 sg13g2_decap_8 FILLER_27_233 ();
 sg13g2_decap_8 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_247 ();
 sg13g2_decap_8 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_261 ();
 sg13g2_decap_8 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_275 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_decap_8 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_27_436 ();
 sg13g2_decap_8 FILLER_27_443 ();
 sg13g2_decap_8 FILLER_27_450 ();
 sg13g2_decap_8 FILLER_27_457 ();
 sg13g2_decap_8 FILLER_27_464 ();
 sg13g2_decap_8 FILLER_27_471 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_8 FILLER_27_485 ();
 sg13g2_decap_8 FILLER_27_492 ();
 sg13g2_decap_8 FILLER_27_499 ();
 sg13g2_decap_8 FILLER_27_506 ();
 sg13g2_decap_8 FILLER_27_513 ();
 sg13g2_decap_8 FILLER_27_520 ();
 sg13g2_decap_8 FILLER_27_527 ();
 sg13g2_decap_8 FILLER_27_534 ();
 sg13g2_decap_8 FILLER_27_541 ();
 sg13g2_decap_8 FILLER_27_548 ();
 sg13g2_decap_8 FILLER_27_555 ();
 sg13g2_decap_8 FILLER_27_562 ();
 sg13g2_decap_8 FILLER_27_569 ();
 sg13g2_decap_8 FILLER_27_576 ();
 sg13g2_decap_8 FILLER_27_583 ();
 sg13g2_decap_8 FILLER_27_590 ();
 sg13g2_decap_8 FILLER_27_597 ();
 sg13g2_decap_8 FILLER_27_604 ();
 sg13g2_decap_8 FILLER_27_611 ();
 sg13g2_decap_8 FILLER_27_618 ();
 sg13g2_decap_8 FILLER_27_625 ();
 sg13g2_decap_8 FILLER_27_632 ();
 sg13g2_decap_8 FILLER_27_639 ();
 sg13g2_decap_8 FILLER_27_646 ();
 sg13g2_decap_8 FILLER_27_653 ();
 sg13g2_decap_8 FILLER_27_660 ();
 sg13g2_decap_8 FILLER_27_667 ();
 sg13g2_decap_8 FILLER_27_674 ();
 sg13g2_decap_8 FILLER_27_681 ();
 sg13g2_decap_8 FILLER_27_688 ();
 sg13g2_decap_8 FILLER_27_695 ();
 sg13g2_decap_8 FILLER_27_702 ();
 sg13g2_decap_8 FILLER_27_709 ();
 sg13g2_decap_8 FILLER_27_716 ();
 sg13g2_decap_8 FILLER_27_723 ();
 sg13g2_decap_8 FILLER_27_730 ();
 sg13g2_decap_8 FILLER_27_737 ();
 sg13g2_decap_8 FILLER_27_744 ();
 sg13g2_decap_8 FILLER_27_751 ();
 sg13g2_decap_8 FILLER_27_758 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_decap_8 FILLER_27_772 ();
 sg13g2_decap_8 FILLER_27_779 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_decap_8 FILLER_27_954 ();
 sg13g2_decap_8 FILLER_27_961 ();
 sg13g2_decap_8 FILLER_27_968 ();
 sg13g2_decap_8 FILLER_27_975 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_4 FILLER_27_1024 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_277 ();
 sg13g2_decap_8 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_8 FILLER_28_424 ();
 sg13g2_decap_8 FILLER_28_431 ();
 sg13g2_decap_8 FILLER_28_438 ();
 sg13g2_decap_8 FILLER_28_445 ();
 sg13g2_decap_8 FILLER_28_452 ();
 sg13g2_decap_8 FILLER_28_459 ();
 sg13g2_decap_8 FILLER_28_466 ();
 sg13g2_decap_8 FILLER_28_473 ();
 sg13g2_decap_8 FILLER_28_480 ();
 sg13g2_decap_8 FILLER_28_487 ();
 sg13g2_decap_8 FILLER_28_494 ();
 sg13g2_decap_8 FILLER_28_501 ();
 sg13g2_decap_8 FILLER_28_508 ();
 sg13g2_decap_8 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_522 ();
 sg13g2_decap_8 FILLER_28_529 ();
 sg13g2_decap_8 FILLER_28_536 ();
 sg13g2_decap_8 FILLER_28_543 ();
 sg13g2_decap_8 FILLER_28_550 ();
 sg13g2_decap_8 FILLER_28_557 ();
 sg13g2_decap_8 FILLER_28_564 ();
 sg13g2_decap_8 FILLER_28_571 ();
 sg13g2_decap_8 FILLER_28_578 ();
 sg13g2_decap_8 FILLER_28_585 ();
 sg13g2_decap_8 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_599 ();
 sg13g2_decap_8 FILLER_28_606 ();
 sg13g2_decap_8 FILLER_28_613 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_decap_8 FILLER_28_634 ();
 sg13g2_decap_8 FILLER_28_641 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_655 ();
 sg13g2_decap_8 FILLER_28_662 ();
 sg13g2_decap_8 FILLER_28_669 ();
 sg13g2_decap_8 FILLER_28_676 ();
 sg13g2_decap_8 FILLER_28_683 ();
 sg13g2_decap_8 FILLER_28_690 ();
 sg13g2_decap_8 FILLER_28_697 ();
 sg13g2_decap_8 FILLER_28_704 ();
 sg13g2_decap_8 FILLER_28_711 ();
 sg13g2_decap_8 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_725 ();
 sg13g2_decap_8 FILLER_28_732 ();
 sg13g2_decap_8 FILLER_28_739 ();
 sg13g2_decap_8 FILLER_28_746 ();
 sg13g2_decap_8 FILLER_28_753 ();
 sg13g2_decap_8 FILLER_28_760 ();
 sg13g2_decap_8 FILLER_28_767 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_decap_8 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_788 ();
 sg13g2_decap_8 FILLER_28_795 ();
 sg13g2_decap_8 FILLER_28_802 ();
 sg13g2_decap_8 FILLER_28_809 ();
 sg13g2_decap_8 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_8 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_28_865 ();
 sg13g2_decap_8 FILLER_28_872 ();
 sg13g2_decap_8 FILLER_28_879 ();
 sg13g2_decap_8 FILLER_28_886 ();
 sg13g2_decap_8 FILLER_28_893 ();
 sg13g2_decap_8 FILLER_28_900 ();
 sg13g2_decap_8 FILLER_28_907 ();
 sg13g2_decap_8 FILLER_28_914 ();
 sg13g2_decap_8 FILLER_28_921 ();
 sg13g2_decap_8 FILLER_28_928 ();
 sg13g2_decap_8 FILLER_28_935 ();
 sg13g2_decap_8 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_949 ();
 sg13g2_decap_8 FILLER_28_956 ();
 sg13g2_decap_8 FILLER_28_963 ();
 sg13g2_decap_8 FILLER_28_970 ();
 sg13g2_decap_8 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_984 ();
 sg13g2_decap_8 FILLER_28_991 ();
 sg13g2_decap_8 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1005 ();
 sg13g2_decap_8 FILLER_28_1012 ();
 sg13g2_decap_8 FILLER_28_1019 ();
 sg13g2_fill_2 FILLER_28_1026 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_decap_8 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_18 ();
 sg13g2_decap_8 FILLER_29_25 ();
 sg13g2_decap_8 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_95 ();
 sg13g2_decap_8 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_109 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_137 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_200 ();
 sg13g2_decap_8 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_417 ();
 sg13g2_decap_8 FILLER_29_424 ();
 sg13g2_decap_8 FILLER_29_431 ();
 sg13g2_decap_8 FILLER_29_438 ();
 sg13g2_decap_8 FILLER_29_445 ();
 sg13g2_decap_8 FILLER_29_452 ();
 sg13g2_decap_8 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_466 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_decap_8 FILLER_29_480 ();
 sg13g2_decap_8 FILLER_29_487 ();
 sg13g2_decap_8 FILLER_29_494 ();
 sg13g2_decap_8 FILLER_29_501 ();
 sg13g2_decap_8 FILLER_29_508 ();
 sg13g2_decap_8 FILLER_29_515 ();
 sg13g2_decap_8 FILLER_29_522 ();
 sg13g2_decap_8 FILLER_29_529 ();
 sg13g2_decap_8 FILLER_29_536 ();
 sg13g2_decap_8 FILLER_29_543 ();
 sg13g2_decap_8 FILLER_29_550 ();
 sg13g2_decap_8 FILLER_29_557 ();
 sg13g2_decap_8 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_571 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_decap_8 FILLER_29_599 ();
 sg13g2_decap_8 FILLER_29_606 ();
 sg13g2_decap_8 FILLER_29_613 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_decap_8 FILLER_29_627 ();
 sg13g2_decap_8 FILLER_29_634 ();
 sg13g2_decap_8 FILLER_29_641 ();
 sg13g2_decap_8 FILLER_29_648 ();
 sg13g2_decap_8 FILLER_29_655 ();
 sg13g2_decap_8 FILLER_29_662 ();
 sg13g2_decap_8 FILLER_29_669 ();
 sg13g2_decap_8 FILLER_29_676 ();
 sg13g2_decap_8 FILLER_29_683 ();
 sg13g2_decap_8 FILLER_29_690 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_decap_8 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_711 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_decap_8 FILLER_29_746 ();
 sg13g2_decap_8 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_decap_8 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_8 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_29_865 ();
 sg13g2_decap_8 FILLER_29_872 ();
 sg13g2_decap_8 FILLER_29_879 ();
 sg13g2_decap_8 FILLER_29_886 ();
 sg13g2_decap_8 FILLER_29_893 ();
 sg13g2_decap_8 FILLER_29_900 ();
 sg13g2_decap_8 FILLER_29_907 ();
 sg13g2_decap_8 FILLER_29_914 ();
 sg13g2_decap_8 FILLER_29_921 ();
 sg13g2_decap_8 FILLER_29_928 ();
 sg13g2_decap_8 FILLER_29_935 ();
 sg13g2_decap_8 FILLER_29_942 ();
 sg13g2_decap_8 FILLER_29_949 ();
 sg13g2_decap_8 FILLER_29_956 ();
 sg13g2_decap_8 FILLER_29_963 ();
 sg13g2_decap_8 FILLER_29_970 ();
 sg13g2_decap_8 FILLER_29_977 ();
 sg13g2_decap_8 FILLER_29_984 ();
 sg13g2_decap_8 FILLER_29_991 ();
 sg13g2_decap_8 FILLER_29_998 ();
 sg13g2_decap_8 FILLER_29_1005 ();
 sg13g2_decap_8 FILLER_29_1012 ();
 sg13g2_decap_8 FILLER_29_1019 ();
 sg13g2_fill_2 FILLER_29_1026 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_decap_8 FILLER_30_875 ();
 sg13g2_decap_8 FILLER_30_882 ();
 sg13g2_decap_8 FILLER_30_889 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_decap_8 FILLER_30_903 ();
 sg13g2_decap_8 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_917 ();
 sg13g2_decap_8 FILLER_30_924 ();
 sg13g2_decap_8 FILLER_30_931 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_8 FILLER_30_945 ();
 sg13g2_decap_8 FILLER_30_952 ();
 sg13g2_decap_8 FILLER_30_959 ();
 sg13g2_decap_8 FILLER_30_966 ();
 sg13g2_decap_8 FILLER_30_973 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_987 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1001 ();
 sg13g2_decap_8 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1015 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_decap_8 FILLER_31_882 ();
 sg13g2_decap_8 FILLER_31_889 ();
 sg13g2_decap_8 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_903 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_966 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_decap_8 FILLER_31_980 ();
 sg13g2_decap_8 FILLER_31_987 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_546 ();
 sg13g2_decap_8 FILLER_32_553 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_decap_8 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_32_868 ();
 sg13g2_decap_8 FILLER_32_875 ();
 sg13g2_decap_8 FILLER_32_882 ();
 sg13g2_decap_8 FILLER_32_889 ();
 sg13g2_decap_8 FILLER_32_896 ();
 sg13g2_decap_8 FILLER_32_903 ();
 sg13g2_decap_8 FILLER_32_910 ();
 sg13g2_decap_8 FILLER_32_917 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_decap_8 FILLER_32_931 ();
 sg13g2_decap_8 FILLER_32_938 ();
 sg13g2_decap_8 FILLER_32_945 ();
 sg13g2_decap_8 FILLER_32_952 ();
 sg13g2_decap_8 FILLER_32_959 ();
 sg13g2_decap_8 FILLER_32_966 ();
 sg13g2_decap_8 FILLER_32_973 ();
 sg13g2_decap_8 FILLER_32_980 ();
 sg13g2_decap_8 FILLER_32_987 ();
 sg13g2_decap_8 FILLER_32_994 ();
 sg13g2_decap_8 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1008 ();
 sg13g2_decap_8 FILLER_32_1015 ();
 sg13g2_decap_8 FILLER_32_1022 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_decap_8 FILLER_33_875 ();
 sg13g2_decap_8 FILLER_33_882 ();
 sg13g2_decap_8 FILLER_33_889 ();
 sg13g2_decap_8 FILLER_33_896 ();
 sg13g2_decap_8 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_decap_8 FILLER_33_938 ();
 sg13g2_decap_8 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_959 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_973 ();
 sg13g2_decap_8 FILLER_33_980 ();
 sg13g2_decap_8 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_511 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_560 ();
 sg13g2_decap_8 FILLER_34_567 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_700 ();
 sg13g2_decap_8 FILLER_34_707 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_decap_8 FILLER_34_721 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_34_868 ();
 sg13g2_decap_8 FILLER_34_875 ();
 sg13g2_decap_8 FILLER_34_882 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_decap_8 FILLER_34_896 ();
 sg13g2_decap_8 FILLER_34_903 ();
 sg13g2_decap_8 FILLER_34_910 ();
 sg13g2_decap_8 FILLER_34_917 ();
 sg13g2_decap_8 FILLER_34_924 ();
 sg13g2_decap_8 FILLER_34_931 ();
 sg13g2_decap_8 FILLER_34_938 ();
 sg13g2_decap_8 FILLER_34_945 ();
 sg13g2_decap_8 FILLER_34_952 ();
 sg13g2_decap_8 FILLER_34_959 ();
 sg13g2_decap_8 FILLER_34_966 ();
 sg13g2_decap_8 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_980 ();
 sg13g2_decap_8 FILLER_34_987 ();
 sg13g2_decap_8 FILLER_34_994 ();
 sg13g2_decap_8 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1008 ();
 sg13g2_decap_8 FILLER_34_1015 ();
 sg13g2_decap_8 FILLER_34_1022 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_567 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_616 ();
 sg13g2_decap_8 FILLER_35_623 ();
 sg13g2_decap_8 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_decap_8 FILLER_35_651 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_decap_8 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_35_868 ();
 sg13g2_decap_8 FILLER_35_875 ();
 sg13g2_decap_8 FILLER_35_882 ();
 sg13g2_decap_8 FILLER_35_889 ();
 sg13g2_decap_8 FILLER_35_896 ();
 sg13g2_decap_8 FILLER_35_903 ();
 sg13g2_decap_8 FILLER_35_910 ();
 sg13g2_decap_8 FILLER_35_917 ();
 sg13g2_decap_8 FILLER_35_924 ();
 sg13g2_decap_8 FILLER_35_931 ();
 sg13g2_decap_8 FILLER_35_938 ();
 sg13g2_decap_8 FILLER_35_945 ();
 sg13g2_decap_8 FILLER_35_952 ();
 sg13g2_decap_8 FILLER_35_959 ();
 sg13g2_decap_8 FILLER_35_966 ();
 sg13g2_decap_8 FILLER_35_973 ();
 sg13g2_decap_8 FILLER_35_980 ();
 sg13g2_decap_8 FILLER_35_987 ();
 sg13g2_decap_8 FILLER_35_994 ();
 sg13g2_decap_8 FILLER_35_1001 ();
 sg13g2_decap_8 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1015 ();
 sg13g2_decap_8 FILLER_35_1022 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_462 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_483 ();
 sg13g2_decap_8 FILLER_36_490 ();
 sg13g2_decap_8 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_511 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_567 ();
 sg13g2_decap_8 FILLER_36_574 ();
 sg13g2_decap_8 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_595 ();
 sg13g2_decap_8 FILLER_36_602 ();
 sg13g2_decap_8 FILLER_36_609 ();
 sg13g2_decap_8 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_630 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_672 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_decap_8 FILLER_36_686 ();
 sg13g2_decap_8 FILLER_36_693 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_decap_8 FILLER_36_707 ();
 sg13g2_decap_8 FILLER_36_714 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_decap_8 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_8 FILLER_36_854 ();
 sg13g2_decap_8 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_36_868 ();
 sg13g2_decap_8 FILLER_36_875 ();
 sg13g2_decap_8 FILLER_36_882 ();
 sg13g2_decap_8 FILLER_36_889 ();
 sg13g2_decap_8 FILLER_36_896 ();
 sg13g2_decap_8 FILLER_36_903 ();
 sg13g2_decap_8 FILLER_36_910 ();
 sg13g2_decap_8 FILLER_36_917 ();
 sg13g2_decap_8 FILLER_36_924 ();
 sg13g2_decap_8 FILLER_36_931 ();
 sg13g2_decap_8 FILLER_36_938 ();
 sg13g2_decap_8 FILLER_36_945 ();
 sg13g2_decap_8 FILLER_36_952 ();
 sg13g2_decap_8 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_966 ();
 sg13g2_decap_8 FILLER_36_973 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_896 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_37_931 ();
 sg13g2_decap_8 FILLER_37_938 ();
 sg13g2_decap_8 FILLER_37_945 ();
 sg13g2_decap_8 FILLER_37_952 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_decap_8 FILLER_37_973 ();
 sg13g2_decap_8 FILLER_37_980 ();
 sg13g2_decap_8 FILLER_37_987 ();
 sg13g2_decap_8 FILLER_37_994 ();
 sg13g2_decap_8 FILLER_37_1001 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_decap_8 FILLER_37_1022 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_448 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_462 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_8 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_decap_8 FILLER_38_497 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_decap_8 FILLER_38_511 ();
 sg13g2_decap_8 FILLER_38_518 ();
 sg13g2_decap_8 FILLER_38_525 ();
 sg13g2_decap_8 FILLER_38_532 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_553 ();
 sg13g2_decap_8 FILLER_38_560 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_decap_8 FILLER_38_602 ();
 sg13g2_decap_8 FILLER_38_609 ();
 sg13g2_decap_8 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_decap_8 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_644 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_8 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_679 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_38_868 ();
 sg13g2_decap_8 FILLER_38_875 ();
 sg13g2_decap_8 FILLER_38_882 ();
 sg13g2_decap_8 FILLER_38_889 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_decap_8 FILLER_38_903 ();
 sg13g2_decap_8 FILLER_38_910 ();
 sg13g2_decap_8 FILLER_38_917 ();
 sg13g2_decap_8 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_38_931 ();
 sg13g2_decap_8 FILLER_38_938 ();
 sg13g2_decap_8 FILLER_38_945 ();
 sg13g2_decap_8 FILLER_38_952 ();
 sg13g2_decap_8 FILLER_38_959 ();
 sg13g2_decap_8 FILLER_38_966 ();
 sg13g2_decap_8 FILLER_38_973 ();
 sg13g2_decap_8 FILLER_38_980 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_decap_8 FILLER_38_1001 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_decap_8 FILLER_38_1015 ();
 sg13g2_decap_8 FILLER_38_1022 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_511 ();
 sg13g2_decap_8 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_525 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_8 FILLER_39_546 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_decap_8 FILLER_39_560 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_8 FILLER_39_581 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_decap_8 FILLER_39_644 ();
 sg13g2_decap_8 FILLER_39_651 ();
 sg13g2_decap_8 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_693 ();
 sg13g2_decap_8 FILLER_39_700 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_756 ();
 sg13g2_decap_8 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_791 ();
 sg13g2_decap_8 FILLER_39_798 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_decap_8 FILLER_39_875 ();
 sg13g2_decap_8 FILLER_39_882 ();
 sg13g2_decap_8 FILLER_39_889 ();
 sg13g2_decap_8 FILLER_39_896 ();
 sg13g2_decap_8 FILLER_39_903 ();
 sg13g2_decap_8 FILLER_39_910 ();
 sg13g2_decap_8 FILLER_39_917 ();
 sg13g2_decap_8 FILLER_39_924 ();
 sg13g2_decap_8 FILLER_39_931 ();
 sg13g2_decap_8 FILLER_39_938 ();
 sg13g2_decap_8 FILLER_39_945 ();
 sg13g2_decap_8 FILLER_39_952 ();
 sg13g2_decap_8 FILLER_39_959 ();
 sg13g2_decap_8 FILLER_39_966 ();
 sg13g2_decap_8 FILLER_39_973 ();
 sg13g2_decap_8 FILLER_39_980 ();
 sg13g2_decap_8 FILLER_39_987 ();
 sg13g2_decap_8 FILLER_39_994 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_8 FILLER_39_1008 ();
 sg13g2_decap_8 FILLER_39_1015 ();
 sg13g2_decap_8 FILLER_39_1022 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_decap_8 FILLER_40_567 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_658 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_decap_8 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_40_868 ();
 sg13g2_decap_8 FILLER_40_875 ();
 sg13g2_decap_8 FILLER_40_882 ();
 sg13g2_decap_8 FILLER_40_889 ();
 sg13g2_decap_8 FILLER_40_896 ();
 sg13g2_decap_8 FILLER_40_903 ();
 sg13g2_decap_8 FILLER_40_910 ();
 sg13g2_decap_8 FILLER_40_917 ();
 sg13g2_decap_8 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_938 ();
 sg13g2_decap_8 FILLER_40_945 ();
 sg13g2_decap_8 FILLER_40_952 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_decap_8 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_987 ();
 sg13g2_decap_8 FILLER_40_994 ();
 sg13g2_decap_8 FILLER_40_1001 ();
 sg13g2_decap_8 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_518 ();
 sg13g2_decap_8 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_8 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_8 FILLER_41_602 ();
 sg13g2_decap_8 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_decap_8 FILLER_41_875 ();
 sg13g2_decap_8 FILLER_41_882 ();
 sg13g2_decap_8 FILLER_41_889 ();
 sg13g2_decap_8 FILLER_41_896 ();
 sg13g2_decap_8 FILLER_41_903 ();
 sg13g2_decap_8 FILLER_41_910 ();
 sg13g2_decap_8 FILLER_41_917 ();
 sg13g2_decap_8 FILLER_41_924 ();
 sg13g2_decap_8 FILLER_41_931 ();
 sg13g2_decap_8 FILLER_41_938 ();
 sg13g2_decap_8 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_952 ();
 sg13g2_decap_8 FILLER_41_959 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_980 ();
 sg13g2_decap_8 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_994 ();
 sg13g2_decap_8 FILLER_41_1001 ();
 sg13g2_decap_8 FILLER_41_1008 ();
 sg13g2_decap_8 FILLER_41_1015 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_8 FILLER_42_511 ();
 sg13g2_decap_8 FILLER_42_518 ();
 sg13g2_decap_8 FILLER_42_525 ();
 sg13g2_decap_8 FILLER_42_532 ();
 sg13g2_decap_8 FILLER_42_539 ();
 sg13g2_decap_8 FILLER_42_546 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_560 ();
 sg13g2_decap_8 FILLER_42_567 ();
 sg13g2_decap_8 FILLER_42_574 ();
 sg13g2_decap_8 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_588 ();
 sg13g2_decap_8 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_602 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_decap_8 FILLER_42_616 ();
 sg13g2_decap_8 FILLER_42_623 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_651 ();
 sg13g2_decap_8 FILLER_42_658 ();
 sg13g2_decap_8 FILLER_42_665 ();
 sg13g2_decap_8 FILLER_42_672 ();
 sg13g2_decap_8 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_8 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_decap_8 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_42_868 ();
 sg13g2_decap_8 FILLER_42_875 ();
 sg13g2_decap_8 FILLER_42_882 ();
 sg13g2_decap_8 FILLER_42_889 ();
 sg13g2_decap_8 FILLER_42_896 ();
 sg13g2_decap_8 FILLER_42_903 ();
 sg13g2_decap_8 FILLER_42_910 ();
 sg13g2_decap_8 FILLER_42_917 ();
 sg13g2_decap_8 FILLER_42_924 ();
 sg13g2_decap_8 FILLER_42_931 ();
 sg13g2_decap_8 FILLER_42_938 ();
 sg13g2_decap_8 FILLER_42_945 ();
 sg13g2_decap_8 FILLER_42_952 ();
 sg13g2_decap_8 FILLER_42_959 ();
 sg13g2_decap_8 FILLER_42_966 ();
 sg13g2_decap_8 FILLER_42_973 ();
 sg13g2_decap_8 FILLER_42_980 ();
 sg13g2_decap_8 FILLER_42_987 ();
 sg13g2_decap_8 FILLER_42_994 ();
 sg13g2_decap_8 FILLER_42_1001 ();
 sg13g2_decap_8 FILLER_42_1008 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_decap_8 FILLER_42_1022 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_decap_8 FILLER_43_504 ();
 sg13g2_decap_8 FILLER_43_511 ();
 sg13g2_decap_8 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_8 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_decap_8 FILLER_43_567 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_8 FILLER_43_581 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_882 ();
 sg13g2_decap_8 FILLER_43_889 ();
 sg13g2_decap_8 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_903 ();
 sg13g2_decap_8 FILLER_43_910 ();
 sg13g2_decap_8 FILLER_43_917 ();
 sg13g2_decap_8 FILLER_43_924 ();
 sg13g2_decap_8 FILLER_43_931 ();
 sg13g2_decap_8 FILLER_43_938 ();
 sg13g2_decap_8 FILLER_43_945 ();
 sg13g2_decap_8 FILLER_43_952 ();
 sg13g2_decap_8 FILLER_43_959 ();
 sg13g2_decap_8 FILLER_43_966 ();
 sg13g2_decap_8 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_980 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_994 ();
 sg13g2_decap_8 FILLER_43_1001 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_decap_8 FILLER_44_483 ();
 sg13g2_decap_8 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_decap_8 FILLER_44_504 ();
 sg13g2_decap_8 FILLER_44_511 ();
 sg13g2_decap_8 FILLER_44_518 ();
 sg13g2_decap_8 FILLER_44_525 ();
 sg13g2_decap_8 FILLER_44_532 ();
 sg13g2_decap_8 FILLER_44_539 ();
 sg13g2_decap_8 FILLER_44_546 ();
 sg13g2_decap_8 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_8 FILLER_44_567 ();
 sg13g2_decap_8 FILLER_44_574 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_decap_8 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_609 ();
 sg13g2_decap_8 FILLER_44_616 ();
 sg13g2_decap_8 FILLER_44_623 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_decap_8 FILLER_44_637 ();
 sg13g2_decap_8 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_651 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_693 ();
 sg13g2_decap_8 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_714 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_decap_8 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_44_868 ();
 sg13g2_decap_8 FILLER_44_875 ();
 sg13g2_decap_8 FILLER_44_882 ();
 sg13g2_decap_8 FILLER_44_889 ();
 sg13g2_decap_8 FILLER_44_896 ();
 sg13g2_decap_8 FILLER_44_903 ();
 sg13g2_decap_8 FILLER_44_910 ();
 sg13g2_decap_8 FILLER_44_917 ();
 sg13g2_decap_8 FILLER_44_924 ();
 sg13g2_decap_8 FILLER_44_931 ();
 sg13g2_decap_8 FILLER_44_938 ();
 sg13g2_decap_8 FILLER_44_945 ();
 sg13g2_decap_8 FILLER_44_952 ();
 sg13g2_decap_8 FILLER_44_959 ();
 sg13g2_decap_8 FILLER_44_966 ();
 sg13g2_decap_8 FILLER_44_973 ();
 sg13g2_decap_8 FILLER_44_980 ();
 sg13g2_decap_8 FILLER_44_987 ();
 sg13g2_decap_8 FILLER_44_994 ();
 sg13g2_decap_8 FILLER_44_1001 ();
 sg13g2_decap_8 FILLER_44_1008 ();
 sg13g2_decap_8 FILLER_44_1015 ();
 sg13g2_decap_8 FILLER_44_1022 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_525 ();
 sg13g2_decap_8 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_decap_8 FILLER_45_553 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_567 ();
 sg13g2_decap_8 FILLER_45_574 ();
 sg13g2_decap_8 FILLER_45_581 ();
 sg13g2_decap_8 FILLER_45_588 ();
 sg13g2_decap_8 FILLER_45_595 ();
 sg13g2_decap_8 FILLER_45_602 ();
 sg13g2_decap_8 FILLER_45_609 ();
 sg13g2_decap_8 FILLER_45_616 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_decap_8 FILLER_45_630 ();
 sg13g2_decap_8 FILLER_45_637 ();
 sg13g2_decap_8 FILLER_45_644 ();
 sg13g2_decap_8 FILLER_45_651 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_672 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_707 ();
 sg13g2_decap_8 FILLER_45_714 ();
 sg13g2_decap_8 FILLER_45_721 ();
 sg13g2_decap_8 FILLER_45_728 ();
 sg13g2_decap_8 FILLER_45_735 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_decap_8 FILLER_45_749 ();
 sg13g2_decap_8 FILLER_45_756 ();
 sg13g2_decap_8 FILLER_45_763 ();
 sg13g2_decap_8 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_777 ();
 sg13g2_decap_8 FILLER_45_784 ();
 sg13g2_decap_8 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_812 ();
 sg13g2_decap_8 FILLER_45_819 ();
 sg13g2_decap_8 FILLER_45_826 ();
 sg13g2_decap_8 FILLER_45_833 ();
 sg13g2_decap_8 FILLER_45_840 ();
 sg13g2_decap_8 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_decap_8 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_45_868 ();
 sg13g2_decap_8 FILLER_45_875 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_8 FILLER_45_889 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_decap_8 FILLER_45_903 ();
 sg13g2_decap_8 FILLER_45_910 ();
 sg13g2_decap_8 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_924 ();
 sg13g2_decap_8 FILLER_45_931 ();
 sg13g2_decap_8 FILLER_45_938 ();
 sg13g2_decap_8 FILLER_45_945 ();
 sg13g2_decap_8 FILLER_45_952 ();
 sg13g2_decap_8 FILLER_45_959 ();
 sg13g2_decap_8 FILLER_45_966 ();
 sg13g2_decap_8 FILLER_45_973 ();
 sg13g2_decap_8 FILLER_45_980 ();
 sg13g2_decap_8 FILLER_45_987 ();
 sg13g2_decap_8 FILLER_45_994 ();
 sg13g2_decap_8 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_8 FILLER_46_889 ();
 sg13g2_decap_8 FILLER_46_896 ();
 sg13g2_decap_8 FILLER_46_903 ();
 sg13g2_decap_8 FILLER_46_910 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_decap_8 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_931 ();
 sg13g2_decap_8 FILLER_46_938 ();
 sg13g2_decap_8 FILLER_46_945 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_994 ();
 sg13g2_decap_8 FILLER_46_1001 ();
 sg13g2_decap_8 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1022 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_48_931 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_945 ();
 sg13g2_decap_8 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_959 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_298 ();
 sg13g2_decap_8 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_312 ();
 sg13g2_decap_8 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_decap_8 FILLER_49_340 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_8 FILLER_49_424 ();
 sg13g2_decap_8 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_494 ();
 sg13g2_decap_8 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_508 ();
 sg13g2_decap_8 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_522 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_550 ();
 sg13g2_decap_8 FILLER_49_557 ();
 sg13g2_decap_8 FILLER_49_564 ();
 sg13g2_decap_8 FILLER_49_571 ();
 sg13g2_decap_8 FILLER_49_578 ();
 sg13g2_decap_8 FILLER_49_585 ();
 sg13g2_decap_8 FILLER_49_592 ();
 sg13g2_decap_8 FILLER_49_599 ();
 sg13g2_decap_8 FILLER_49_606 ();
 sg13g2_decap_8 FILLER_49_613 ();
 sg13g2_decap_8 FILLER_49_620 ();
 sg13g2_decap_8 FILLER_49_627 ();
 sg13g2_decap_8 FILLER_49_634 ();
 sg13g2_decap_8 FILLER_49_641 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_decap_8 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_662 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_decap_8 FILLER_49_683 ();
 sg13g2_decap_8 FILLER_49_690 ();
 sg13g2_decap_8 FILLER_49_697 ();
 sg13g2_decap_8 FILLER_49_704 ();
 sg13g2_decap_8 FILLER_49_711 ();
 sg13g2_decap_8 FILLER_49_718 ();
 sg13g2_decap_8 FILLER_49_725 ();
 sg13g2_decap_8 FILLER_49_732 ();
 sg13g2_decap_8 FILLER_49_739 ();
 sg13g2_decap_8 FILLER_49_746 ();
 sg13g2_decap_8 FILLER_49_753 ();
 sg13g2_decap_8 FILLER_49_760 ();
 sg13g2_decap_8 FILLER_49_767 ();
 sg13g2_decap_8 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_781 ();
 sg13g2_decap_8 FILLER_49_788 ();
 sg13g2_decap_8 FILLER_49_795 ();
 sg13g2_decap_8 FILLER_49_802 ();
 sg13g2_decap_8 FILLER_49_809 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_decap_8 FILLER_49_823 ();
 sg13g2_decap_8 FILLER_49_830 ();
 sg13g2_decap_8 FILLER_49_837 ();
 sg13g2_decap_8 FILLER_49_844 ();
 sg13g2_decap_8 FILLER_49_851 ();
 sg13g2_decap_8 FILLER_49_858 ();
 sg13g2_decap_8 FILLER_49_865 ();
 sg13g2_decap_8 FILLER_49_872 ();
 sg13g2_decap_8 FILLER_49_879 ();
 sg13g2_decap_8 FILLER_49_886 ();
 sg13g2_decap_8 FILLER_49_893 ();
 sg13g2_decap_8 FILLER_49_900 ();
 sg13g2_decap_8 FILLER_49_907 ();
 sg13g2_decap_8 FILLER_49_914 ();
 sg13g2_decap_8 FILLER_49_921 ();
 sg13g2_decap_8 FILLER_49_928 ();
 sg13g2_decap_8 FILLER_49_935 ();
 sg13g2_decap_8 FILLER_49_942 ();
 sg13g2_decap_8 FILLER_49_949 ();
 sg13g2_decap_8 FILLER_49_956 ();
 sg13g2_decap_8 FILLER_49_963 ();
 sg13g2_decap_8 FILLER_49_970 ();
 sg13g2_decap_8 FILLER_49_977 ();
 sg13g2_decap_8 FILLER_49_984 ();
 sg13g2_decap_8 FILLER_49_991 ();
 sg13g2_decap_8 FILLER_49_998 ();
 sg13g2_decap_8 FILLER_49_1005 ();
 sg13g2_decap_8 FILLER_49_1012 ();
 sg13g2_decap_8 FILLER_49_1019 ();
 sg13g2_fill_2 FILLER_49_1026 ();
 sg13g2_fill_1 FILLER_49_1028 ();
 assign uio_oe[0] = net26;
 assign uio_oe[1] = net27;
 assign uio_oe[2] = net28;
 assign uio_oe[3] = net29;
 assign uio_oe[4] = net30;
 assign uio_oe[5] = net31;
 assign uio_oe[6] = net32;
 assign uio_oe[7] = net33;
endmodule
