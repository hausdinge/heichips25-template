VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO heichips25_internal
  CLASS BLOCK ;
  FOREIGN heichips25_internal ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 21.580 3.150 23.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 97.180 3.150 99.380 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 172.780 3.150 174.980 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 248.380 3.150 250.580 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 323.980 3.150 326.180 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 399.580 3.150 401.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 475.180 3.560 477.380 193.000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 15.380 3.560 17.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 90.980 3.560 93.180 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 166.580 3.560 168.780 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 242.180 3.560 244.380 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 317.780 3.560 319.980 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 393.380 3.560 395.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 468.980 3.560 471.180 193.000 ;
    END
  END VPWR
  PIN analog_adc
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 499.600 165.700 500.000 166.100 ;
    END
  END analog_adc
  PIN analog_pin0
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.654400 ;
    PORT
      LAYER Metal3 ;
        RECT 499.600 32.980 500.000 33.380 ;
    END
  END analog_pin0
  PIN analog_pin1
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.654400 ;
    PORT
      LAYER Metal3 ;
        RECT 499.600 99.340 500.000 99.740 ;
    END
  END analog_pin1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.901600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.340 0.400 183.740 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.140 0.400 179.540 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.540 0.400 187.940 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 111.940 0.400 112.340 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.140 0.400 116.540 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.340 0.400 120.740 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.540 0.400 124.940 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.740 0.400 129.140 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.940 0.400 133.340 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.140 0.400 137.540 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.340 0.400 141.740 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.540 0.400 145.940 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.740 0.400 150.140 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.940 0.400 154.340 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.140 0.400 158.540 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.340 0.400 162.740 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.540 0.400 166.940 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.740 0.400 171.140 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.940 0.400 175.340 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.340 0.400 78.740 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.540 0.400 82.940 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.740 0.400 87.140 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.940 0.400 91.340 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.140 0.400 95.540 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.340 0.400 99.740 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.540 0.400 103.940 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.740 0.400 108.140 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.740 0.400 45.140 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.940 0.400 49.340 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.140 0.400 53.540 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.340 0.400 57.740 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.540 0.400 61.940 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 65.740 0.400 66.140 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.940 0.400 70.340 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.140 0.400 74.540 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.140 0.400 11.540 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.340 0.400 15.740 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.540 0.400 19.940 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.740 0.400 24.140 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.940 0.400 28.340 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.140 0.400 32.540 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.340 0.400 36.740 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.540 0.400 40.940 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 496.800 192.930 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 496.800 193.000 ;
      LAYER Metal2 ;
        RECT 2.775 3.635 494.505 192.925 ;
      LAYER Metal3 ;
        RECT 0.400 188.150 499.825 192.880 ;
        RECT 0.610 187.330 499.825 188.150 ;
        RECT 0.400 183.950 499.825 187.330 ;
        RECT 0.610 183.130 499.825 183.950 ;
        RECT 0.400 179.750 499.825 183.130 ;
        RECT 0.610 178.930 499.825 179.750 ;
        RECT 0.400 175.550 499.825 178.930 ;
        RECT 0.610 174.730 499.825 175.550 ;
        RECT 0.400 171.350 499.825 174.730 ;
        RECT 0.610 170.530 499.825 171.350 ;
        RECT 0.400 167.150 499.825 170.530 ;
        RECT 0.610 166.330 499.825 167.150 ;
        RECT 0.400 166.310 499.825 166.330 ;
        RECT 0.400 165.490 499.390 166.310 ;
        RECT 0.400 162.950 499.825 165.490 ;
        RECT 0.610 162.130 499.825 162.950 ;
        RECT 0.400 158.750 499.825 162.130 ;
        RECT 0.610 157.930 499.825 158.750 ;
        RECT 0.400 154.550 499.825 157.930 ;
        RECT 0.610 153.730 499.825 154.550 ;
        RECT 0.400 150.350 499.825 153.730 ;
        RECT 0.610 149.530 499.825 150.350 ;
        RECT 0.400 146.150 499.825 149.530 ;
        RECT 0.610 145.330 499.825 146.150 ;
        RECT 0.400 141.950 499.825 145.330 ;
        RECT 0.610 141.130 499.825 141.950 ;
        RECT 0.400 137.750 499.825 141.130 ;
        RECT 0.610 136.930 499.825 137.750 ;
        RECT 0.400 133.550 499.825 136.930 ;
        RECT 0.610 132.730 499.825 133.550 ;
        RECT 0.400 129.350 499.825 132.730 ;
        RECT 0.610 128.530 499.825 129.350 ;
        RECT 0.400 125.150 499.825 128.530 ;
        RECT 0.610 124.330 499.825 125.150 ;
        RECT 0.400 120.950 499.825 124.330 ;
        RECT 0.610 120.130 499.825 120.950 ;
        RECT 0.400 116.750 499.825 120.130 ;
        RECT 0.610 115.930 499.825 116.750 ;
        RECT 0.400 112.550 499.825 115.930 ;
        RECT 0.610 111.730 499.825 112.550 ;
        RECT 0.400 108.350 499.825 111.730 ;
        RECT 0.610 107.530 499.825 108.350 ;
        RECT 0.400 104.150 499.825 107.530 ;
        RECT 0.610 103.330 499.825 104.150 ;
        RECT 0.400 99.950 499.825 103.330 ;
        RECT 0.610 99.130 499.390 99.950 ;
        RECT 0.400 95.750 499.825 99.130 ;
        RECT 0.610 94.930 499.825 95.750 ;
        RECT 0.400 91.550 499.825 94.930 ;
        RECT 0.610 90.730 499.825 91.550 ;
        RECT 0.400 87.350 499.825 90.730 ;
        RECT 0.610 86.530 499.825 87.350 ;
        RECT 0.400 83.150 499.825 86.530 ;
        RECT 0.610 82.330 499.825 83.150 ;
        RECT 0.400 78.950 499.825 82.330 ;
        RECT 0.610 78.130 499.825 78.950 ;
        RECT 0.400 74.750 499.825 78.130 ;
        RECT 0.610 73.930 499.825 74.750 ;
        RECT 0.400 70.550 499.825 73.930 ;
        RECT 0.610 69.730 499.825 70.550 ;
        RECT 0.400 66.350 499.825 69.730 ;
        RECT 0.610 65.530 499.825 66.350 ;
        RECT 0.400 62.150 499.825 65.530 ;
        RECT 0.610 61.330 499.825 62.150 ;
        RECT 0.400 57.950 499.825 61.330 ;
        RECT 0.610 57.130 499.825 57.950 ;
        RECT 0.400 53.750 499.825 57.130 ;
        RECT 0.610 52.930 499.825 53.750 ;
        RECT 0.400 49.550 499.825 52.930 ;
        RECT 0.610 48.730 499.825 49.550 ;
        RECT 0.400 45.350 499.825 48.730 ;
        RECT 0.610 44.530 499.825 45.350 ;
        RECT 0.400 41.150 499.825 44.530 ;
        RECT 0.610 40.330 499.825 41.150 ;
        RECT 0.400 36.950 499.825 40.330 ;
        RECT 0.610 36.130 499.825 36.950 ;
        RECT 0.400 33.590 499.825 36.130 ;
        RECT 0.400 32.770 499.390 33.590 ;
        RECT 0.400 32.750 499.825 32.770 ;
        RECT 0.610 31.930 499.825 32.750 ;
        RECT 0.400 28.550 499.825 31.930 ;
        RECT 0.610 27.730 499.825 28.550 ;
        RECT 0.400 24.350 499.825 27.730 ;
        RECT 0.610 23.530 499.825 24.350 ;
        RECT 0.400 20.150 499.825 23.530 ;
        RECT 0.610 19.330 499.825 20.150 ;
        RECT 0.400 15.950 499.825 19.330 ;
        RECT 0.610 15.130 499.825 15.950 ;
        RECT 0.400 11.750 499.825 15.130 ;
        RECT 0.610 10.930 499.825 11.750 ;
        RECT 0.400 3.680 499.825 10.930 ;
      LAYER Metal4 ;
        RECT 4.215 3.635 499.780 192.925 ;
      LAYER Metal5 ;
        RECT 4.175 3.470 495.025 193.090 ;
      LAYER TopMetal1 ;
        RECT 331.420 28.160 337.620 162.940 ;
  END
END heichips25_internal
END LIBRARY

