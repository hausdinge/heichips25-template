magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771642464
<< metal1 >>
rect 576 38576 83328 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 83328 38576
rect 576 38512 83328 38536
rect 643 38156 701 38157
rect 643 38116 652 38156
rect 692 38116 701 38156
rect 643 38115 701 38116
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 576 37820 83328 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 83328 37820
rect 576 37756 83328 37780
rect 576 37064 83328 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 83328 37064
rect 576 37000 83328 37024
rect 576 36308 83328 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 83328 36308
rect 576 36244 83328 36268
rect 12163 35888 12221 35889
rect 12163 35848 12172 35888
rect 12212 35848 12221 35888
rect 12163 35847 12221 35848
rect 12451 35888 12509 35889
rect 12451 35848 12460 35888
rect 12500 35848 12509 35888
rect 12451 35847 12509 35848
rect 13323 35888 13365 35897
rect 13323 35848 13324 35888
rect 13364 35848 13365 35888
rect 13323 35839 13365 35848
rect 576 35552 83328 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 83328 35552
rect 576 35488 83328 35512
rect 32619 35216 32661 35225
rect 32619 35176 32620 35216
rect 32660 35176 32661 35216
rect 32619 35167 32661 35176
rect 32715 35216 32757 35225
rect 32715 35176 32716 35216
rect 32756 35176 32757 35216
rect 32715 35167 32757 35176
rect 32995 35216 33053 35217
rect 32995 35176 33004 35216
rect 33044 35176 33053 35216
rect 32995 35175 33053 35176
rect 33763 35216 33821 35217
rect 33763 35176 33772 35216
rect 33812 35176 33821 35216
rect 33763 35175 33821 35176
rect 34059 35216 34101 35225
rect 34059 35176 34060 35216
rect 34100 35176 34101 35216
rect 34059 35167 34101 35176
rect 34155 35216 34197 35225
rect 34155 35176 34156 35216
rect 34196 35176 34197 35216
rect 34155 35167 34197 35176
rect 50275 35216 50333 35217
rect 50275 35176 50284 35216
rect 50324 35176 50333 35216
rect 50275 35175 50333 35176
rect 15043 35132 15101 35133
rect 15043 35092 15052 35132
rect 15092 35092 15101 35132
rect 15043 35091 15101 35092
rect 82243 35132 82301 35133
rect 82243 35092 82252 35132
rect 82292 35092 82301 35132
rect 82243 35091 82301 35092
rect 15243 34964 15285 34973
rect 15243 34924 15244 34964
rect 15284 34924 15285 34964
rect 15243 34915 15285 34924
rect 32323 34964 32381 34965
rect 32323 34924 32332 34964
rect 32372 34924 32381 34964
rect 32323 34923 32381 34924
rect 34435 34964 34493 34965
rect 34435 34924 34444 34964
rect 34484 34924 34493 34964
rect 34435 34923 34493 34924
rect 82443 34964 82485 34973
rect 82443 34924 82444 34964
rect 82484 34924 82485 34964
rect 82443 34915 82485 34924
rect 576 34796 83328 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 83328 34796
rect 576 34732 83328 34756
rect 22723 34544 22781 34545
rect 22723 34504 22732 34544
rect 22772 34504 22781 34544
rect 22723 34503 22781 34504
rect 28963 34544 29021 34545
rect 28963 34504 28972 34544
rect 29012 34504 29021 34544
rect 28963 34503 29021 34504
rect 34723 34544 34781 34545
rect 34723 34504 34732 34544
rect 34772 34504 34781 34544
rect 34723 34503 34781 34504
rect 38179 34544 38237 34545
rect 38179 34504 38188 34544
rect 38228 34504 38237 34544
rect 38179 34503 38237 34504
rect 49987 34544 50045 34545
rect 49987 34504 49996 34544
rect 50036 34504 50045 34544
rect 49987 34503 50045 34504
rect 50571 34544 50613 34553
rect 50571 34504 50572 34544
rect 50612 34504 50613 34544
rect 50571 34495 50613 34504
rect 52195 34544 52253 34545
rect 52195 34504 52204 34544
rect 52244 34504 52253 34544
rect 52195 34503 52253 34504
rect 83203 34544 83261 34545
rect 83203 34504 83212 34544
rect 83252 34504 83261 34544
rect 83203 34503 83261 34504
rect 20803 34460 20861 34461
rect 20803 34420 20812 34460
rect 20852 34420 20861 34460
rect 20803 34419 20861 34420
rect 21187 34460 21245 34461
rect 21187 34420 21196 34460
rect 21236 34420 21245 34460
rect 21187 34419 21245 34420
rect 21571 34460 21629 34461
rect 21571 34420 21580 34460
rect 21620 34420 21629 34460
rect 21571 34419 21629 34420
rect 22915 34460 22973 34461
rect 22915 34420 22924 34460
rect 22964 34420 22973 34460
rect 22915 34419 22973 34420
rect 45571 34460 45629 34461
rect 45571 34420 45580 34460
rect 45620 34420 45629 34460
rect 45571 34419 45629 34420
rect 15051 34376 15093 34385
rect 15051 34336 15052 34376
rect 15092 34336 15093 34376
rect 15051 34327 15093 34336
rect 15811 34376 15869 34377
rect 15811 34336 15820 34376
rect 15860 34336 15869 34376
rect 15811 34335 15869 34336
rect 16675 34376 16733 34377
rect 16675 34336 16684 34376
rect 16724 34336 16733 34376
rect 16675 34335 16733 34336
rect 18403 34376 18461 34377
rect 18403 34336 18412 34376
rect 18452 34336 18461 34376
rect 18403 34335 18461 34336
rect 19267 34376 19325 34377
rect 19267 34336 19276 34376
rect 19316 34336 19325 34376
rect 19267 34335 19325 34336
rect 22051 34376 22109 34377
rect 22051 34336 22060 34376
rect 22100 34336 22109 34376
rect 22051 34335 22109 34336
rect 22347 34376 22389 34385
rect 22347 34336 22348 34376
rect 22388 34336 22389 34376
rect 22347 34327 22389 34336
rect 29355 34376 29397 34385
rect 29355 34336 29356 34376
rect 29396 34336 29397 34376
rect 29355 34327 29397 34336
rect 29635 34376 29693 34377
rect 29635 34336 29644 34376
rect 29684 34336 29693 34376
rect 29635 34335 29693 34336
rect 32331 34376 32373 34385
rect 32331 34336 32332 34376
rect 32372 34336 32373 34376
rect 32331 34327 32373 34336
rect 32707 34376 32765 34377
rect 32707 34336 32716 34376
rect 32756 34336 32765 34376
rect 32707 34335 32765 34336
rect 33571 34376 33629 34377
rect 33571 34336 33580 34376
rect 33620 34336 33629 34376
rect 33571 34335 33629 34336
rect 36931 34376 36989 34377
rect 36931 34336 36940 34376
rect 36980 34336 36989 34376
rect 36931 34335 36989 34336
rect 37891 34376 37949 34377
rect 37891 34336 37900 34376
rect 37940 34336 37949 34376
rect 37891 34335 37949 34336
rect 38571 34376 38613 34385
rect 38571 34336 38572 34376
rect 38612 34336 38613 34376
rect 38571 34327 38613 34336
rect 38851 34376 38909 34377
rect 38851 34336 38860 34376
rect 38900 34336 38909 34376
rect 38851 34335 38909 34336
rect 49315 34376 49373 34377
rect 49315 34336 49324 34376
rect 49364 34336 49373 34376
rect 49315 34335 49373 34336
rect 49611 34376 49653 34385
rect 49611 34336 49612 34376
rect 49652 34336 49653 34376
rect 49611 34327 49653 34336
rect 50275 34376 50333 34377
rect 50275 34336 50284 34376
rect 50324 34336 50333 34376
rect 50275 34335 50333 34336
rect 51523 34376 51581 34377
rect 51523 34336 51532 34376
rect 51572 34336 51581 34376
rect 51523 34335 51581 34336
rect 51819 34376 51861 34385
rect 51819 34336 51820 34376
rect 51860 34336 51861 34376
rect 51819 34327 51861 34336
rect 81187 34376 81245 34377
rect 81187 34336 81196 34376
rect 81236 34336 81245 34376
rect 81187 34335 81245 34336
rect 82051 34376 82109 34377
rect 82051 34336 82060 34376
rect 82100 34336 82109 34376
rect 82051 34335 82109 34336
rect 15435 34292 15477 34301
rect 15435 34252 15436 34292
rect 15476 34252 15477 34292
rect 15435 34243 15477 34252
rect 18027 34292 18069 34301
rect 18027 34252 18028 34292
rect 18068 34252 18069 34292
rect 18027 34243 18069 34252
rect 22443 34292 22485 34301
rect 22443 34252 22444 34292
rect 22484 34252 22485 34292
rect 22443 34243 22485 34252
rect 29259 34292 29301 34301
rect 29259 34252 29260 34292
rect 29300 34252 29301 34292
rect 29259 34243 29301 34252
rect 38475 34292 38517 34301
rect 38475 34252 38476 34292
rect 38516 34252 38517 34292
rect 38475 34243 38517 34252
rect 49707 34292 49749 34301
rect 49707 34252 49708 34292
rect 49748 34252 49749 34292
rect 49707 34243 49749 34252
rect 51915 34292 51957 34301
rect 51915 34252 51916 34292
rect 51956 34252 51957 34292
rect 51915 34243 51957 34252
rect 80811 34292 80853 34301
rect 80811 34252 80812 34292
rect 80852 34252 80853 34292
rect 80811 34243 80853 34252
rect 14667 34208 14709 34217
rect 14667 34168 14668 34208
rect 14708 34168 14709 34208
rect 14667 34159 14709 34168
rect 17827 34208 17885 34209
rect 17827 34168 17836 34208
rect 17876 34168 17885 34208
rect 17827 34167 17885 34168
rect 20419 34208 20477 34209
rect 20419 34168 20428 34208
rect 20468 34168 20477 34208
rect 20419 34167 20477 34168
rect 21003 34208 21045 34217
rect 21003 34168 21004 34208
rect 21044 34168 21045 34208
rect 21003 34159 21045 34168
rect 21387 34208 21429 34217
rect 21387 34168 21388 34208
rect 21428 34168 21429 34208
rect 21387 34159 21429 34168
rect 21771 34208 21813 34217
rect 21771 34168 21772 34208
rect 21812 34168 21813 34208
rect 21771 34159 21813 34168
rect 23115 34208 23157 34217
rect 23115 34168 23116 34208
rect 23156 34168 23157 34208
rect 23115 34159 23157 34168
rect 45387 34208 45429 34217
rect 45387 34168 45388 34208
rect 45428 34168 45429 34208
rect 45387 34159 45429 34168
rect 50763 34208 50805 34217
rect 50763 34168 50764 34208
rect 50804 34168 50805 34208
rect 50763 34159 50805 34168
rect 576 34040 83328 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 83328 34040
rect 576 33976 83328 34000
rect 29539 33872 29597 33873
rect 29539 33832 29548 33872
rect 29588 33832 29597 33872
rect 29539 33831 29597 33832
rect 40291 33872 40349 33873
rect 40291 33832 40300 33872
rect 40340 33832 40349 33872
rect 40291 33831 40349 33832
rect 52483 33872 52541 33873
rect 52483 33832 52492 33872
rect 52532 33832 52541 33872
rect 52483 33831 52541 33832
rect 17355 33788 17397 33797
rect 17355 33748 17356 33788
rect 17396 33748 17397 33788
rect 17355 33739 17397 33748
rect 21099 33788 21141 33797
rect 21099 33748 21100 33788
rect 21140 33748 21141 33788
rect 21099 33739 21141 33748
rect 25323 33788 25365 33797
rect 25323 33748 25324 33788
rect 25364 33748 25365 33788
rect 25323 33739 25365 33748
rect 37899 33788 37941 33797
rect 37899 33748 37900 33788
rect 37940 33748 37941 33788
rect 37899 33739 37941 33748
rect 50091 33788 50133 33797
rect 50091 33748 50092 33788
rect 50132 33748 50133 33788
rect 50091 33739 50133 33748
rect 81867 33788 81909 33797
rect 81867 33748 81868 33788
rect 81908 33748 81909 33788
rect 81867 33739 81909 33748
rect 13995 33704 14037 33713
rect 13995 33664 13996 33704
rect 14036 33664 14037 33704
rect 13995 33655 14037 33664
rect 14371 33704 14429 33705
rect 14371 33664 14380 33704
rect 14420 33664 14429 33704
rect 14371 33663 14429 33664
rect 15235 33704 15293 33705
rect 15235 33664 15244 33704
rect 15284 33664 15293 33704
rect 15235 33663 15293 33664
rect 16963 33704 17021 33705
rect 16963 33664 16972 33704
rect 17012 33664 17021 33704
rect 20707 33704 20765 33705
rect 16963 33663 17021 33664
rect 17259 33662 17301 33671
rect 20707 33664 20716 33704
rect 20756 33664 20765 33704
rect 20707 33663 20765 33664
rect 21003 33704 21045 33713
rect 21003 33664 21004 33704
rect 21044 33664 21045 33704
rect 17259 33622 17260 33662
rect 17300 33622 17301 33662
rect 21003 33655 21045 33664
rect 21771 33704 21813 33713
rect 21771 33664 21772 33704
rect 21812 33664 21813 33704
rect 21771 33655 21813 33664
rect 22627 33704 22685 33705
rect 22627 33664 22636 33704
rect 22676 33664 22685 33704
rect 22627 33663 22685 33664
rect 24067 33704 24125 33705
rect 24067 33664 24076 33704
rect 24116 33664 24125 33704
rect 24067 33663 24125 33664
rect 24931 33704 24989 33705
rect 24931 33664 24940 33704
rect 24980 33664 24989 33704
rect 24931 33663 24989 33664
rect 25603 33704 25661 33705
rect 25603 33664 25612 33704
rect 25652 33664 25661 33704
rect 25603 33663 25661 33664
rect 26563 33704 26621 33705
rect 26563 33664 26572 33704
rect 26612 33664 26621 33704
rect 26563 33663 26621 33664
rect 27147 33704 27189 33713
rect 27147 33664 27148 33704
rect 27188 33664 27189 33704
rect 27147 33655 27189 33664
rect 27523 33704 27581 33705
rect 27523 33664 27532 33704
rect 27572 33664 27581 33704
rect 27523 33663 27581 33664
rect 28387 33704 28445 33705
rect 28387 33664 28396 33704
rect 28436 33664 28445 33704
rect 28387 33663 28445 33664
rect 30211 33704 30269 33705
rect 30211 33664 30220 33704
rect 30260 33664 30269 33704
rect 30211 33663 30269 33664
rect 30507 33704 30549 33713
rect 30507 33664 30508 33704
rect 30548 33664 30549 33704
rect 30507 33655 30549 33664
rect 30603 33704 30645 33713
rect 30603 33664 30604 33704
rect 30644 33664 30645 33704
rect 30603 33655 30645 33664
rect 31083 33704 31125 33713
rect 31083 33664 31084 33704
rect 31124 33664 31125 33704
rect 31083 33655 31125 33664
rect 31459 33704 31517 33705
rect 31459 33664 31468 33704
rect 31508 33664 31517 33704
rect 31459 33663 31517 33664
rect 32323 33704 32381 33705
rect 32323 33664 32332 33704
rect 32372 33664 32381 33704
rect 32323 33663 32381 33664
rect 33763 33704 33821 33705
rect 33763 33664 33772 33704
rect 33812 33664 33821 33704
rect 33763 33663 33821 33664
rect 34059 33704 34101 33713
rect 34059 33664 34060 33704
rect 34100 33664 34101 33704
rect 34059 33655 34101 33664
rect 34155 33704 34197 33713
rect 34155 33664 34156 33704
rect 34196 33664 34197 33704
rect 34155 33655 34197 33664
rect 35307 33704 35349 33713
rect 35307 33664 35308 33704
rect 35348 33664 35349 33704
rect 35307 33655 35349 33664
rect 35683 33704 35741 33705
rect 35683 33664 35692 33704
rect 35732 33664 35741 33704
rect 35683 33663 35741 33664
rect 36547 33704 36605 33705
rect 36547 33664 36556 33704
rect 36596 33664 36605 33704
rect 36547 33663 36605 33664
rect 38275 33704 38333 33705
rect 38275 33664 38284 33704
rect 38324 33664 38333 33704
rect 38275 33663 38333 33664
rect 39139 33704 39197 33705
rect 39139 33664 39148 33704
rect 39188 33664 39197 33704
rect 39139 33663 39197 33664
rect 41643 33704 41685 33713
rect 41643 33664 41644 33704
rect 41684 33664 41685 33704
rect 41643 33655 41685 33664
rect 42019 33704 42077 33705
rect 42019 33664 42028 33704
rect 42068 33664 42077 33704
rect 42019 33663 42077 33664
rect 42883 33704 42941 33705
rect 42883 33664 42892 33704
rect 42932 33664 42941 33704
rect 42883 33663 42941 33664
rect 44907 33704 44949 33713
rect 44907 33664 44908 33704
rect 44948 33664 44949 33704
rect 44907 33655 44949 33664
rect 45283 33704 45341 33705
rect 45283 33664 45292 33704
rect 45332 33664 45341 33704
rect 45283 33663 45341 33664
rect 46147 33704 46205 33705
rect 46147 33664 46156 33704
rect 46196 33664 46205 33704
rect 46147 33663 46205 33664
rect 47499 33704 47541 33713
rect 47499 33664 47500 33704
rect 47540 33664 47541 33704
rect 47499 33655 47541 33664
rect 47875 33704 47933 33705
rect 47875 33664 47884 33704
rect 47924 33664 47933 33704
rect 47875 33663 47933 33664
rect 48739 33704 48797 33705
rect 48739 33664 48748 33704
rect 48788 33664 48797 33704
rect 48739 33663 48797 33664
rect 50467 33704 50525 33705
rect 50467 33664 50476 33704
rect 50516 33664 50525 33704
rect 50467 33663 50525 33664
rect 51331 33704 51389 33705
rect 51331 33664 51340 33704
rect 51380 33664 51389 33704
rect 51331 33663 51389 33664
rect 52675 33704 52733 33705
rect 52675 33664 52684 33704
rect 52724 33664 52733 33704
rect 52675 33663 52733 33664
rect 81963 33704 82005 33713
rect 81963 33664 81964 33704
rect 82004 33664 82005 33704
rect 81963 33655 82005 33664
rect 82243 33704 82301 33705
rect 82243 33664 82252 33704
rect 82292 33664 82301 33704
rect 82243 33663 82301 33664
rect 17259 33613 17301 33622
rect 33483 33620 33525 33629
rect 33483 33580 33484 33620
rect 33524 33580 33525 33620
rect 33483 33571 33525 33580
rect 17635 33536 17693 33537
rect 17635 33496 17644 33536
rect 17684 33496 17693 33536
rect 17635 33495 17693 33496
rect 30883 33536 30941 33537
rect 30883 33496 30892 33536
rect 30932 33496 30941 33536
rect 30883 33495 30941 33496
rect 34435 33536 34493 33537
rect 34435 33496 34444 33536
rect 34484 33496 34493 33536
rect 34435 33495 34493 33496
rect 81571 33536 81629 33537
rect 81571 33496 81580 33536
rect 81620 33496 81629 33536
rect 81571 33495 81629 33496
rect 16387 33452 16445 33453
rect 16387 33412 16396 33452
rect 16436 33412 16445 33452
rect 16387 33411 16445 33412
rect 21379 33452 21437 33453
rect 21379 33412 21388 33452
rect 21428 33412 21437 33452
rect 21379 33411 21437 33412
rect 21963 33452 22005 33461
rect 21963 33412 21964 33452
rect 22004 33412 22005 33452
rect 21963 33403 22005 33412
rect 22915 33452 22973 33453
rect 22915 33412 22924 33452
rect 22964 33412 22973 33452
rect 22915 33411 22973 33412
rect 29539 33452 29597 33453
rect 29539 33412 29548 33452
rect 29588 33412 29597 33452
rect 29539 33411 29597 33412
rect 37699 33452 37757 33453
rect 37699 33412 37708 33452
rect 37748 33412 37757 33452
rect 37699 33411 37757 33412
rect 44035 33452 44093 33453
rect 44035 33412 44044 33452
rect 44084 33412 44093 33452
rect 44035 33411 44093 33412
rect 47299 33452 47357 33453
rect 47299 33412 47308 33452
rect 47348 33412 47357 33452
rect 47299 33411 47357 33412
rect 49891 33452 49949 33453
rect 49891 33412 49900 33452
rect 49940 33412 49949 33452
rect 49891 33411 49949 33412
rect 52483 33452 52541 33453
rect 52483 33412 52492 33452
rect 52532 33412 52541 33452
rect 52483 33411 52541 33412
rect 576 33284 83328 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 83328 33284
rect 576 33220 83328 33244
rect 12259 33116 12317 33117
rect 12259 33076 12268 33116
rect 12308 33076 12317 33116
rect 12259 33075 12317 33076
rect 14467 33116 14525 33117
rect 14467 33076 14476 33116
rect 14516 33076 14525 33116
rect 14467 33075 14525 33076
rect 15331 33116 15389 33117
rect 15331 33076 15340 33116
rect 15380 33076 15389 33116
rect 15331 33075 15389 33076
rect 20515 33116 20573 33117
rect 20515 33076 20524 33116
rect 20564 33076 20573 33116
rect 20515 33075 20573 33076
rect 23683 33116 23741 33117
rect 23683 33076 23692 33116
rect 23732 33076 23741 33116
rect 23683 33075 23741 33076
rect 27139 33116 27197 33117
rect 27139 33076 27148 33116
rect 27188 33076 27197 33116
rect 27139 33075 27197 33076
rect 31747 33116 31805 33117
rect 31747 33076 31756 33116
rect 31796 33076 31805 33116
rect 31747 33075 31805 33076
rect 36739 33116 36797 33117
rect 36739 33076 36748 33116
rect 36788 33076 36797 33116
rect 36739 33075 36797 33076
rect 41251 33116 41309 33117
rect 41251 33076 41260 33116
rect 41300 33076 41309 33116
rect 41251 33075 41309 33076
rect 42315 33116 42357 33125
rect 42315 33076 42316 33116
rect 42356 33076 42357 33116
rect 42315 33067 42357 33076
rect 45283 33116 45341 33117
rect 45283 33076 45292 33116
rect 45332 33076 45341 33116
rect 45283 33075 45341 33076
rect 47203 33116 47261 33117
rect 47203 33076 47212 33116
rect 47252 33076 47261 33116
rect 47203 33075 47261 33076
rect 9571 33032 9629 33033
rect 9571 32992 9580 33032
rect 9620 32992 9629 33032
rect 9571 32991 9629 32992
rect 17923 33032 17981 33033
rect 17923 32992 17932 33032
rect 17972 32992 17981 33032
rect 17923 32991 17981 32992
rect 43083 33032 43125 33041
rect 43083 32992 43084 33032
rect 43124 32992 43125 33032
rect 43083 32983 43125 32992
rect 69771 33032 69813 33041
rect 69771 32992 69772 33032
rect 69812 32992 69813 33032
rect 69771 32983 69813 32992
rect 42115 32948 42173 32949
rect 42115 32908 42124 32948
rect 42164 32908 42173 32948
rect 42115 32907 42173 32908
rect 5731 32864 5789 32865
rect 5731 32824 5740 32864
rect 5780 32824 5789 32864
rect 5731 32823 5789 32824
rect 6595 32864 6653 32865
rect 6595 32824 6604 32864
rect 6644 32824 6653 32864
rect 6595 32823 6653 32824
rect 8899 32864 8957 32865
rect 8899 32824 8908 32864
rect 8948 32824 8957 32864
rect 8899 32823 8957 32824
rect 9195 32864 9237 32873
rect 9195 32824 9196 32864
rect 9236 32824 9237 32864
rect 9195 32815 9237 32824
rect 9291 32864 9333 32873
rect 9291 32824 9292 32864
rect 9332 32824 9333 32864
rect 9291 32815 9333 32824
rect 9867 32864 9909 32873
rect 9867 32824 9868 32864
rect 9908 32824 9909 32864
rect 9867 32815 9909 32824
rect 10243 32864 10301 32865
rect 10243 32824 10252 32864
rect 10292 32824 10301 32864
rect 10243 32823 10301 32824
rect 11107 32864 11165 32865
rect 11107 32824 11116 32864
rect 11156 32824 11165 32864
rect 11107 32823 11165 32824
rect 13795 32864 13853 32865
rect 13795 32824 13804 32864
rect 13844 32824 13853 32864
rect 13795 32823 13853 32824
rect 14091 32864 14133 32873
rect 14091 32824 14092 32864
rect 14132 32824 14133 32864
rect 14091 32815 14133 32824
rect 15723 32864 15765 32873
rect 15723 32824 15724 32864
rect 15764 32824 15765 32864
rect 15723 32815 15765 32824
rect 16003 32864 16061 32865
rect 16003 32824 16012 32864
rect 16052 32824 16061 32864
rect 16003 32823 16061 32824
rect 17215 32864 17257 32873
rect 17215 32824 17216 32864
rect 17256 32824 17257 32864
rect 17215 32815 17257 32824
rect 17547 32864 17589 32873
rect 17547 32824 17548 32864
rect 17588 32824 17589 32864
rect 17547 32815 17589 32824
rect 17643 32864 17685 32873
rect 17643 32824 17644 32864
rect 17684 32824 17685 32864
rect 17643 32815 17685 32824
rect 18123 32864 18165 32873
rect 18123 32824 18124 32864
rect 18164 32824 18165 32864
rect 18123 32815 18165 32824
rect 18499 32864 18557 32865
rect 18499 32824 18508 32864
rect 18548 32824 18557 32864
rect 18499 32823 18557 32824
rect 19363 32864 19421 32865
rect 19363 32824 19372 32864
rect 19412 32824 19421 32864
rect 19363 32823 19421 32824
rect 21291 32864 21333 32873
rect 21291 32824 21292 32864
rect 21332 32824 21333 32864
rect 21291 32815 21333 32824
rect 21667 32864 21725 32865
rect 21667 32824 21676 32864
rect 21716 32824 21725 32864
rect 21667 32823 21725 32824
rect 22531 32864 22589 32865
rect 22531 32824 22540 32864
rect 22580 32824 22589 32864
rect 22531 32823 22589 32824
rect 25507 32864 25565 32865
rect 25507 32824 25516 32864
rect 25556 32824 25565 32864
rect 25507 32823 25565 32824
rect 27531 32864 27573 32873
rect 27531 32824 27532 32864
rect 27572 32824 27573 32864
rect 27531 32815 27573 32824
rect 27811 32864 27869 32865
rect 27811 32824 27820 32864
rect 27860 32824 27869 32864
rect 27811 32823 27869 32824
rect 29355 32864 29397 32873
rect 29355 32824 29356 32864
rect 29396 32824 29397 32864
rect 29355 32815 29397 32824
rect 29731 32864 29789 32865
rect 29731 32824 29740 32864
rect 29780 32824 29789 32864
rect 29731 32823 29789 32824
rect 30595 32864 30653 32865
rect 30595 32824 30604 32864
rect 30644 32824 30653 32864
rect 30595 32823 30653 32824
rect 33091 32864 33149 32865
rect 33091 32824 33100 32864
rect 33140 32824 33149 32864
rect 33091 32823 33149 32824
rect 33963 32864 34005 32873
rect 33963 32824 33964 32864
rect 34004 32824 34005 32864
rect 33963 32815 34005 32824
rect 34347 32864 34389 32873
rect 34347 32824 34348 32864
rect 34388 32824 34389 32864
rect 34347 32815 34389 32824
rect 34723 32864 34781 32865
rect 34723 32824 34732 32864
rect 34772 32824 34781 32864
rect 34723 32823 34781 32824
rect 35587 32864 35645 32865
rect 35587 32824 35596 32864
rect 35636 32824 35645 32864
rect 35587 32823 35645 32824
rect 36931 32864 36989 32865
rect 36931 32824 36940 32864
rect 36980 32824 36989 32864
rect 36931 32823 36989 32824
rect 37315 32864 37373 32865
rect 37315 32824 37324 32864
rect 37364 32824 37373 32864
rect 37315 32823 37373 32824
rect 38763 32864 38805 32873
rect 38763 32824 38764 32864
rect 38804 32824 38805 32864
rect 38763 32815 38805 32824
rect 40579 32864 40637 32865
rect 40579 32824 40588 32864
rect 40628 32824 40637 32864
rect 40579 32823 40637 32824
rect 40875 32864 40917 32873
rect 40875 32824 40876 32864
rect 40916 32824 40917 32864
rect 40875 32815 40917 32824
rect 40971 32864 41013 32873
rect 40971 32824 40972 32864
rect 41012 32824 41013 32864
rect 40971 32815 41013 32824
rect 44707 32864 44765 32865
rect 44707 32824 44716 32864
rect 44756 32824 44765 32864
rect 44707 32823 44765 32824
rect 45579 32864 45621 32873
rect 45579 32824 45580 32864
rect 45620 32824 45621 32864
rect 45579 32815 45621 32824
rect 45675 32864 45717 32873
rect 45675 32824 45676 32864
rect 45716 32824 45717 32864
rect 45675 32815 45717 32824
rect 45955 32864 46013 32865
rect 45955 32824 45964 32864
rect 46004 32824 46013 32864
rect 45955 32823 46013 32824
rect 47595 32864 47637 32873
rect 47595 32824 47596 32864
rect 47636 32824 47637 32864
rect 47595 32815 47637 32824
rect 47875 32864 47933 32865
rect 47875 32824 47884 32864
rect 47924 32824 47933 32864
rect 47875 32823 47933 32824
rect 49123 32864 49181 32865
rect 49123 32824 49132 32864
rect 49172 32824 49181 32864
rect 49123 32823 49181 32824
rect 50283 32864 50325 32873
rect 50283 32824 50284 32864
rect 50324 32824 50325 32864
rect 50283 32815 50325 32824
rect 50755 32864 50813 32865
rect 50755 32824 50764 32864
rect 50804 32824 50813 32864
rect 50755 32823 50813 32824
rect 51715 32864 51773 32865
rect 51715 32824 51724 32864
rect 51764 32824 51773 32864
rect 51715 32823 51773 32824
rect 51915 32864 51957 32873
rect 51915 32824 51916 32864
rect 51956 32824 51957 32864
rect 51915 32815 51957 32824
rect 52291 32864 52349 32865
rect 52291 32824 52300 32864
rect 52340 32824 52349 32864
rect 52291 32823 52349 32824
rect 53155 32864 53213 32865
rect 53155 32824 53164 32864
rect 53204 32824 53213 32864
rect 53155 32823 53213 32824
rect 64963 32864 65021 32865
rect 64963 32824 64972 32864
rect 65012 32824 65021 32864
rect 64963 32823 65021 32824
rect 65251 32864 65309 32865
rect 65251 32824 65260 32864
rect 65300 32824 65309 32864
rect 65251 32823 65309 32824
rect 66123 32864 66165 32873
rect 66123 32824 66124 32864
rect 66164 32824 66165 32864
rect 66123 32815 66165 32824
rect 70051 32864 70109 32865
rect 70051 32824 70060 32864
rect 70100 32824 70109 32864
rect 70051 32823 70109 32824
rect 5355 32780 5397 32789
rect 5355 32740 5356 32780
rect 5396 32740 5397 32780
rect 5355 32731 5397 32740
rect 14187 32780 14229 32789
rect 14187 32740 14188 32780
rect 14228 32740 14229 32780
rect 14187 32731 14229 32740
rect 15627 32780 15669 32789
rect 15627 32740 15628 32780
rect 15668 32740 15669 32780
rect 15627 32731 15669 32740
rect 27435 32780 27477 32789
rect 27435 32740 27436 32780
rect 27476 32740 27477 32780
rect 27435 32731 27477 32740
rect 47499 32780 47541 32789
rect 47499 32740 47500 32780
rect 47540 32740 47541 32780
rect 47499 32731 47541 32740
rect 7747 32696 7805 32697
rect 7747 32656 7756 32696
rect 7796 32656 7805 32696
rect 7747 32655 7805 32656
rect 12259 32696 12317 32697
rect 12259 32656 12268 32696
rect 12308 32656 12317 32696
rect 12259 32655 12317 32656
rect 23683 32696 23741 32697
rect 23683 32656 23692 32696
rect 23732 32656 23741 32696
rect 23683 32655 23741 32656
rect 31747 32696 31805 32697
rect 31747 32656 31756 32696
rect 31796 32656 31805 32696
rect 31747 32655 31805 32656
rect 42699 32696 42741 32705
rect 42699 32656 42700 32696
rect 42740 32656 42741 32696
rect 42699 32647 42741 32656
rect 48651 32696 48693 32705
rect 48651 32656 48652 32696
rect 48692 32656 48693 32696
rect 48651 32647 48693 32656
rect 49899 32696 49941 32705
rect 49899 32656 49900 32696
rect 49940 32656 49941 32696
rect 49899 32647 49941 32656
rect 54307 32696 54365 32697
rect 54307 32656 54316 32696
rect 54356 32656 54365 32696
rect 54307 32655 54365 32656
rect 65739 32696 65781 32705
rect 65739 32656 65740 32696
rect 65780 32656 65781 32696
rect 65739 32647 65781 32656
rect 576 32528 83328 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 83328 32528
rect 576 32464 83328 32488
rect 80811 32192 80853 32201
rect 80811 32152 80812 32192
rect 80852 32152 80853 32192
rect 80811 32143 80853 32152
rect 81187 32192 81245 32193
rect 81187 32152 81196 32192
rect 81236 32152 81245 32192
rect 81187 32151 81245 32152
rect 82051 32192 82109 32193
rect 82051 32152 82060 32192
rect 82100 32152 82109 32192
rect 82051 32151 82109 32152
rect 1891 32108 1949 32109
rect 1891 32068 1900 32108
rect 1940 32068 1949 32108
rect 1891 32067 1949 32068
rect 83203 32024 83261 32025
rect 83203 31984 83212 32024
rect 83252 31984 83261 32024
rect 83203 31983 83261 31984
rect 2091 31940 2133 31949
rect 2091 31900 2092 31940
rect 2132 31900 2133 31940
rect 2091 31891 2133 31900
rect 576 31772 5952 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 5952 31772
rect 576 31708 5952 31732
rect 74016 31772 83328 31796
rect 74016 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 83328 31772
rect 74016 31708 83328 31732
rect 1515 31604 1557 31613
rect 1515 31564 1516 31604
rect 1556 31564 1557 31604
rect 1515 31555 1557 31564
rect 4963 31604 5021 31605
rect 4963 31564 4972 31604
rect 5012 31564 5021 31604
rect 4963 31563 5021 31564
rect 81379 31604 81437 31605
rect 81379 31564 81388 31604
rect 81428 31564 81437 31604
rect 81379 31563 81437 31564
rect 1899 31520 1941 31529
rect 1899 31480 1900 31520
rect 1940 31480 1941 31520
rect 1899 31471 1941 31480
rect 1315 31436 1373 31437
rect 1315 31396 1324 31436
rect 1364 31396 1373 31436
rect 1315 31395 1373 31396
rect 1699 31436 1757 31437
rect 1699 31396 1708 31436
rect 1748 31396 1757 31436
rect 1699 31395 1757 31396
rect 2755 31352 2813 31353
rect 2755 31312 2764 31352
rect 2804 31312 2813 31352
rect 2755 31311 2813 31312
rect 3619 31352 3677 31353
rect 3619 31312 3628 31352
rect 3668 31312 3677 31352
rect 3619 31311 3677 31312
rect 5259 31352 5301 31361
rect 5259 31312 5260 31352
rect 5300 31312 5301 31352
rect 5259 31303 5301 31312
rect 5355 31348 5397 31357
rect 5355 31308 5356 31348
rect 5396 31308 5397 31348
rect 5671 31352 5729 31353
rect 5671 31312 5680 31352
rect 5720 31312 5729 31352
rect 5671 31311 5729 31312
rect 81675 31352 81717 31361
rect 81675 31312 81676 31352
rect 81716 31312 81717 31352
rect 5355 31299 5397 31308
rect 81675 31303 81717 31312
rect 81771 31352 81813 31361
rect 81771 31312 81772 31352
rect 81812 31312 81813 31352
rect 81771 31303 81813 31312
rect 82051 31352 82109 31353
rect 82051 31312 82060 31352
rect 82100 31312 82109 31352
rect 82051 31311 82109 31312
rect 2379 31268 2421 31277
rect 2379 31228 2380 31268
rect 2420 31228 2421 31268
rect 2379 31219 2421 31228
rect 4771 31184 4829 31185
rect 4771 31144 4780 31184
rect 4820 31144 4829 31184
rect 4771 31143 4829 31144
rect 576 31016 5952 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 5952 31016
rect 576 30952 5952 30976
rect 74016 31016 83328 31040
rect 74016 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 83328 31016
rect 74016 30952 83328 30976
rect 1227 30680 1269 30689
rect 1227 30640 1228 30680
rect 1268 30640 1269 30680
rect 1227 30631 1269 30640
rect 1603 30680 1661 30681
rect 1603 30640 1612 30680
rect 1652 30640 1661 30680
rect 1603 30639 1661 30640
rect 2467 30680 2525 30681
rect 2467 30640 2476 30680
rect 2516 30640 2525 30680
rect 2467 30639 2525 30640
rect 78307 30680 78365 30681
rect 78307 30640 78316 30680
rect 78356 30640 78365 30680
rect 78307 30639 78365 30640
rect 78699 30680 78741 30689
rect 78699 30640 78700 30680
rect 78740 30640 78741 30680
rect 78699 30631 78741 30640
rect 81859 30680 81917 30681
rect 81859 30640 81868 30680
rect 81908 30640 81917 30680
rect 81859 30639 81917 30640
rect 82243 30680 82301 30681
rect 82243 30640 82252 30680
rect 82292 30640 82301 30680
rect 82243 30639 82301 30640
rect 82539 30512 82581 30521
rect 82539 30472 82540 30512
rect 82580 30472 82581 30512
rect 82539 30463 82581 30472
rect 3619 30428 3677 30429
rect 3619 30388 3628 30428
rect 3668 30388 3677 30428
rect 3619 30387 3677 30388
rect 78891 30428 78933 30437
rect 78891 30388 78892 30428
rect 78932 30388 78933 30428
rect 78891 30379 78933 30388
rect 576 30260 5952 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 5952 30260
rect 576 30196 5952 30220
rect 74016 30260 83328 30284
rect 74016 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 83328 30260
rect 74016 30196 83328 30220
rect 1891 30092 1949 30093
rect 1891 30052 1900 30092
rect 1940 30052 1949 30092
rect 1891 30051 1949 30052
rect 2091 29924 2133 29933
rect 2091 29884 2092 29924
rect 2132 29884 2133 29924
rect 2091 29875 2133 29884
rect 1219 29840 1277 29841
rect 1219 29800 1228 29840
rect 1268 29800 1277 29840
rect 1219 29799 1277 29800
rect 1515 29840 1557 29849
rect 1515 29800 1516 29840
rect 1556 29800 1557 29840
rect 1515 29791 1557 29800
rect 2179 29840 2237 29841
rect 2179 29800 2188 29840
rect 2228 29800 2237 29840
rect 2179 29799 2237 29800
rect 2379 29840 2421 29849
rect 2379 29800 2380 29840
rect 2420 29800 2421 29840
rect 2379 29791 2421 29800
rect 2475 29840 2517 29849
rect 2475 29800 2476 29840
rect 2516 29800 2517 29840
rect 2475 29791 2517 29800
rect 2571 29840 2613 29849
rect 2571 29800 2572 29840
rect 2612 29800 2613 29840
rect 2571 29791 2613 29800
rect 2667 29840 2709 29849
rect 2667 29800 2668 29840
rect 2708 29800 2709 29840
rect 2667 29791 2709 29800
rect 3811 29840 3869 29841
rect 3811 29800 3820 29840
rect 3860 29800 3869 29840
rect 3811 29799 3869 29800
rect 4675 29840 4733 29841
rect 4675 29800 4684 29840
rect 4724 29800 4733 29840
rect 4675 29799 4733 29800
rect 1611 29756 1653 29765
rect 1611 29716 1612 29756
rect 1652 29716 1653 29756
rect 1611 29707 1653 29716
rect 3435 29756 3477 29765
rect 3435 29716 3436 29756
rect 3476 29716 3477 29756
rect 3435 29707 3477 29716
rect 5827 29672 5885 29673
rect 5827 29632 5836 29672
rect 5876 29632 5885 29672
rect 5827 29631 5885 29632
rect 576 29504 5952 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 5952 29504
rect 576 29440 5952 29464
rect 74016 29504 83328 29528
rect 74016 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 83328 29504
rect 74016 29440 83328 29464
rect 2667 29336 2709 29345
rect 2667 29296 2668 29336
rect 2708 29296 2709 29336
rect 2667 29287 2709 29296
rect 2755 29336 2813 29337
rect 2755 29296 2764 29336
rect 2804 29296 2813 29336
rect 2755 29295 2813 29296
rect 3523 29336 3581 29337
rect 3523 29296 3532 29336
rect 3572 29296 3581 29336
rect 3523 29295 3581 29296
rect 3811 29336 3869 29337
rect 3811 29296 3820 29336
rect 3860 29296 3869 29336
rect 3811 29295 3869 29296
rect 2851 29252 2909 29253
rect 2851 29212 2860 29252
rect 2900 29212 2909 29252
rect 2851 29211 2909 29212
rect 1515 29168 1557 29177
rect 1515 29128 1516 29168
rect 1556 29128 1557 29168
rect 1515 29119 1557 29128
rect 1707 29168 1749 29177
rect 1707 29128 1708 29168
rect 1748 29128 1749 29168
rect 1707 29119 1749 29128
rect 1899 29168 1941 29177
rect 1899 29128 1900 29168
rect 1940 29128 1941 29168
rect 1899 29119 1941 29128
rect 2091 29168 2133 29177
rect 2091 29128 2092 29168
rect 2132 29128 2133 29168
rect 2091 29119 2133 29128
rect 2179 29168 2237 29169
rect 2179 29128 2188 29168
rect 2228 29128 2237 29168
rect 2179 29127 2237 29128
rect 2955 29168 2997 29177
rect 2955 29128 2956 29168
rect 2996 29128 2997 29168
rect 2955 29119 2997 29128
rect 3051 29168 3093 29177
rect 3051 29128 3052 29168
rect 3092 29128 3093 29168
rect 3051 29119 3093 29128
rect 3331 29168 3389 29169
rect 3331 29128 3340 29168
rect 3380 29128 3389 29168
rect 3331 29127 3389 29128
rect 3435 29168 3477 29177
rect 3435 29128 3436 29168
rect 3476 29128 3477 29168
rect 3435 29119 3477 29128
rect 3627 29168 3669 29177
rect 3627 29128 3628 29168
rect 3668 29128 3669 29168
rect 3627 29119 3669 29128
rect 3907 29168 3965 29169
rect 3907 29128 3916 29168
rect 3956 29128 3965 29168
rect 3907 29127 3965 29128
rect 4579 29168 4637 29169
rect 4579 29128 4588 29168
rect 4628 29128 4637 29168
rect 4579 29127 4637 29128
rect 4771 29168 4829 29169
rect 4771 29128 4780 29168
rect 4820 29128 4829 29168
rect 4771 29127 4829 29128
rect 5643 29168 5685 29177
rect 5643 29128 5644 29168
rect 5684 29128 5685 29168
rect 5643 29119 5685 29128
rect 1899 29000 1941 29009
rect 1899 28960 1900 29000
rect 1940 28960 1941 29000
rect 1899 28951 1941 28960
rect 1515 28916 1557 28925
rect 1515 28876 1516 28916
rect 1556 28876 1557 28916
rect 1515 28867 1557 28876
rect 4099 28916 4157 28917
rect 4099 28876 4108 28916
rect 4148 28876 4157 28916
rect 4099 28875 4157 28876
rect 5067 28916 5109 28925
rect 5067 28876 5068 28916
rect 5108 28876 5109 28916
rect 5067 28867 5109 28876
rect 576 28748 5952 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 5952 28748
rect 576 28684 5952 28708
rect 74016 28748 83328 28772
rect 74016 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 83328 28748
rect 74016 28684 83328 28708
rect 3139 28580 3197 28581
rect 3139 28540 3148 28580
rect 3188 28540 3197 28580
rect 3139 28539 3197 28540
rect 3907 28496 3965 28497
rect 3907 28456 3916 28496
rect 3956 28456 3965 28496
rect 3907 28455 3965 28456
rect 747 28328 789 28337
rect 747 28288 748 28328
rect 788 28288 789 28328
rect 747 28279 789 28288
rect 1123 28328 1181 28329
rect 1123 28288 1132 28328
rect 1172 28288 1181 28328
rect 1123 28287 1181 28288
rect 1987 28328 2045 28329
rect 1987 28288 1996 28328
rect 2036 28288 2045 28328
rect 1987 28287 2045 28288
rect 3435 28328 3477 28337
rect 3435 28288 3436 28328
rect 3476 28288 3477 28328
rect 3435 28279 3477 28288
rect 3531 28328 3573 28337
rect 3531 28288 3532 28328
rect 3572 28288 3573 28328
rect 3531 28279 3573 28288
rect 3627 28328 3669 28337
rect 3627 28288 3628 28328
rect 3668 28288 3669 28328
rect 3627 28279 3669 28288
rect 3723 28328 3765 28337
rect 3723 28288 3724 28328
rect 3764 28288 3765 28328
rect 3723 28279 3765 28288
rect 4107 28328 4149 28337
rect 4107 28288 4108 28328
rect 4148 28288 4149 28328
rect 4107 28279 4149 28288
rect 4299 28328 4341 28337
rect 4299 28288 4300 28328
rect 4340 28288 4341 28328
rect 4299 28279 4341 28288
rect 4579 28328 4637 28329
rect 4579 28288 4588 28328
rect 4628 28288 4637 28328
rect 4579 28287 4637 28288
rect 4771 28328 4829 28329
rect 4771 28288 4780 28328
rect 4820 28288 4829 28328
rect 4771 28287 4829 28288
rect 5643 28328 5685 28337
rect 5643 28288 5644 28328
rect 5684 28288 5685 28328
rect 5643 28279 5685 28288
rect 4203 28160 4245 28169
rect 4203 28120 4204 28160
rect 4244 28120 4245 28160
rect 4203 28111 4245 28120
rect 4491 28160 4533 28169
rect 4491 28120 4492 28160
rect 4532 28120 4533 28160
rect 4491 28111 4533 28120
rect 576 27992 5952 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 5952 27992
rect 576 27928 5952 27952
rect 74016 27992 83328 28016
rect 74016 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 83328 27992
rect 74016 27928 83328 27952
rect 2083 27824 2141 27825
rect 2083 27784 2092 27824
rect 2132 27784 2141 27824
rect 2083 27783 2141 27784
rect 2755 27824 2813 27825
rect 2755 27784 2764 27824
rect 2804 27784 2813 27824
rect 2755 27783 2813 27784
rect 83203 27824 83261 27825
rect 83203 27784 83212 27824
rect 83252 27784 83261 27824
rect 83203 27783 83261 27784
rect 1795 27740 1853 27741
rect 1795 27700 1804 27740
rect 1844 27700 1853 27740
rect 1795 27699 1853 27700
rect 1995 27656 2037 27665
rect 1995 27616 1996 27656
rect 2036 27616 2037 27656
rect 1995 27607 2037 27616
rect 2091 27656 2133 27665
rect 2091 27616 2092 27656
rect 2132 27616 2133 27656
rect 2091 27607 2133 27616
rect 2851 27656 2909 27657
rect 2851 27616 2860 27656
rect 2900 27616 2909 27656
rect 2851 27615 2909 27616
rect 4579 27656 4637 27657
rect 4579 27616 4588 27656
rect 4628 27616 4637 27656
rect 4579 27615 4637 27616
rect 5443 27656 5501 27657
rect 5443 27616 5452 27656
rect 5492 27616 5501 27656
rect 5443 27615 5501 27616
rect 5835 27656 5877 27665
rect 5835 27616 5836 27656
rect 5876 27616 5877 27656
rect 5835 27607 5877 27616
rect 80811 27656 80853 27665
rect 80811 27616 80812 27656
rect 80852 27616 80853 27656
rect 80811 27607 80853 27616
rect 81187 27656 81245 27657
rect 81187 27616 81196 27656
rect 81236 27616 81245 27656
rect 81187 27615 81245 27616
rect 82051 27656 82109 27657
rect 82051 27616 82060 27656
rect 82100 27616 82109 27656
rect 82051 27615 82109 27616
rect 3435 27572 3477 27581
rect 3435 27532 3436 27572
rect 3476 27532 3477 27572
rect 3435 27523 3477 27532
rect 3043 27488 3101 27489
rect 3043 27448 3052 27488
rect 3092 27448 3101 27488
rect 3043 27447 3101 27448
rect 576 27236 5952 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 5952 27236
rect 576 27172 5952 27196
rect 74016 27236 83328 27260
rect 74016 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 83328 27236
rect 74016 27172 83328 27196
rect 4683 27068 4725 27077
rect 4683 27028 4684 27068
rect 4724 27028 4725 27068
rect 4683 27019 4725 27028
rect 81379 27068 81437 27069
rect 81379 27028 81388 27068
rect 81428 27028 81437 27068
rect 81379 27027 81437 27028
rect 4099 26984 4157 26985
rect 4099 26944 4108 26984
rect 4148 26944 4157 26984
rect 4099 26943 4157 26944
rect 1027 26900 1085 26901
rect 1027 26860 1036 26900
rect 1076 26860 1085 26900
rect 1027 26859 1085 26860
rect 1411 26816 1469 26817
rect 1411 26776 1420 26816
rect 1460 26776 1469 26816
rect 1411 26775 1469 26776
rect 1515 26816 1557 26825
rect 1515 26776 1516 26816
rect 1556 26776 1557 26816
rect 1515 26767 1557 26776
rect 1707 26816 1749 26825
rect 1707 26776 1708 26816
rect 1748 26776 1749 26816
rect 1707 26767 1749 26776
rect 2379 26816 2421 26825
rect 2379 26776 2380 26816
rect 2420 26776 2421 26816
rect 2379 26767 2421 26776
rect 2667 26816 2709 26825
rect 2667 26776 2668 26816
rect 2708 26776 2709 26816
rect 2667 26767 2709 26776
rect 3339 26816 3381 26825
rect 3339 26776 3340 26816
rect 3380 26776 3381 26816
rect 3339 26767 3381 26776
rect 3435 26816 3477 26825
rect 3435 26776 3436 26816
rect 3476 26776 3477 26816
rect 3435 26767 3477 26776
rect 3531 26816 3573 26825
rect 3531 26776 3532 26816
rect 3572 26776 3573 26816
rect 3531 26767 3573 26776
rect 3627 26816 3669 26825
rect 3627 26776 3628 26816
rect 3668 26776 3669 26816
rect 3627 26767 3669 26776
rect 4003 26816 4061 26817
rect 4003 26776 4012 26816
rect 4052 26776 4061 26816
rect 4003 26775 4061 26776
rect 4107 26816 4149 26825
rect 4107 26776 4108 26816
rect 4148 26776 4149 26816
rect 4107 26767 4149 26776
rect 4291 26816 4349 26817
rect 4291 26776 4300 26816
rect 4340 26776 4349 26816
rect 4291 26775 4349 26776
rect 4491 26816 4533 26825
rect 4491 26776 4492 26816
rect 4532 26776 4533 26816
rect 4491 26767 4533 26776
rect 4683 26816 4725 26825
rect 4683 26776 4684 26816
rect 4724 26776 4725 26816
rect 4683 26767 4725 26776
rect 81675 26816 81717 26825
rect 81675 26776 81676 26816
rect 81716 26776 81717 26816
rect 81675 26767 81717 26776
rect 81771 26816 81813 26825
rect 81771 26776 81772 26816
rect 81812 26776 81813 26816
rect 81771 26767 81813 26776
rect 82051 26816 82109 26817
rect 82051 26776 82060 26816
rect 82100 26776 82109 26816
rect 82051 26775 82109 26776
rect 1227 26648 1269 26657
rect 1227 26608 1228 26648
rect 1268 26608 1269 26648
rect 1227 26599 1269 26608
rect 1603 26648 1661 26649
rect 1603 26608 1612 26648
rect 1652 26608 1661 26648
rect 1603 26607 1661 26608
rect 2571 26648 2613 26657
rect 2571 26608 2572 26648
rect 2612 26608 2613 26648
rect 2571 26599 2613 26608
rect 3811 26648 3869 26649
rect 3811 26608 3820 26648
rect 3860 26608 3869 26648
rect 3811 26607 3869 26608
rect 576 26480 5952 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 5952 26480
rect 576 26416 5952 26440
rect 74016 26480 83328 26504
rect 74016 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 83328 26480
rect 74016 26416 83328 26440
rect 3043 26312 3101 26313
rect 3043 26272 3052 26312
rect 3092 26272 3101 26312
rect 3043 26271 3101 26272
rect 3331 26312 3389 26313
rect 3331 26272 3340 26312
rect 3380 26272 3389 26312
rect 3331 26271 3389 26272
rect 651 26228 693 26237
rect 651 26188 652 26228
rect 692 26188 693 26228
rect 651 26179 693 26188
rect 3427 26228 3485 26229
rect 3427 26188 3436 26228
rect 3476 26188 3485 26228
rect 3427 26187 3485 26188
rect 1027 26144 1085 26145
rect 1027 26104 1036 26144
rect 1076 26104 1085 26144
rect 1027 26103 1085 26104
rect 1891 26144 1949 26145
rect 1891 26104 1900 26144
rect 1940 26104 1949 26144
rect 1891 26103 1949 26104
rect 3531 26144 3573 26153
rect 3531 26104 3532 26144
rect 3572 26104 3573 26144
rect 3531 26095 3573 26104
rect 3627 26144 3669 26153
rect 3627 26104 3628 26144
rect 3668 26104 3669 26144
rect 3627 26095 3669 26104
rect 3819 26144 3861 26153
rect 3819 26104 3820 26144
rect 3860 26104 3861 26144
rect 3819 26095 3861 26104
rect 3915 26144 3957 26153
rect 3915 26104 3916 26144
rect 3956 26104 3957 26144
rect 3915 26095 3957 26104
rect 4107 26144 4149 26153
rect 4107 26104 4108 26144
rect 4148 26104 4149 26144
rect 4107 26095 4149 26104
rect 4299 26144 4341 26153
rect 4299 26104 4300 26144
rect 4340 26104 4341 26144
rect 4299 26095 4341 26104
rect 4491 26144 4533 26153
rect 4491 26104 4492 26144
rect 4532 26104 4533 26144
rect 4491 26095 4533 26104
rect 4683 26144 4725 26153
rect 4683 26104 4684 26144
rect 4724 26104 4725 26144
rect 4683 26095 4725 26104
rect 4875 26144 4917 26153
rect 4875 26104 4876 26144
rect 4916 26104 4917 26144
rect 4875 26095 4917 26104
rect 3339 25976 3381 25985
rect 3339 25936 3340 25976
rect 3380 25936 3381 25976
rect 3339 25927 3381 25936
rect 3907 25976 3965 25977
rect 3907 25936 3916 25976
rect 3956 25936 3965 25976
rect 3907 25935 3965 25936
rect 4299 25892 4341 25901
rect 4299 25852 4300 25892
rect 4340 25852 4341 25892
rect 4299 25843 4341 25852
rect 4875 25892 4917 25901
rect 4875 25852 4876 25892
rect 4916 25852 4917 25892
rect 4875 25843 4917 25852
rect 576 25724 5952 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 5952 25724
rect 576 25660 5952 25684
rect 74016 25724 83328 25748
rect 74016 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 83328 25724
rect 74016 25660 83328 25684
rect 1707 25556 1749 25565
rect 1707 25516 1708 25556
rect 1748 25516 1749 25556
rect 1707 25507 1749 25516
rect 643 25388 701 25389
rect 643 25348 652 25388
rect 692 25348 701 25388
rect 643 25347 701 25348
rect 1707 25304 1749 25313
rect 1707 25264 1708 25304
rect 1748 25264 1749 25304
rect 1707 25255 1749 25264
rect 1899 25304 1941 25313
rect 1899 25264 1900 25304
rect 1940 25264 1941 25304
rect 1899 25255 1941 25264
rect 1987 25304 2045 25305
rect 1987 25264 1996 25304
rect 2036 25264 2045 25304
rect 1987 25263 2045 25264
rect 3811 25304 3869 25305
rect 3811 25264 3820 25304
rect 3860 25264 3869 25304
rect 3811 25263 3869 25264
rect 4675 25304 4733 25305
rect 4675 25264 4684 25304
rect 4724 25264 4733 25304
rect 4675 25263 4733 25264
rect 3435 25220 3477 25229
rect 3435 25180 3436 25220
rect 3476 25180 3477 25220
rect 3435 25171 3477 25180
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 5827 25136 5885 25137
rect 5827 25096 5836 25136
rect 5876 25096 5885 25136
rect 5827 25095 5885 25096
rect 576 24968 5952 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 5952 24968
rect 576 24904 5952 24928
rect 74016 24968 83328 24992
rect 74016 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 83328 24968
rect 74016 24904 83328 24928
rect 843 24800 885 24809
rect 843 24760 844 24800
rect 884 24760 885 24800
rect 843 24751 885 24760
rect 4299 24800 4341 24809
rect 4299 24760 4300 24800
rect 4340 24760 4341 24800
rect 4299 24751 4341 24760
rect 3235 24716 3293 24717
rect 3235 24676 3244 24716
rect 3284 24676 3293 24716
rect 3235 24675 3293 24676
rect 2179 24632 2237 24633
rect 2179 24592 2188 24632
rect 2228 24592 2237 24632
rect 2179 24591 2237 24592
rect 3331 24632 3389 24633
rect 3331 24592 3340 24632
rect 3380 24592 3389 24632
rect 3331 24591 3389 24592
rect 3715 24632 3773 24633
rect 3715 24592 3724 24632
rect 3764 24592 3773 24632
rect 3715 24591 3773 24592
rect 3915 24632 3957 24641
rect 3915 24592 3916 24632
rect 3956 24592 3957 24632
rect 3915 24583 3957 24592
rect 4107 24632 4149 24641
rect 4107 24592 4108 24632
rect 4148 24592 4149 24632
rect 4107 24583 4149 24592
rect 4387 24632 4445 24633
rect 4387 24592 4396 24632
rect 4436 24592 4445 24632
rect 4387 24591 4445 24592
rect 79747 24632 79805 24633
rect 79747 24592 79756 24632
rect 79796 24592 79805 24632
rect 79747 24591 79805 24592
rect 643 24548 701 24549
rect 643 24508 652 24548
rect 692 24508 701 24548
rect 643 24507 701 24508
rect 1027 24548 1085 24549
rect 1027 24508 1036 24548
rect 1076 24508 1085 24548
rect 1027 24507 1085 24508
rect 81763 24548 81821 24549
rect 81763 24508 81772 24548
rect 81812 24508 81821 24548
rect 81763 24507 81821 24508
rect 4107 24464 4149 24473
rect 4107 24424 4108 24464
rect 4148 24424 4149 24464
rect 4107 24415 4149 24424
rect 1227 24380 1269 24389
rect 1227 24340 1228 24380
rect 1268 24340 1269 24380
rect 1227 24331 1269 24340
rect 2091 24380 2133 24389
rect 2091 24340 2092 24380
rect 2132 24340 2133 24380
rect 2091 24331 2133 24340
rect 576 24212 5952 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 5952 24212
rect 576 24148 5952 24172
rect 74016 24212 83328 24236
rect 74016 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 83328 24212
rect 74016 24148 83328 24172
rect 5251 24044 5309 24045
rect 5251 24004 5260 24044
rect 5300 24004 5309 24044
rect 5251 24003 5309 24004
rect 1323 23960 1365 23969
rect 1323 23920 1324 23960
rect 1364 23920 1365 23960
rect 1323 23911 1365 23920
rect 2859 23834 2901 23843
rect 843 23792 885 23801
rect 843 23752 844 23792
rect 884 23752 885 23792
rect 843 23743 885 23752
rect 1035 23792 1077 23801
rect 1035 23752 1036 23792
rect 1076 23752 1077 23792
rect 1035 23743 1077 23752
rect 1131 23785 1173 23794
rect 1131 23745 1132 23785
rect 1172 23745 1173 23785
rect 1131 23736 1173 23745
rect 1611 23792 1653 23801
rect 1611 23752 1612 23792
rect 1652 23752 1653 23792
rect 1611 23743 1653 23752
rect 1699 23792 1757 23793
rect 1699 23752 1708 23792
rect 1748 23752 1757 23792
rect 1699 23751 1757 23752
rect 1995 23792 2037 23801
rect 1995 23752 1996 23792
rect 2036 23752 2037 23792
rect 1995 23743 2037 23752
rect 2091 23792 2133 23801
rect 2091 23752 2092 23792
rect 2132 23752 2133 23792
rect 2859 23794 2860 23834
rect 2900 23794 2901 23834
rect 2859 23785 2901 23794
rect 3235 23792 3293 23793
rect 2091 23743 2133 23752
rect 3235 23752 3244 23792
rect 3284 23752 3293 23792
rect 3235 23751 3293 23752
rect 4099 23792 4157 23793
rect 4099 23752 4108 23792
rect 4148 23752 4157 23792
rect 4099 23751 4157 23752
rect 1803 23620 1845 23629
rect 1803 23580 1804 23620
rect 1844 23580 1845 23620
rect 2275 23624 2333 23625
rect 2275 23584 2284 23624
rect 2324 23584 2333 23624
rect 2275 23583 2333 23584
rect 1803 23571 1845 23580
rect 576 23456 5952 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 5952 23456
rect 576 23392 5952 23416
rect 74016 23456 83328 23480
rect 74016 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 83328 23456
rect 74016 23392 83328 23416
rect 3043 23288 3101 23289
rect 3043 23248 3052 23288
rect 3092 23248 3101 23288
rect 3043 23247 3101 23248
rect 4395 23288 4437 23297
rect 4395 23248 4396 23288
rect 4436 23248 4437 23288
rect 4395 23239 4437 23248
rect 651 23120 693 23129
rect 651 23080 652 23120
rect 692 23080 693 23120
rect 651 23071 693 23080
rect 1027 23120 1085 23121
rect 1027 23080 1036 23120
rect 1076 23080 1085 23120
rect 1027 23079 1085 23080
rect 1891 23120 1949 23121
rect 1891 23080 1900 23120
rect 1940 23080 1949 23120
rect 1891 23079 1949 23080
rect 4195 23036 4253 23037
rect 4195 22996 4204 23036
rect 4244 22996 4253 23036
rect 4195 22995 4253 22996
rect 4579 23036 4637 23037
rect 4579 22996 4588 23036
rect 4628 22996 4637 23036
rect 4579 22995 4637 22996
rect 4779 22868 4821 22877
rect 4779 22828 4780 22868
rect 4820 22828 4821 22868
rect 4779 22819 4821 22828
rect 576 22700 5952 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 5952 22700
rect 576 22636 5952 22660
rect 74016 22700 83328 22724
rect 74016 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 83328 22700
rect 74016 22636 83328 22660
rect 1227 22532 1269 22541
rect 1227 22492 1228 22532
rect 1268 22492 1269 22532
rect 1227 22483 1269 22492
rect 1027 22364 1085 22365
rect 1027 22324 1036 22364
rect 1076 22324 1085 22364
rect 1027 22323 1085 22324
rect 3811 22280 3869 22281
rect 3811 22240 3820 22280
rect 3860 22240 3869 22280
rect 3811 22239 3869 22240
rect 4675 22280 4733 22281
rect 4675 22240 4684 22280
rect 4724 22240 4733 22280
rect 4675 22239 4733 22240
rect 3435 22196 3477 22205
rect 3435 22156 3436 22196
rect 3476 22156 3477 22196
rect 3435 22147 3477 22156
rect 643 22112 701 22113
rect 643 22072 652 22112
rect 692 22072 701 22112
rect 643 22071 701 22072
rect 5827 22112 5885 22113
rect 5827 22072 5836 22112
rect 5876 22072 5885 22112
rect 5827 22071 5885 22072
rect 576 21944 5952 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 5952 21944
rect 576 21880 5952 21904
rect 74016 21944 99360 21968
rect 74016 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 74016 21880 99360 21904
rect 4299 21692 4341 21701
rect 4299 21652 4300 21692
rect 4340 21652 4341 21692
rect 4299 21643 4341 21652
rect 4395 21608 4437 21617
rect 4395 21568 4396 21608
rect 4436 21568 4437 21608
rect 4395 21559 4437 21568
rect 4675 21608 4733 21609
rect 4675 21568 4684 21608
rect 4724 21568 4733 21608
rect 4675 21567 4733 21568
rect 4003 21440 4061 21441
rect 4003 21400 4012 21440
rect 4052 21400 4061 21440
rect 4003 21399 4061 21400
rect 576 21188 5952 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 5952 21188
rect 576 21124 5952 21148
rect 74016 21188 99360 21212
rect 74016 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 74016 21124 99360 21148
rect 5155 21020 5213 21021
rect 5155 20980 5164 21020
rect 5204 20980 5213 21020
rect 5155 20979 5213 20980
rect 3139 20768 3197 20769
rect 3139 20728 3148 20768
rect 3188 20728 3197 20768
rect 3139 20727 3197 20728
rect 4003 20768 4061 20769
rect 4003 20728 4012 20768
rect 4052 20728 4061 20768
rect 4003 20727 4061 20728
rect 2763 20684 2805 20693
rect 2763 20644 2764 20684
rect 2804 20644 2805 20684
rect 2763 20635 2805 20644
rect 643 20600 701 20601
rect 643 20560 652 20600
rect 692 20560 701 20600
rect 643 20559 701 20560
rect 576 20432 5952 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 5952 20432
rect 576 20368 5952 20392
rect 74016 20432 99360 20456
rect 74016 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 74016 20368 99360 20392
rect 643 20264 701 20265
rect 643 20224 652 20264
rect 692 20224 701 20264
rect 643 20223 701 20224
rect 2763 20180 2805 20189
rect 2763 20140 2764 20180
rect 2804 20140 2805 20180
rect 2763 20131 2805 20140
rect 81387 20180 81429 20189
rect 81387 20140 81388 20180
rect 81428 20140 81429 20180
rect 81387 20131 81429 20140
rect 2859 20096 2901 20105
rect 2859 20056 2860 20096
rect 2900 20056 2901 20096
rect 2859 20047 2901 20056
rect 3139 20096 3197 20097
rect 3139 20056 3148 20096
rect 3188 20056 3197 20096
rect 3139 20055 3197 20056
rect 3435 20096 3477 20105
rect 3435 20056 3436 20096
rect 3476 20056 3477 20096
rect 3435 20047 3477 20056
rect 3811 20096 3869 20097
rect 3811 20056 3820 20096
rect 3860 20056 3869 20096
rect 3811 20055 3869 20056
rect 4675 20096 4733 20097
rect 4675 20056 4684 20096
rect 4724 20056 4733 20096
rect 4675 20055 4733 20056
rect 80995 20096 81053 20097
rect 80995 20056 81004 20096
rect 81044 20056 81053 20096
rect 80995 20055 81053 20056
rect 81291 20096 81333 20105
rect 81291 20056 81292 20096
rect 81332 20056 81333 20096
rect 81291 20047 81333 20056
rect 81867 20096 81909 20105
rect 81867 20056 81868 20096
rect 81908 20056 81909 20096
rect 81867 20047 81909 20056
rect 82243 20096 82301 20097
rect 82243 20056 82252 20096
rect 82292 20056 82301 20096
rect 82243 20055 82301 20056
rect 83107 20096 83165 20097
rect 83107 20056 83116 20096
rect 83156 20056 83165 20096
rect 83107 20055 83165 20056
rect 5835 20012 5877 20021
rect 5835 19972 5836 20012
rect 5876 19972 5877 20012
rect 5835 19963 5877 19972
rect 84267 20012 84309 20021
rect 84267 19972 84268 20012
rect 84308 19972 84309 20012
rect 84267 19963 84309 19972
rect 2467 19928 2525 19929
rect 2467 19888 2476 19928
rect 2516 19888 2525 19928
rect 2467 19887 2525 19888
rect 81667 19928 81725 19929
rect 81667 19888 81676 19928
rect 81716 19888 81725 19928
rect 81667 19887 81725 19888
rect 576 19676 5952 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 5952 19676
rect 576 19612 5952 19636
rect 74016 19676 99360 19700
rect 74016 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 74016 19612 99360 19636
rect 4291 19508 4349 19509
rect 4291 19468 4300 19508
rect 4340 19468 4349 19508
rect 4291 19467 4349 19468
rect 81483 19508 81525 19517
rect 81483 19468 81484 19508
rect 81524 19468 81525 19508
rect 81483 19459 81525 19468
rect 2083 19340 2141 19341
rect 2083 19300 2092 19340
rect 2132 19300 2141 19340
rect 2083 19299 2141 19300
rect 81283 19340 81341 19341
rect 81283 19300 81292 19340
rect 81332 19300 81341 19340
rect 81283 19299 81341 19300
rect 4587 19256 4629 19265
rect 4587 19216 4588 19256
rect 4628 19216 4629 19256
rect 4587 19207 4629 19216
rect 4683 19256 4725 19265
rect 4683 19216 4684 19256
rect 4724 19216 4725 19256
rect 4683 19207 4725 19216
rect 4963 19256 5021 19257
rect 4963 19216 4972 19256
rect 5012 19216 5021 19256
rect 4963 19215 5021 19216
rect 643 19088 701 19089
rect 643 19048 652 19088
rect 692 19048 701 19088
rect 643 19047 701 19048
rect 1899 19088 1941 19097
rect 1899 19048 1900 19088
rect 1940 19048 1941 19088
rect 1899 19039 1941 19048
rect 81483 19088 81525 19097
rect 81483 19048 81484 19088
rect 81524 19048 81525 19088
rect 81483 19039 81525 19048
rect 576 18920 5952 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 5952 18920
rect 576 18856 5952 18880
rect 74016 18920 81984 18944
rect 74016 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 81984 18920
rect 74016 18856 81984 18880
rect 843 18584 885 18593
rect 843 18544 844 18584
rect 884 18544 885 18584
rect 843 18535 885 18544
rect 1219 18584 1277 18585
rect 1219 18544 1228 18584
rect 1268 18544 1277 18584
rect 1219 18543 1277 18544
rect 2083 18584 2141 18585
rect 2083 18544 2092 18584
rect 2132 18544 2141 18584
rect 2083 18543 2141 18544
rect 3435 18584 3477 18593
rect 3435 18544 3436 18584
rect 3476 18544 3477 18584
rect 3435 18535 3477 18544
rect 3811 18584 3869 18585
rect 3811 18544 3820 18584
rect 3860 18544 3869 18584
rect 3811 18543 3869 18544
rect 4675 18584 4733 18585
rect 4675 18544 4684 18584
rect 4724 18544 4733 18584
rect 4675 18543 4733 18544
rect 3235 18332 3293 18333
rect 3235 18292 3244 18332
rect 3284 18292 3293 18332
rect 3235 18291 3293 18292
rect 5827 18332 5885 18333
rect 5827 18292 5836 18332
rect 5876 18292 5885 18332
rect 5827 18291 5885 18292
rect 576 18164 5952 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 5952 18164
rect 576 18100 5952 18124
rect 74016 18164 81984 18188
rect 74016 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 81984 18164
rect 74016 18100 81984 18124
rect 1603 17996 1661 17997
rect 1603 17956 1612 17996
rect 1652 17956 1661 17996
rect 1603 17955 1661 17956
rect 3907 17996 3965 17997
rect 3907 17956 3916 17996
rect 3956 17956 3965 17996
rect 3907 17955 3965 17956
rect 1411 17828 1469 17829
rect 1411 17788 1420 17828
rect 1460 17788 1469 17828
rect 1411 17787 1469 17788
rect 2659 17828 2717 17829
rect 2659 17788 2668 17828
rect 2708 17788 2717 17828
rect 2659 17787 2717 17788
rect 3235 17828 3293 17829
rect 3235 17788 3244 17828
rect 3284 17788 3293 17828
rect 3235 17787 3293 17788
rect 1899 17744 1941 17753
rect 1899 17704 1900 17744
rect 1940 17704 1941 17744
rect 1899 17695 1941 17704
rect 1995 17744 2037 17753
rect 1995 17704 1996 17744
rect 2036 17704 2037 17744
rect 1995 17695 2037 17704
rect 2275 17744 2333 17745
rect 2275 17704 2284 17744
rect 2324 17704 2333 17744
rect 2275 17703 2333 17704
rect 4299 17744 4341 17753
rect 4299 17704 4300 17744
rect 4340 17704 4341 17744
rect 4299 17695 4341 17704
rect 4579 17744 4637 17745
rect 4579 17704 4588 17744
rect 4628 17704 4637 17744
rect 4579 17703 4637 17704
rect 4203 17660 4245 17669
rect 4203 17620 4204 17660
rect 4244 17620 4245 17660
rect 4203 17611 4245 17620
rect 643 17576 701 17577
rect 643 17536 652 17576
rect 692 17536 701 17576
rect 643 17535 701 17536
rect 1227 17576 1269 17585
rect 1227 17536 1228 17576
rect 1268 17536 1269 17576
rect 1227 17527 1269 17536
rect 2859 17576 2901 17585
rect 2859 17536 2860 17576
rect 2900 17536 2901 17576
rect 2859 17527 2901 17536
rect 3051 17576 3093 17585
rect 3051 17536 3052 17576
rect 3092 17536 3093 17576
rect 3051 17527 3093 17536
rect 576 17408 5952 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 5952 17408
rect 576 17344 5952 17368
rect 74016 17408 81984 17432
rect 74016 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 81984 17408
rect 74016 17344 81984 17368
rect 643 17240 701 17241
rect 643 17200 652 17240
rect 692 17200 701 17240
rect 643 17199 701 17200
rect 1027 17240 1085 17241
rect 1027 17200 1036 17240
rect 1076 17200 1085 17240
rect 1027 17199 1085 17200
rect 1995 17072 2037 17081
rect 1995 17032 1996 17072
rect 2036 17032 2037 17072
rect 1995 17023 2037 17032
rect 2371 17072 2429 17073
rect 2371 17032 2380 17072
rect 2420 17032 2429 17072
rect 2371 17031 2429 17032
rect 3235 17072 3293 17073
rect 3235 17032 3244 17072
rect 3284 17032 3293 17072
rect 3235 17031 3293 17032
rect 74179 17072 74237 17073
rect 74179 17032 74188 17072
rect 74228 17032 74237 17072
rect 74179 17031 74237 17032
rect 75619 16988 75677 16989
rect 75619 16948 75628 16988
rect 75668 16948 75677 16988
rect 75619 16947 75677 16948
rect 4387 16820 4445 16821
rect 4387 16780 4396 16820
rect 4436 16780 4445 16820
rect 4387 16779 4445 16780
rect 576 16652 5952 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 5952 16652
rect 576 16588 5952 16612
rect 74016 16652 81984 16676
rect 74016 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 81984 16652
rect 74016 16588 81984 16612
rect 1603 16484 1661 16485
rect 1603 16444 1612 16484
rect 1652 16444 1661 16484
rect 1603 16443 1661 16444
rect 2571 16484 2613 16493
rect 2571 16444 2572 16484
rect 2612 16444 2613 16484
rect 2571 16435 2613 16444
rect 5827 16484 5885 16485
rect 5827 16444 5836 16484
rect 5876 16444 5885 16484
rect 5827 16443 5885 16444
rect 1219 16316 1277 16317
rect 1219 16276 1228 16316
rect 1268 16276 1277 16316
rect 1219 16275 1277 16276
rect 2755 16316 2813 16317
rect 2755 16276 2764 16316
rect 2804 16276 2813 16316
rect 2755 16275 2813 16276
rect 1899 16232 1941 16241
rect 1899 16192 1900 16232
rect 1940 16192 1941 16232
rect 1899 16183 1941 16192
rect 1995 16232 2037 16241
rect 1995 16192 1996 16232
rect 2036 16192 2037 16232
rect 1995 16183 2037 16192
rect 2275 16232 2333 16233
rect 2275 16192 2284 16232
rect 2324 16192 2333 16232
rect 2275 16191 2333 16192
rect 3811 16232 3869 16233
rect 3811 16192 3820 16232
rect 3860 16192 3869 16232
rect 3811 16191 3869 16192
rect 4675 16232 4733 16233
rect 4675 16192 4684 16232
rect 4724 16192 4733 16232
rect 4675 16191 4733 16192
rect 3435 16148 3477 16157
rect 3435 16108 3436 16148
rect 3476 16108 3477 16148
rect 3435 16099 3477 16108
rect 643 16064 701 16065
rect 643 16024 652 16064
rect 692 16024 701 16064
rect 643 16023 701 16024
rect 1419 16064 1461 16073
rect 1419 16024 1420 16064
rect 1460 16024 1461 16064
rect 1419 16015 1461 16024
rect 2571 16064 2613 16073
rect 2571 16024 2572 16064
rect 2612 16024 2613 16064
rect 2571 16015 2613 16024
rect 576 15896 5952 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 5952 15896
rect 576 15832 5952 15856
rect 74016 15896 81984 15920
rect 74016 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 81984 15896
rect 74016 15832 81984 15856
rect 81859 15728 81917 15729
rect 81859 15688 81868 15728
rect 81908 15688 81917 15728
rect 81859 15687 81917 15688
rect 4491 15644 4533 15653
rect 4491 15604 4492 15644
rect 4532 15604 4533 15644
rect 4491 15595 4533 15604
rect 1419 15560 1461 15569
rect 1419 15520 1420 15560
rect 1460 15520 1461 15560
rect 1419 15511 1461 15520
rect 1515 15560 1557 15569
rect 1515 15520 1516 15560
rect 1556 15520 1557 15560
rect 1515 15511 1557 15520
rect 1611 15560 1653 15569
rect 1611 15520 1612 15560
rect 1652 15520 1653 15560
rect 1611 15511 1653 15520
rect 1987 15560 2045 15561
rect 1987 15520 1996 15560
rect 2036 15520 2045 15560
rect 1987 15519 2045 15520
rect 2187 15560 2229 15569
rect 2187 15520 2188 15560
rect 2228 15520 2229 15560
rect 2187 15511 2229 15520
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 4867 15560 4925 15561
rect 4867 15520 4876 15560
rect 4916 15520 4925 15560
rect 4867 15519 4925 15520
rect 79467 15560 79509 15569
rect 79467 15520 79468 15560
rect 79508 15520 79509 15560
rect 79467 15511 79509 15520
rect 79843 15560 79901 15561
rect 79843 15520 79852 15560
rect 79892 15520 79901 15560
rect 79843 15519 79901 15520
rect 80707 15560 80765 15561
rect 80707 15520 80716 15560
rect 80756 15520 80765 15560
rect 80707 15519 80765 15520
rect 835 15476 893 15477
rect 835 15436 844 15476
rect 884 15436 893 15476
rect 835 15435 893 15436
rect 2091 15476 2133 15485
rect 2091 15436 2092 15476
rect 2132 15436 2133 15476
rect 2091 15427 2133 15436
rect 1795 15392 1853 15393
rect 1795 15352 1804 15392
rect 1844 15352 1853 15392
rect 1795 15351 1853 15352
rect 4195 15392 4253 15393
rect 4195 15352 4204 15392
rect 4244 15352 4253 15392
rect 4195 15351 4253 15352
rect 651 15308 693 15317
rect 651 15268 652 15308
rect 692 15268 693 15308
rect 651 15259 693 15268
rect 576 15140 5952 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 5952 15140
rect 576 15076 5952 15100
rect 74016 15140 81984 15164
rect 74016 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 81984 15140
rect 74016 15076 81984 15100
rect 3235 14972 3293 14973
rect 3235 14932 3244 14972
rect 3284 14932 3293 14972
rect 3235 14931 3293 14932
rect 80419 14972 80477 14973
rect 80419 14932 80428 14972
rect 80468 14932 80477 14972
rect 80419 14931 80477 14932
rect 1219 14720 1277 14721
rect 1219 14680 1228 14720
rect 1268 14680 1277 14720
rect 1219 14679 1277 14680
rect 2083 14720 2141 14721
rect 2083 14680 2092 14720
rect 2132 14680 2141 14720
rect 2083 14679 2141 14680
rect 3811 14720 3869 14721
rect 3811 14680 3820 14720
rect 3860 14680 3869 14720
rect 3811 14679 3869 14680
rect 4675 14720 4733 14721
rect 4675 14680 4684 14720
rect 4724 14680 4733 14720
rect 4675 14679 4733 14680
rect 80715 14720 80757 14729
rect 80715 14680 80716 14720
rect 80756 14680 80757 14720
rect 80715 14671 80757 14680
rect 80811 14720 80853 14729
rect 80811 14680 80812 14720
rect 80852 14680 80853 14720
rect 80811 14671 80853 14680
rect 81091 14720 81149 14721
rect 81091 14680 81100 14720
rect 81140 14680 81149 14720
rect 81091 14679 81149 14680
rect 843 14636 885 14645
rect 843 14596 844 14636
rect 884 14596 885 14636
rect 843 14587 885 14596
rect 3435 14636 3477 14645
rect 3435 14596 3436 14636
rect 3476 14596 3477 14636
rect 3435 14587 3477 14596
rect 5827 14552 5885 14553
rect 5827 14512 5836 14552
rect 5876 14512 5885 14552
rect 5827 14511 5885 14512
rect 576 14384 5952 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 5952 14384
rect 576 14320 5952 14344
rect 74016 14384 81984 14408
rect 74016 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 81984 14384
rect 74016 14320 81984 14344
rect 1611 14132 1653 14141
rect 1611 14092 1612 14132
rect 1652 14092 1653 14132
rect 1611 14083 1653 14092
rect 3915 14132 3957 14141
rect 3915 14092 3916 14132
rect 3956 14092 3957 14132
rect 3915 14083 3957 14092
rect 1707 14048 1749 14057
rect 1707 14008 1708 14048
rect 1748 14008 1749 14048
rect 1707 13999 1749 14008
rect 1987 14048 2045 14049
rect 1987 14008 1996 14048
rect 2036 14008 2045 14048
rect 1987 14007 2045 14008
rect 4011 14048 4053 14057
rect 4011 14008 4012 14048
rect 4052 14008 4053 14048
rect 4011 13999 4053 14008
rect 4291 14048 4349 14049
rect 4291 14008 4300 14048
rect 4340 14008 4349 14048
rect 4291 14007 4349 14008
rect 835 13964 893 13965
rect 835 13924 844 13964
rect 884 13924 893 13964
rect 835 13923 893 13924
rect 76387 13964 76445 13965
rect 76387 13924 76396 13964
rect 76436 13924 76445 13964
rect 76387 13923 76445 13924
rect 651 13880 693 13889
rect 651 13840 652 13880
rect 692 13840 693 13880
rect 651 13831 693 13840
rect 1315 13880 1373 13881
rect 1315 13840 1324 13880
rect 1364 13840 1373 13880
rect 1315 13839 1373 13840
rect 3619 13880 3677 13881
rect 3619 13840 3628 13880
rect 3668 13840 3677 13880
rect 3619 13839 3677 13840
rect 76203 13796 76245 13805
rect 76203 13756 76204 13796
rect 76244 13756 76245 13796
rect 76203 13747 76245 13756
rect 576 13628 5952 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 5952 13628
rect 576 13564 5952 13588
rect 74016 13628 81984 13652
rect 74016 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 81984 13628
rect 74016 13564 81984 13588
rect 1899 13460 1941 13469
rect 1899 13420 1900 13460
rect 1940 13420 1941 13460
rect 1899 13411 1941 13420
rect 5827 13460 5885 13461
rect 5827 13420 5836 13460
rect 5876 13420 5885 13460
rect 5827 13419 5885 13420
rect 81859 13460 81917 13461
rect 81859 13420 81868 13460
rect 81908 13420 81917 13460
rect 81859 13419 81917 13420
rect 76579 13376 76637 13377
rect 76579 13336 76588 13376
rect 76628 13336 76637 13376
rect 76579 13335 76637 13336
rect 835 13292 893 13293
rect 835 13252 844 13292
rect 884 13252 893 13292
rect 835 13251 893 13252
rect 1515 13208 1557 13217
rect 1515 13168 1516 13208
rect 1556 13168 1557 13208
rect 1515 13159 1557 13168
rect 1707 13208 1749 13217
rect 1707 13168 1708 13208
rect 1748 13168 1749 13208
rect 3811 13208 3869 13209
rect 1707 13159 1749 13168
rect 1987 13197 2045 13198
rect 1987 13157 1996 13197
rect 2036 13157 2045 13197
rect 3811 13168 3820 13208
rect 3860 13168 3869 13208
rect 3811 13167 3869 13168
rect 4675 13208 4733 13209
rect 4675 13168 4684 13208
rect 4724 13168 4733 13208
rect 4675 13167 4733 13168
rect 75907 13208 75965 13209
rect 75907 13168 75916 13208
rect 75956 13168 75965 13208
rect 75907 13167 75965 13168
rect 76203 13208 76245 13217
rect 76203 13168 76204 13208
rect 76244 13168 76245 13208
rect 76203 13159 76245 13168
rect 76779 13208 76821 13217
rect 76779 13168 76780 13208
rect 76820 13168 76821 13208
rect 76779 13159 76821 13168
rect 77155 13208 77213 13209
rect 77155 13168 77164 13208
rect 77204 13168 77213 13208
rect 77155 13167 77213 13168
rect 78019 13208 78077 13209
rect 78019 13168 78028 13208
rect 78068 13168 78077 13208
rect 78019 13167 78077 13168
rect 79843 13208 79901 13209
rect 79843 13168 79852 13208
rect 79892 13168 79901 13208
rect 79843 13167 79901 13168
rect 80707 13208 80765 13209
rect 80707 13168 80716 13208
rect 80756 13168 80765 13208
rect 80707 13167 80765 13168
rect 1987 13156 2045 13157
rect 3435 13124 3477 13133
rect 3435 13084 3436 13124
rect 3476 13084 3477 13124
rect 3435 13075 3477 13084
rect 76299 13124 76341 13133
rect 76299 13084 76300 13124
rect 76340 13084 76341 13124
rect 76299 13075 76341 13084
rect 79467 13124 79509 13133
rect 79467 13084 79468 13124
rect 79508 13084 79509 13124
rect 79467 13075 79509 13084
rect 651 13040 693 13049
rect 651 13000 652 13040
rect 692 13000 693 13040
rect 651 12991 693 13000
rect 1611 13040 1653 13049
rect 1611 13000 1612 13040
rect 1652 13000 1653 13040
rect 1611 12991 1653 13000
rect 75627 13040 75669 13049
rect 75627 13000 75628 13040
rect 75668 13000 75669 13040
rect 75627 12991 75669 13000
rect 79171 13040 79229 13041
rect 79171 13000 79180 13040
rect 79220 13000 79229 13040
rect 79171 12999 79229 13000
rect 81859 13040 81917 13041
rect 81859 13000 81868 13040
rect 81908 13000 81917 13040
rect 81859 12999 81917 13000
rect 576 12872 5952 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 5952 12872
rect 576 12808 5952 12832
rect 74016 12872 81984 12896
rect 74016 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 81984 12872
rect 74016 12808 81984 12832
rect 77259 12704 77301 12713
rect 77259 12664 77260 12704
rect 77300 12664 77301 12704
rect 77259 12655 77301 12664
rect 4203 12620 4245 12629
rect 4203 12580 4204 12620
rect 4244 12580 4245 12620
rect 4203 12571 4245 12580
rect 80235 12620 80277 12629
rect 80235 12580 80236 12620
rect 80276 12580 80277 12620
rect 80235 12571 80277 12580
rect 843 12536 885 12545
rect 843 12496 844 12536
rect 884 12496 885 12536
rect 843 12487 885 12496
rect 1131 12536 1173 12545
rect 1131 12496 1132 12536
rect 1172 12496 1173 12536
rect 1131 12487 1173 12496
rect 1323 12536 1365 12545
rect 1323 12496 1324 12536
rect 1364 12496 1365 12536
rect 1323 12487 1365 12496
rect 1699 12536 1757 12537
rect 1699 12496 1708 12536
rect 1748 12496 1757 12536
rect 1699 12495 1757 12496
rect 2563 12536 2621 12537
rect 2563 12496 2572 12536
rect 2612 12496 2621 12536
rect 2563 12495 2621 12496
rect 4299 12536 4341 12545
rect 4299 12496 4300 12536
rect 4340 12496 4341 12536
rect 4299 12487 4341 12496
rect 4579 12536 4637 12537
rect 4579 12496 4588 12536
rect 4628 12496 4637 12536
rect 4579 12495 4637 12496
rect 79075 12536 79133 12537
rect 79075 12496 79084 12536
rect 79124 12496 79133 12536
rect 79075 12495 79133 12496
rect 79371 12536 79413 12545
rect 79371 12496 79372 12536
rect 79412 12496 79413 12536
rect 79371 12487 79413 12496
rect 79467 12536 79509 12545
rect 79467 12496 79468 12536
rect 79508 12496 79509 12536
rect 79467 12487 79509 12496
rect 80331 12536 80373 12545
rect 80331 12496 80332 12536
rect 80372 12496 80373 12536
rect 80331 12487 80373 12496
rect 80611 12536 80669 12537
rect 80611 12496 80620 12536
rect 80660 12496 80669 12536
rect 80611 12495 80669 12496
rect 939 12452 981 12461
rect 939 12412 940 12452
rect 980 12412 981 12452
rect 939 12403 981 12412
rect 77443 12452 77501 12453
rect 77443 12412 77452 12452
rect 77492 12412 77501 12452
rect 77443 12411 77501 12412
rect 3907 12368 3965 12369
rect 3907 12328 3916 12368
rect 3956 12328 3965 12368
rect 3907 12327 3965 12328
rect 79939 12368 79997 12369
rect 79939 12328 79948 12368
rect 79988 12328 79997 12368
rect 79939 12327 79997 12328
rect 3715 12284 3773 12285
rect 3715 12244 3724 12284
rect 3764 12244 3773 12284
rect 3715 12243 3773 12244
rect 79747 12284 79805 12285
rect 79747 12244 79756 12284
rect 79796 12244 79805 12284
rect 79747 12243 79805 12244
rect 576 12116 5952 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 5952 12116
rect 576 12052 5952 12076
rect 74016 12116 81984 12140
rect 74016 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 81984 12116
rect 74016 12052 81984 12076
rect 651 11948 693 11957
rect 651 11908 652 11948
rect 692 11908 693 11948
rect 651 11899 693 11908
rect 1315 11948 1373 11949
rect 1315 11908 1324 11948
rect 1364 11908 1373 11948
rect 1315 11907 1373 11908
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 5835 11780 5877 11789
rect 5835 11740 5836 11780
rect 5876 11740 5877 11780
rect 5835 11731 5877 11740
rect 81867 11780 81909 11789
rect 81867 11740 81868 11780
rect 81908 11740 81909 11780
rect 81867 11731 81909 11740
rect 1611 11696 1653 11705
rect 1611 11656 1612 11696
rect 1652 11656 1653 11696
rect 1611 11647 1653 11656
rect 1707 11696 1749 11705
rect 1707 11656 1708 11696
rect 1748 11656 1749 11696
rect 1707 11647 1749 11656
rect 1987 11696 2045 11697
rect 1987 11656 1996 11696
rect 2036 11656 2045 11696
rect 1987 11655 2045 11656
rect 3811 11696 3869 11697
rect 3811 11656 3820 11696
rect 3860 11656 3869 11696
rect 3811 11655 3869 11656
rect 4675 11696 4733 11697
rect 4675 11656 4684 11696
rect 4724 11656 4733 11696
rect 4675 11655 4733 11656
rect 79467 11696 79509 11705
rect 79467 11656 79468 11696
rect 79508 11656 79509 11696
rect 79467 11647 79509 11656
rect 79843 11696 79901 11697
rect 79843 11656 79852 11696
rect 79892 11656 79901 11696
rect 79843 11655 79901 11656
rect 80707 11696 80765 11697
rect 80707 11656 80716 11696
rect 80756 11656 80765 11696
rect 80707 11655 80765 11656
rect 3435 11612 3477 11621
rect 3435 11572 3436 11612
rect 3476 11572 3477 11612
rect 3435 11563 3477 11572
rect 576 11360 5952 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 5952 11360
rect 576 11296 5952 11320
rect 74016 11360 81984 11384
rect 74016 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 81984 11360
rect 74016 11296 81984 11320
rect 651 11192 693 11201
rect 651 11152 652 11192
rect 692 11152 693 11192
rect 651 11143 693 11152
rect 1699 11192 1757 11193
rect 1699 11152 1708 11192
rect 1748 11152 1757 11192
rect 1699 11151 1757 11152
rect 1411 11108 1469 11109
rect 1411 11068 1420 11108
rect 1460 11068 1469 11108
rect 1411 11067 1469 11068
rect 4011 11108 4053 11117
rect 4011 11068 4012 11108
rect 4052 11068 4053 11108
rect 4011 11059 4053 11068
rect 1603 11024 1661 11025
rect 1603 10984 1612 11024
rect 1652 10984 1661 11024
rect 1603 10983 1661 10984
rect 4107 11024 4149 11033
rect 4107 10984 4108 11024
rect 4148 10984 4149 11024
rect 4107 10975 4149 10984
rect 4387 11024 4445 11025
rect 4387 10984 4396 11024
rect 4436 10984 4445 11024
rect 4387 10983 4445 10984
rect 80139 11024 80181 11033
rect 80139 10984 80140 11024
rect 80180 10984 80181 11024
rect 80139 10975 80181 10984
rect 80235 11024 80277 11033
rect 80235 10984 80236 11024
rect 80276 10984 80277 11024
rect 80235 10975 80277 10984
rect 80515 11024 80573 11025
rect 80515 10984 80524 11024
rect 80564 10984 80573 11024
rect 80515 10983 80573 10984
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 1219 10940 1277 10941
rect 1219 10900 1228 10940
rect 1268 10900 1277 10940
rect 1219 10899 1277 10900
rect 3715 10856 3773 10857
rect 3715 10816 3724 10856
rect 3764 10816 3773 10856
rect 3715 10815 3773 10816
rect 1035 10772 1077 10781
rect 1035 10732 1036 10772
rect 1076 10732 1077 10772
rect 1035 10723 1077 10732
rect 79843 10772 79901 10773
rect 79843 10732 79852 10772
rect 79892 10732 79901 10772
rect 79843 10731 79901 10732
rect 576 10604 5952 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 5952 10604
rect 576 10540 5952 10564
rect 74016 10604 81984 10628
rect 74016 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 81984 10604
rect 74016 10540 81984 10564
rect 5827 10436 5885 10437
rect 5827 10396 5836 10436
rect 5876 10396 5885 10436
rect 5827 10395 5885 10396
rect 3243 10268 3285 10277
rect 3243 10228 3244 10268
rect 3284 10228 3285 10268
rect 3243 10219 3285 10228
rect 81867 10268 81909 10277
rect 81867 10228 81868 10268
rect 81908 10228 81909 10268
rect 81867 10219 81909 10228
rect 1219 10184 1277 10185
rect 1219 10144 1228 10184
rect 1268 10144 1277 10184
rect 1219 10143 1277 10144
rect 2083 10184 2141 10185
rect 2083 10144 2092 10184
rect 2132 10144 2141 10184
rect 2083 10143 2141 10144
rect 3811 10184 3869 10185
rect 3811 10144 3820 10184
rect 3860 10144 3869 10184
rect 3811 10143 3869 10144
rect 4675 10184 4733 10185
rect 4675 10144 4684 10184
rect 4724 10144 4733 10184
rect 4675 10143 4733 10144
rect 79467 10184 79509 10193
rect 79467 10144 79468 10184
rect 79508 10144 79509 10184
rect 79467 10135 79509 10144
rect 79843 10184 79901 10185
rect 79843 10144 79852 10184
rect 79892 10144 79901 10184
rect 79843 10143 79901 10144
rect 80707 10184 80765 10185
rect 80707 10144 80716 10184
rect 80756 10144 80765 10184
rect 80707 10143 80765 10144
rect 843 10100 885 10109
rect 843 10060 844 10100
rect 884 10060 885 10100
rect 843 10051 885 10060
rect 3435 10100 3477 10109
rect 3435 10060 3436 10100
rect 3476 10060 3477 10100
rect 3435 10051 3477 10060
rect 576 9848 5952 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 5952 9848
rect 576 9784 5952 9808
rect 74016 9848 81984 9872
rect 74016 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 81984 9848
rect 74016 9784 81984 9808
rect 651 9680 693 9689
rect 651 9640 652 9680
rect 692 9640 693 9680
rect 651 9631 693 9640
rect 1027 9680 1085 9681
rect 1027 9640 1036 9680
rect 1076 9640 1085 9680
rect 1027 9639 1085 9640
rect 1315 9680 1373 9681
rect 1315 9640 1324 9680
rect 1364 9640 1373 9680
rect 1315 9639 1373 9640
rect 1803 9596 1845 9605
rect 1803 9556 1804 9596
rect 1844 9556 1845 9596
rect 1803 9547 1845 9556
rect 4299 9596 4341 9605
rect 4299 9556 4300 9596
rect 4340 9556 4341 9596
rect 4299 9547 4341 9556
rect 1219 9512 1277 9513
rect 1219 9472 1228 9512
rect 1268 9472 1277 9512
rect 1219 9471 1277 9472
rect 1899 9512 1941 9521
rect 1899 9472 1900 9512
rect 1940 9472 1941 9512
rect 1899 9463 1941 9472
rect 2179 9512 2237 9513
rect 2179 9472 2188 9512
rect 2228 9472 2237 9512
rect 2179 9471 2237 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4675 9512 4733 9513
rect 4675 9472 4684 9512
rect 4724 9472 4733 9512
rect 4675 9471 4733 9472
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 1507 9344 1565 9345
rect 1507 9304 1516 9344
rect 1556 9304 1565 9344
rect 1507 9303 1565 9304
rect 4003 9344 4061 9345
rect 4003 9304 4012 9344
rect 4052 9304 4061 9344
rect 4003 9303 4061 9304
rect 576 9092 5952 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 5952 9092
rect 576 9028 5952 9052
rect 74016 9092 81984 9116
rect 74016 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 81984 9092
rect 74016 9028 81984 9052
rect 651 8924 693 8933
rect 651 8884 652 8924
rect 692 8884 693 8924
rect 651 8875 693 8884
rect 5251 8924 5309 8925
rect 5251 8884 5260 8924
rect 5300 8884 5309 8924
rect 5251 8883 5309 8884
rect 1411 8840 1469 8841
rect 1411 8800 1420 8840
rect 1460 8800 1469 8840
rect 1411 8799 1469 8800
rect 2659 8840 2717 8841
rect 2659 8800 2668 8840
rect 2708 8800 2717 8840
rect 2659 8799 2717 8800
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 1603 8672 1661 8673
rect 1603 8632 1612 8672
rect 1652 8632 1661 8672
rect 1603 8631 1661 8632
rect 1987 8672 2045 8673
rect 1987 8632 1996 8672
rect 2036 8632 2045 8672
rect 1987 8631 2045 8632
rect 2283 8672 2325 8681
rect 2283 8632 2284 8672
rect 2324 8632 2325 8672
rect 2283 8623 2325 8632
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 2859 8672 2901 8681
rect 2859 8632 2860 8672
rect 2900 8632 2901 8672
rect 2859 8623 2901 8632
rect 3235 8672 3293 8673
rect 3235 8632 3244 8672
rect 3284 8632 3293 8672
rect 3235 8631 3293 8632
rect 4099 8672 4157 8673
rect 4099 8632 4108 8672
rect 4148 8632 4157 8672
rect 4099 8631 4157 8632
rect 1027 8504 1085 8505
rect 1027 8464 1036 8504
rect 1076 8464 1085 8504
rect 1027 8463 1085 8464
rect 1699 8504 1757 8505
rect 1699 8464 1708 8504
rect 1748 8464 1757 8504
rect 1699 8463 1757 8464
rect 576 8336 5952 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 5952 8336
rect 576 8272 5952 8296
rect 74016 8336 81984 8360
rect 74016 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 81984 8336
rect 74016 8272 81984 8296
rect 643 8168 701 8169
rect 643 8128 652 8168
rect 692 8128 701 8168
rect 643 8127 701 8128
rect 3435 8000 3477 8009
rect 3435 7960 3436 8000
rect 3476 7960 3477 8000
rect 3435 7951 3477 7960
rect 3811 8000 3869 8001
rect 3811 7960 3820 8000
rect 3860 7960 3869 8000
rect 3811 7959 3869 7960
rect 4675 8000 4733 8001
rect 4675 7960 4684 8000
rect 4724 7960 4733 8000
rect 4675 7959 4733 7960
rect 5827 7748 5885 7749
rect 5827 7708 5836 7748
rect 5876 7708 5885 7748
rect 5827 7707 5885 7708
rect 576 7580 5952 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 5952 7580
rect 576 7516 5952 7540
rect 74016 7580 81984 7604
rect 74016 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 81984 7580
rect 74016 7516 81984 7540
rect 3523 7412 3581 7413
rect 3523 7372 3532 7412
rect 3572 7372 3581 7412
rect 3523 7371 3581 7372
rect 1323 7160 1365 7169
rect 1323 7120 1324 7160
rect 1364 7120 1365 7160
rect 1323 7111 1365 7120
rect 1411 7160 1469 7161
rect 1411 7120 1420 7160
rect 1460 7120 1469 7160
rect 1411 7119 1469 7120
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 1699 7160 1757 7161
rect 1699 7120 1708 7160
rect 1748 7120 1757 7160
rect 1699 7119 1757 7120
rect 1987 7160 2045 7161
rect 1987 7120 1996 7160
rect 2036 7120 2045 7160
rect 1987 7119 2045 7120
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 3915 7160 3957 7169
rect 3915 7120 3916 7160
rect 3956 7120 3957 7160
rect 3915 7111 3957 7120
rect 4195 7160 4253 7161
rect 4195 7120 4204 7160
rect 4244 7120 4253 7160
rect 4195 7119 4253 7120
rect 1899 7076 1941 7085
rect 1899 7036 1900 7076
rect 1940 7036 1941 7076
rect 1899 7027 1941 7036
rect 643 6992 701 6993
rect 643 6952 652 6992
rect 692 6952 701 6992
rect 643 6951 701 6952
rect 576 6824 5952 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 5952 6824
rect 576 6760 5952 6784
rect 74016 6824 81984 6848
rect 74016 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 81984 6824
rect 74016 6760 81984 6784
rect 81859 6656 81917 6657
rect 81859 6616 81868 6656
rect 81908 6616 81917 6656
rect 81859 6615 81917 6616
rect 79467 6488 79509 6497
rect 79467 6448 79468 6488
rect 79508 6448 79509 6488
rect 79467 6439 79509 6448
rect 79843 6488 79901 6489
rect 79843 6448 79852 6488
rect 79892 6448 79901 6488
rect 79843 6447 79901 6448
rect 80707 6488 80765 6489
rect 80707 6448 80716 6488
rect 80756 6448 80765 6488
rect 80707 6447 80765 6448
rect 81859 6236 81917 6237
rect 81859 6196 81868 6236
rect 81908 6196 81917 6236
rect 81859 6195 81917 6196
rect 576 6068 5952 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 5952 6068
rect 576 6004 5952 6028
rect 74016 6068 81984 6092
rect 74016 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 81984 6068
rect 74016 6004 81984 6028
rect 80131 5900 80189 5901
rect 80131 5860 80140 5900
rect 80180 5860 80189 5900
rect 80131 5859 80189 5860
rect 5835 5732 5877 5741
rect 5835 5692 5836 5732
rect 5876 5692 5877 5732
rect 5835 5683 5877 5692
rect 3811 5648 3869 5649
rect 3811 5608 3820 5648
rect 3860 5608 3869 5648
rect 3811 5607 3869 5608
rect 4675 5648 4733 5649
rect 4675 5608 4684 5648
rect 4724 5608 4733 5648
rect 4675 5607 4733 5608
rect 80427 5648 80469 5657
rect 80427 5608 80428 5648
rect 80468 5608 80469 5648
rect 80427 5599 80469 5608
rect 80523 5648 80565 5657
rect 80523 5608 80524 5648
rect 80564 5608 80565 5648
rect 80523 5599 80565 5608
rect 80803 5648 80861 5649
rect 80803 5608 80812 5648
rect 80852 5608 80861 5648
rect 80803 5607 80861 5608
rect 3435 5564 3477 5573
rect 3435 5524 3436 5564
rect 3476 5524 3477 5564
rect 3435 5515 3477 5524
rect 643 5480 701 5481
rect 643 5440 652 5480
rect 692 5440 701 5480
rect 643 5439 701 5440
rect 576 5312 5952 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 5952 5312
rect 576 5248 5952 5272
rect 74016 5312 81984 5336
rect 74016 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 81984 5312
rect 74016 5248 81984 5272
rect 643 5144 701 5145
rect 643 5104 652 5144
rect 692 5104 701 5144
rect 643 5103 701 5104
rect 4491 5060 4533 5069
rect 4491 5020 4492 5060
rect 4532 5020 4533 5060
rect 4491 5011 4533 5020
rect 4587 4976 4629 4985
rect 4587 4936 4588 4976
rect 4628 4936 4629 4976
rect 4587 4927 4629 4936
rect 4867 4976 4925 4977
rect 4867 4936 4876 4976
rect 4916 4936 4925 4976
rect 4867 4935 4925 4936
rect 80139 4976 80181 4985
rect 80139 4936 80140 4976
rect 80180 4936 80181 4976
rect 80139 4927 80181 4936
rect 80235 4976 80277 4985
rect 80235 4936 80236 4976
rect 80276 4936 80277 4976
rect 80235 4927 80277 4936
rect 80515 4976 80573 4977
rect 80515 4936 80524 4976
rect 80564 4936 80573 4976
rect 80515 4935 80573 4936
rect 4195 4808 4253 4809
rect 4195 4768 4204 4808
rect 4244 4768 4253 4808
rect 4195 4767 4253 4768
rect 79843 4724 79901 4725
rect 79843 4684 79852 4724
rect 79892 4684 79901 4724
rect 79843 4683 79901 4684
rect 576 4556 5952 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 5952 4556
rect 576 4492 5952 4516
rect 74016 4556 81984 4580
rect 74016 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 81984 4556
rect 74016 4492 81984 4516
rect 81859 4388 81917 4389
rect 81859 4348 81868 4388
rect 81908 4348 81917 4388
rect 81859 4347 81917 4348
rect 79467 4136 79509 4145
rect 79467 4096 79468 4136
rect 79508 4096 79509 4136
rect 79467 4087 79509 4096
rect 79843 4136 79901 4137
rect 79843 4096 79852 4136
rect 79892 4096 79901 4136
rect 79843 4095 79901 4096
rect 80707 4136 80765 4137
rect 80707 4096 80716 4136
rect 80756 4096 80765 4136
rect 80707 4095 80765 4096
rect 643 3968 701 3969
rect 643 3928 652 3968
rect 692 3928 701 3968
rect 643 3927 701 3928
rect 81859 3968 81917 3969
rect 81859 3928 81868 3968
rect 81908 3928 81917 3968
rect 81859 3927 81917 3928
rect 576 3800 81984 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 81984 3800
rect 576 3736 81984 3760
rect 643 3632 701 3633
rect 643 3592 652 3632
rect 692 3592 701 3632
rect 643 3591 701 3592
rect 16195 3632 16253 3633
rect 16195 3592 16204 3632
rect 16244 3592 16253 3632
rect 16195 3591 16253 3592
rect 19267 3632 19325 3633
rect 19267 3592 19276 3632
rect 19316 3592 19325 3632
rect 19267 3591 19325 3592
rect 25027 3632 25085 3633
rect 25027 3592 25036 3632
rect 25076 3592 25085 3632
rect 25027 3591 25085 3592
rect 13323 3548 13365 3557
rect 13323 3508 13324 3548
rect 13364 3508 13365 3548
rect 13323 3499 13365 3508
rect 20331 3548 20373 3557
rect 20331 3508 20332 3548
rect 20372 3508 20373 3548
rect 20331 3499 20373 3508
rect 22155 3548 22197 3557
rect 22155 3508 22156 3548
rect 22196 3508 22197 3548
rect 22155 3499 22197 3508
rect 28779 3548 28821 3557
rect 28779 3508 28780 3548
rect 28820 3508 28821 3548
rect 28779 3499 28821 3508
rect 33291 3548 33333 3557
rect 33291 3508 33292 3548
rect 33332 3508 33333 3548
rect 33291 3499 33333 3508
rect 46443 3548 46485 3557
rect 46443 3508 46444 3548
rect 46484 3508 46485 3548
rect 46443 3499 46485 3508
rect 49035 3548 49077 3557
rect 49035 3508 49036 3548
rect 49076 3508 49077 3548
rect 49035 3499 49077 3508
rect 52203 3548 52245 3557
rect 52203 3508 52204 3548
rect 52244 3508 52245 3548
rect 52203 3499 52245 3508
rect 54987 3548 55029 3557
rect 54987 3508 54988 3548
rect 55028 3508 55029 3548
rect 54987 3499 55029 3508
rect 17251 3477 17309 3478
rect 12931 3464 12989 3465
rect 12931 3424 12940 3464
rect 12980 3424 12989 3464
rect 12931 3423 12989 3424
rect 13227 3464 13269 3473
rect 13227 3424 13228 3464
rect 13268 3424 13269 3464
rect 13227 3415 13269 3424
rect 13803 3464 13845 3473
rect 13803 3424 13804 3464
rect 13844 3424 13845 3464
rect 13803 3415 13845 3424
rect 14179 3464 14237 3465
rect 14179 3424 14188 3464
rect 14228 3424 14237 3464
rect 14179 3423 14237 3424
rect 15043 3464 15101 3465
rect 15043 3424 15052 3464
rect 15092 3424 15101 3464
rect 15043 3423 15101 3424
rect 16875 3464 16917 3473
rect 16875 3424 16876 3464
rect 16916 3424 16917 3464
rect 17251 3437 17260 3477
rect 17300 3437 17309 3477
rect 17251 3436 17309 3437
rect 18115 3464 18173 3465
rect 16875 3415 16917 3424
rect 18115 3424 18124 3464
rect 18164 3424 18173 3464
rect 18115 3423 18173 3424
rect 20427 3464 20469 3473
rect 20427 3424 20428 3464
rect 20468 3424 20469 3464
rect 20427 3415 20469 3424
rect 20707 3464 20765 3465
rect 20707 3424 20716 3464
rect 20756 3424 20765 3464
rect 20707 3423 20765 3424
rect 21763 3464 21821 3465
rect 21763 3424 21772 3464
rect 21812 3424 21821 3464
rect 21763 3423 21821 3424
rect 22059 3464 22101 3473
rect 22059 3424 22060 3464
rect 22100 3424 22101 3464
rect 22059 3415 22101 3424
rect 22635 3464 22677 3473
rect 22635 3424 22636 3464
rect 22676 3424 22677 3464
rect 22635 3415 22677 3424
rect 23011 3464 23069 3465
rect 23011 3424 23020 3464
rect 23060 3424 23069 3464
rect 23011 3423 23069 3424
rect 23875 3464 23933 3465
rect 23875 3424 23884 3464
rect 23924 3424 23933 3464
rect 23875 3423 23933 3424
rect 28387 3464 28445 3465
rect 28387 3424 28396 3464
rect 28436 3424 28445 3464
rect 28387 3423 28445 3424
rect 28683 3464 28725 3473
rect 28683 3424 28684 3464
rect 28724 3424 28725 3464
rect 28683 3415 28725 3424
rect 30787 3464 30845 3465
rect 30787 3424 30796 3464
rect 30836 3424 30845 3464
rect 30787 3423 30845 3424
rect 31179 3464 31221 3473
rect 31179 3424 31180 3464
rect 31220 3424 31221 3464
rect 31179 3415 31221 3424
rect 33387 3464 33429 3473
rect 33387 3424 33388 3464
rect 33428 3424 33429 3464
rect 33387 3415 33429 3424
rect 33667 3464 33725 3465
rect 33667 3424 33676 3464
rect 33716 3424 33725 3464
rect 33667 3423 33725 3424
rect 33955 3464 34013 3465
rect 33955 3424 33964 3464
rect 34004 3424 34013 3464
rect 33955 3423 34013 3424
rect 34347 3464 34389 3473
rect 34347 3424 34348 3464
rect 34388 3424 34389 3464
rect 34347 3415 34389 3424
rect 34627 3464 34685 3465
rect 34627 3424 34636 3464
rect 34676 3424 34685 3464
rect 34627 3423 34685 3424
rect 34923 3464 34965 3473
rect 34923 3424 34924 3464
rect 34964 3424 34965 3464
rect 34923 3415 34965 3424
rect 35019 3464 35061 3473
rect 35019 3424 35020 3464
rect 35060 3424 35061 3464
rect 35019 3415 35061 3424
rect 36643 3464 36701 3465
rect 36643 3424 36652 3464
rect 36692 3424 36701 3464
rect 36643 3423 36701 3424
rect 37035 3464 37077 3473
rect 37035 3424 37036 3464
rect 37076 3424 37077 3464
rect 37035 3415 37077 3424
rect 37219 3464 37277 3465
rect 37219 3424 37228 3464
rect 37268 3424 37277 3464
rect 37219 3423 37277 3424
rect 37611 3464 37653 3473
rect 37611 3424 37612 3464
rect 37652 3424 37653 3464
rect 37611 3415 37653 3424
rect 37803 3464 37845 3473
rect 37803 3424 37804 3464
rect 37844 3424 37845 3464
rect 37803 3415 37845 3424
rect 38179 3464 38237 3465
rect 38179 3424 38188 3464
rect 38228 3424 38237 3464
rect 38179 3423 38237 3424
rect 39243 3464 39285 3473
rect 39243 3424 39244 3464
rect 39284 3424 39285 3464
rect 39243 3415 39285 3424
rect 39339 3464 39381 3473
rect 39339 3424 39340 3464
rect 39380 3424 39381 3464
rect 39339 3415 39381 3424
rect 39619 3464 39677 3465
rect 39619 3424 39628 3464
rect 39668 3424 39677 3464
rect 39619 3423 39677 3424
rect 42691 3464 42749 3465
rect 42691 3424 42700 3464
rect 42740 3424 42749 3464
rect 42691 3423 42749 3424
rect 46051 3464 46109 3465
rect 46051 3424 46060 3464
rect 46100 3424 46109 3464
rect 46051 3423 46109 3424
rect 46347 3464 46389 3473
rect 46347 3424 46348 3464
rect 46388 3424 46389 3464
rect 46347 3415 46389 3424
rect 48643 3464 48701 3465
rect 48643 3424 48652 3464
rect 48692 3424 48701 3464
rect 48643 3423 48701 3424
rect 48939 3464 48981 3473
rect 48939 3424 48940 3464
rect 48980 3424 48981 3464
rect 48939 3415 48981 3424
rect 51811 3464 51869 3465
rect 51811 3424 51820 3464
rect 51860 3424 51869 3464
rect 51811 3423 51869 3424
rect 52107 3464 52149 3473
rect 52107 3424 52108 3464
rect 52148 3424 52149 3464
rect 52107 3415 52149 3424
rect 54595 3464 54653 3465
rect 54595 3424 54604 3464
rect 54644 3424 54653 3464
rect 54595 3423 54653 3424
rect 54891 3464 54933 3473
rect 54891 3424 54892 3464
rect 54932 3424 54933 3464
rect 54891 3415 54933 3424
rect 21283 3380 21341 3381
rect 21283 3340 21292 3380
rect 21332 3340 21341 3380
rect 21283 3339 21341 3340
rect 30891 3380 30933 3389
rect 30891 3340 30892 3380
rect 30932 3340 30933 3380
rect 30891 3331 30933 3340
rect 31083 3380 31125 3389
rect 31083 3340 31084 3380
rect 31124 3340 31125 3380
rect 31083 3331 31125 3340
rect 32803 3380 32861 3381
rect 32803 3340 32812 3380
rect 32852 3340 32861 3380
rect 32803 3339 32861 3340
rect 34059 3380 34101 3389
rect 34059 3340 34060 3380
rect 34100 3340 34101 3380
rect 34059 3331 34101 3340
rect 34251 3380 34293 3389
rect 34251 3340 34252 3380
rect 34292 3340 34293 3380
rect 34251 3331 34293 3340
rect 36747 3380 36789 3389
rect 36747 3340 36748 3380
rect 36788 3340 36789 3380
rect 36747 3331 36789 3340
rect 36939 3380 36981 3389
rect 36939 3340 36940 3380
rect 36980 3340 36981 3380
rect 36939 3331 36981 3340
rect 37323 3380 37365 3389
rect 37323 3340 37324 3380
rect 37364 3340 37365 3380
rect 37323 3331 37365 3340
rect 37515 3380 37557 3389
rect 37515 3340 37516 3380
rect 37556 3340 37557 3380
rect 37515 3331 37557 3340
rect 37899 3380 37941 3389
rect 37899 3340 37900 3380
rect 37940 3340 37941 3380
rect 37899 3331 37941 3340
rect 38091 3380 38133 3389
rect 38091 3340 38092 3380
rect 38132 3340 38133 3380
rect 38091 3331 38133 3340
rect 42403 3380 42461 3381
rect 42403 3340 42412 3380
rect 42452 3340 42461 3380
rect 42403 3339 42461 3340
rect 44523 3380 44565 3389
rect 44523 3340 44524 3380
rect 44564 3340 44565 3380
rect 44523 3331 44565 3340
rect 45187 3380 45245 3381
rect 45187 3340 45196 3380
rect 45236 3340 45245 3380
rect 45187 3339 45245 3340
rect 13603 3296 13661 3297
rect 13603 3256 13612 3296
rect 13652 3256 13661 3296
rect 13603 3255 13661 3256
rect 22435 3296 22493 3297
rect 22435 3256 22444 3296
rect 22484 3256 22493 3296
rect 22435 3255 22493 3256
rect 30987 3296 31029 3305
rect 30987 3256 30988 3296
rect 31028 3256 31029 3296
rect 30987 3247 31029 3256
rect 34155 3296 34197 3305
rect 34155 3256 34156 3296
rect 34196 3256 34197 3296
rect 34155 3247 34197 3256
rect 36843 3296 36885 3305
rect 36843 3256 36844 3296
rect 36884 3256 36885 3296
rect 36843 3247 36885 3256
rect 37419 3296 37461 3305
rect 37419 3256 37420 3296
rect 37460 3256 37461 3296
rect 37419 3247 37461 3256
rect 37995 3296 38037 3305
rect 37995 3256 37996 3296
rect 38036 3256 38037 3296
rect 37995 3247 38037 3256
rect 20035 3212 20093 3213
rect 20035 3172 20044 3212
rect 20084 3172 20093 3212
rect 20035 3171 20093 3172
rect 21483 3212 21525 3221
rect 21483 3172 21484 3212
rect 21524 3172 21525 3212
rect 21483 3163 21525 3172
rect 29059 3212 29117 3213
rect 29059 3172 29068 3212
rect 29108 3172 29117 3212
rect 29059 3171 29117 3172
rect 32619 3212 32661 3221
rect 32619 3172 32620 3212
rect 32660 3172 32661 3212
rect 32619 3163 32661 3172
rect 32995 3212 33053 3213
rect 32995 3172 33004 3212
rect 33044 3172 33053 3212
rect 32995 3171 33053 3172
rect 35299 3212 35357 3213
rect 35299 3172 35308 3212
rect 35348 3172 35357 3212
rect 35299 3171 35357 3172
rect 38947 3212 39005 3213
rect 38947 3172 38956 3212
rect 38996 3172 39005 3212
rect 38947 3171 39005 3172
rect 42219 3212 42261 3221
rect 42219 3172 42220 3212
rect 42260 3172 42261 3212
rect 42219 3163 42261 3172
rect 45003 3212 45045 3221
rect 45003 3172 45004 3212
rect 45044 3172 45045 3212
rect 45003 3163 45045 3172
rect 46723 3212 46781 3213
rect 46723 3172 46732 3212
rect 46772 3172 46781 3212
rect 46723 3171 46781 3172
rect 49315 3212 49373 3213
rect 49315 3172 49324 3212
rect 49364 3172 49373 3212
rect 49315 3171 49373 3172
rect 52483 3212 52541 3213
rect 52483 3172 52492 3212
rect 52532 3172 52541 3212
rect 52483 3171 52541 3172
rect 55267 3212 55325 3213
rect 55267 3172 55276 3212
rect 55316 3172 55325 3212
rect 55267 3171 55325 3172
rect 576 3044 81984 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 81984 3044
rect 576 2980 81984 3004
rect 16867 2876 16925 2877
rect 16867 2836 16876 2876
rect 16916 2836 16925 2876
rect 16867 2835 16925 2836
rect 22531 2876 22589 2877
rect 22531 2836 22540 2876
rect 22580 2836 22589 2876
rect 22531 2835 22589 2836
rect 23211 2876 23253 2885
rect 23211 2836 23212 2876
rect 23252 2836 23253 2876
rect 23211 2827 23253 2836
rect 32043 2876 32085 2885
rect 32043 2836 32044 2876
rect 32084 2836 32085 2876
rect 32043 2827 32085 2836
rect 35203 2876 35261 2877
rect 35203 2836 35212 2876
rect 35252 2836 35261 2876
rect 35203 2835 35261 2836
rect 38179 2876 38237 2877
rect 38179 2836 38188 2876
rect 38228 2836 38237 2876
rect 38179 2835 38237 2836
rect 41347 2876 41405 2877
rect 41347 2836 41356 2876
rect 41396 2836 41405 2876
rect 41347 2835 41405 2836
rect 49123 2876 49181 2877
rect 49123 2836 49132 2876
rect 49172 2836 49181 2876
rect 49123 2835 49181 2836
rect 52003 2876 52061 2877
rect 52003 2836 52012 2876
rect 52052 2836 52061 2876
rect 52003 2835 52061 2836
rect 55171 2876 55229 2877
rect 55171 2836 55180 2876
rect 55220 2836 55229 2876
rect 55171 2835 55229 2836
rect 57763 2876 57821 2877
rect 57763 2836 57772 2876
rect 57812 2836 57821 2876
rect 57763 2835 57821 2836
rect 25795 2792 25853 2793
rect 25795 2752 25804 2792
rect 25844 2752 25853 2792
rect 25795 2751 25853 2752
rect 31171 2792 31229 2793
rect 31171 2752 31180 2792
rect 31220 2752 31229 2792
rect 31171 2751 31229 2752
rect 43075 2792 43133 2793
rect 43075 2752 43084 2792
rect 43124 2752 43133 2792
rect 43075 2751 43133 2752
rect 23395 2708 23453 2709
rect 23395 2668 23404 2708
rect 23444 2668 23453 2708
rect 23395 2667 23453 2668
rect 32227 2708 32285 2709
rect 32227 2668 32236 2708
rect 32276 2668 32285 2708
rect 32227 2667 32285 2668
rect 43275 2708 43317 2717
rect 43275 2668 43276 2708
rect 43316 2668 43317 2708
rect 43275 2659 43317 2668
rect 17163 2624 17205 2633
rect 17163 2584 17164 2624
rect 17204 2584 17205 2624
rect 17163 2575 17205 2584
rect 17259 2624 17301 2633
rect 17259 2584 17260 2624
rect 17300 2584 17301 2624
rect 17259 2575 17301 2584
rect 17539 2624 17597 2625
rect 17539 2584 17548 2624
rect 17588 2584 17597 2624
rect 17539 2583 17597 2584
rect 20139 2624 20181 2633
rect 20139 2584 20140 2624
rect 20180 2584 20181 2624
rect 20139 2575 20181 2584
rect 20515 2624 20573 2625
rect 20515 2584 20524 2624
rect 20564 2584 20573 2624
rect 20515 2583 20573 2584
rect 21379 2624 21437 2625
rect 21379 2584 21388 2624
rect 21428 2584 21437 2624
rect 21379 2583 21437 2584
rect 25123 2624 25181 2625
rect 25123 2584 25132 2624
rect 25172 2584 25181 2624
rect 25123 2583 25181 2584
rect 25419 2624 25461 2633
rect 25419 2584 25420 2624
rect 25460 2584 25461 2624
rect 25419 2575 25461 2584
rect 25995 2624 26037 2633
rect 25995 2584 25996 2624
rect 26036 2584 26037 2624
rect 25995 2575 26037 2584
rect 26371 2624 26429 2625
rect 26371 2584 26380 2624
rect 26420 2584 26429 2624
rect 26371 2583 26429 2584
rect 27235 2624 27293 2625
rect 27235 2584 27244 2624
rect 27284 2584 27293 2624
rect 27235 2583 27293 2584
rect 28779 2624 28821 2633
rect 28779 2584 28780 2624
rect 28820 2584 28821 2624
rect 28779 2575 28821 2584
rect 29155 2624 29213 2625
rect 29155 2584 29164 2624
rect 29204 2584 29213 2624
rect 29155 2583 29213 2584
rect 30019 2624 30077 2625
rect 30019 2584 30028 2624
rect 30068 2584 30077 2624
rect 30019 2583 30077 2584
rect 32811 2624 32853 2633
rect 32811 2584 32812 2624
rect 32852 2584 32853 2624
rect 32811 2575 32853 2584
rect 33187 2624 33245 2625
rect 33187 2584 33196 2624
rect 33236 2584 33245 2624
rect 33187 2583 33245 2584
rect 34051 2624 34109 2625
rect 34051 2584 34060 2624
rect 34100 2584 34109 2624
rect 34051 2583 34109 2584
rect 35787 2624 35829 2633
rect 35787 2584 35788 2624
rect 35828 2584 35829 2624
rect 35787 2575 35829 2584
rect 36163 2624 36221 2625
rect 36163 2584 36172 2624
rect 36212 2584 36221 2624
rect 36163 2583 36221 2584
rect 37027 2624 37085 2625
rect 37027 2584 37036 2624
rect 37076 2584 37085 2624
rect 37027 2583 37085 2584
rect 38955 2624 38997 2633
rect 38955 2584 38956 2624
rect 38996 2584 38997 2624
rect 38955 2575 38997 2584
rect 39331 2624 39389 2625
rect 39331 2584 39340 2624
rect 39380 2584 39389 2624
rect 39331 2583 39389 2584
rect 40195 2624 40253 2625
rect 40195 2584 40204 2624
rect 40244 2584 40253 2624
rect 40195 2583 40253 2584
rect 42403 2624 42461 2625
rect 42403 2584 42412 2624
rect 42452 2584 42461 2624
rect 42403 2583 42461 2584
rect 42699 2624 42741 2633
rect 42699 2584 42700 2624
rect 42740 2584 42741 2624
rect 42699 2575 42741 2584
rect 42795 2624 42837 2633
rect 42795 2584 42796 2624
rect 42836 2584 42837 2624
rect 42795 2575 42837 2584
rect 44419 2624 44477 2625
rect 44419 2584 44428 2624
rect 44468 2584 44477 2624
rect 44419 2583 44477 2584
rect 45283 2624 45341 2625
rect 45283 2584 45292 2624
rect 45332 2584 45341 2624
rect 45283 2583 45341 2584
rect 45675 2624 45717 2633
rect 45675 2584 45676 2624
rect 45716 2584 45717 2624
rect 45675 2575 45717 2584
rect 46731 2624 46773 2633
rect 46731 2584 46732 2624
rect 46772 2584 46773 2624
rect 46731 2575 46773 2584
rect 47107 2624 47165 2625
rect 47107 2584 47116 2624
rect 47156 2584 47165 2624
rect 47107 2583 47165 2584
rect 47971 2624 48029 2625
rect 47971 2584 47980 2624
rect 48020 2584 48029 2624
rect 47971 2583 48029 2584
rect 49611 2624 49653 2633
rect 49611 2584 49612 2624
rect 49652 2584 49653 2624
rect 49611 2575 49653 2584
rect 49987 2624 50045 2625
rect 49987 2584 49996 2624
rect 50036 2584 50045 2624
rect 49987 2583 50045 2584
rect 50851 2624 50909 2625
rect 50851 2584 50860 2624
rect 50900 2584 50909 2624
rect 50851 2583 50909 2584
rect 52779 2624 52821 2633
rect 52779 2584 52780 2624
rect 52820 2584 52821 2624
rect 52779 2575 52821 2584
rect 53155 2624 53213 2625
rect 53155 2584 53164 2624
rect 53204 2584 53213 2624
rect 53155 2583 53213 2584
rect 54044 2624 54102 2625
rect 54044 2584 54053 2624
rect 54093 2584 54102 2624
rect 54044 2583 54102 2584
rect 55371 2624 55413 2633
rect 55371 2584 55372 2624
rect 55412 2584 55413 2624
rect 55371 2575 55413 2584
rect 55747 2624 55805 2625
rect 55747 2584 55756 2624
rect 55796 2584 55805 2624
rect 55747 2583 55805 2584
rect 56611 2624 56669 2625
rect 56611 2584 56620 2624
rect 56660 2584 56669 2624
rect 56611 2583 56669 2584
rect 79843 2624 79901 2625
rect 79843 2584 79852 2624
rect 79892 2584 79901 2624
rect 79843 2583 79901 2584
rect 80707 2624 80765 2625
rect 80707 2584 80716 2624
rect 80756 2584 80765 2624
rect 80707 2583 80765 2584
rect 25515 2540 25557 2549
rect 25515 2500 25516 2540
rect 25556 2500 25557 2540
rect 25515 2491 25557 2500
rect 79467 2540 79509 2549
rect 79467 2500 79468 2540
rect 79508 2500 79509 2540
rect 79467 2491 79509 2500
rect 643 2456 701 2457
rect 643 2416 652 2456
rect 692 2416 701 2456
rect 643 2415 701 2416
rect 23211 2456 23253 2465
rect 23211 2416 23212 2456
rect 23252 2416 23253 2456
rect 23211 2407 23253 2416
rect 28387 2456 28445 2457
rect 28387 2416 28396 2456
rect 28436 2416 28445 2456
rect 28387 2415 28445 2416
rect 81859 2456 81917 2457
rect 81859 2416 81868 2456
rect 81908 2416 81917 2456
rect 81859 2415 81917 2416
rect 576 2288 81984 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 81984 2288
rect 576 2224 81984 2248
rect 26467 2120 26525 2121
rect 26467 2080 26476 2120
rect 26516 2080 26525 2120
rect 26467 2079 26525 2080
rect 30115 2120 30173 2121
rect 30115 2080 30124 2120
rect 30164 2080 30173 2120
rect 30115 2079 30173 2080
rect 34531 2120 34589 2121
rect 34531 2080 34540 2120
rect 34580 2080 34589 2120
rect 34531 2079 34589 2080
rect 34819 2120 34877 2121
rect 34819 2080 34828 2120
rect 34868 2080 34877 2120
rect 34819 2079 34877 2080
rect 40099 2120 40157 2121
rect 40099 2080 40108 2120
rect 40148 2080 40157 2120
rect 40099 2079 40157 2080
rect 42115 2120 42173 2121
rect 42115 2080 42124 2120
rect 42164 2080 42173 2120
rect 42115 2079 42173 2080
rect 44899 2120 44957 2121
rect 44899 2080 44908 2120
rect 44948 2080 44957 2120
rect 44899 2079 44957 2080
rect 22539 2036 22581 2045
rect 22539 1996 22540 2036
rect 22580 1996 22581 2036
rect 22539 1987 22581 1996
rect 23499 2036 23541 2045
rect 23499 1996 23500 2036
rect 23540 1996 23541 2036
rect 23499 1987 23541 1996
rect 31659 2036 31701 2045
rect 31659 1996 31660 2036
rect 31700 1996 31701 2036
rect 31659 1987 31701 1996
rect 41643 2036 41685 2045
rect 41643 1996 41644 2036
rect 41684 1996 41685 2036
rect 41643 1987 41685 1996
rect 19747 1952 19805 1953
rect 19747 1912 19756 1952
rect 19796 1912 19805 1952
rect 19747 1911 19805 1912
rect 20611 1952 20669 1953
rect 20611 1912 20620 1952
rect 20660 1912 20669 1952
rect 20611 1911 20669 1912
rect 21003 1952 21045 1961
rect 21003 1912 21004 1952
rect 21044 1912 21045 1952
rect 21003 1903 21045 1912
rect 22147 1952 22205 1953
rect 22147 1912 22156 1952
rect 22196 1912 22205 1952
rect 22147 1911 22205 1912
rect 22443 1952 22485 1961
rect 22443 1912 22444 1952
rect 22484 1912 22485 1952
rect 22443 1903 22485 1912
rect 23107 1952 23165 1953
rect 23107 1912 23116 1952
rect 23156 1912 23165 1952
rect 23107 1911 23165 1912
rect 23403 1952 23445 1961
rect 23403 1912 23404 1952
rect 23444 1912 23445 1952
rect 23403 1903 23445 1912
rect 24075 1952 24117 1961
rect 24075 1912 24076 1952
rect 24116 1912 24117 1952
rect 24075 1903 24117 1912
rect 24451 1952 24509 1953
rect 24451 1912 24460 1952
rect 24500 1912 24509 1952
rect 24451 1911 24509 1912
rect 25315 1952 25373 1953
rect 25315 1912 25324 1952
rect 25364 1912 25373 1952
rect 25315 1911 25373 1912
rect 26851 1952 26909 1953
rect 26851 1912 26860 1952
rect 26900 1912 26909 1952
rect 26851 1911 26909 1912
rect 27147 1952 27189 1961
rect 27147 1912 27148 1952
rect 27188 1912 27189 1952
rect 27147 1903 27189 1912
rect 27243 1952 27285 1961
rect 27243 1912 27244 1952
rect 27284 1912 27285 1952
rect 27243 1903 27285 1912
rect 27723 1952 27765 1961
rect 27723 1912 27724 1952
rect 27764 1912 27765 1952
rect 27723 1903 27765 1912
rect 28099 1952 28157 1953
rect 28099 1912 28108 1952
rect 28148 1912 28157 1952
rect 28099 1911 28157 1912
rect 28963 1952 29021 1953
rect 28963 1912 28972 1952
rect 29012 1912 29021 1952
rect 28963 1911 29021 1912
rect 31267 1952 31325 1953
rect 31267 1912 31276 1952
rect 31316 1912 31325 1952
rect 31267 1911 31325 1912
rect 31563 1952 31605 1961
rect 31563 1912 31564 1952
rect 31604 1912 31605 1952
rect 31563 1903 31605 1912
rect 32139 1952 32181 1961
rect 32139 1912 32140 1952
rect 32180 1912 32181 1952
rect 32139 1903 32181 1912
rect 32515 1952 32573 1953
rect 32515 1912 32524 1952
rect 32564 1912 32573 1952
rect 32515 1911 32573 1912
rect 33379 1952 33437 1953
rect 33379 1912 33388 1952
rect 33428 1912 33437 1952
rect 33379 1911 33437 1912
rect 35971 1952 36029 1953
rect 35971 1912 35980 1952
rect 36020 1912 36029 1952
rect 35971 1911 36029 1912
rect 36835 1952 36893 1953
rect 36835 1912 36844 1952
rect 36884 1912 36893 1952
rect 36835 1911 36893 1912
rect 37227 1952 37269 1961
rect 37227 1912 37228 1952
rect 37268 1912 37269 1952
rect 37227 1903 37269 1912
rect 37707 1952 37749 1961
rect 37707 1912 37708 1952
rect 37748 1912 37749 1952
rect 37707 1903 37749 1912
rect 38083 1952 38141 1953
rect 38083 1912 38092 1952
rect 38132 1912 38141 1952
rect 38083 1911 38141 1912
rect 38947 1952 39005 1953
rect 38947 1912 38956 1952
rect 38996 1912 39005 1952
rect 38947 1911 39005 1912
rect 41251 1952 41309 1953
rect 41251 1912 41260 1952
rect 41300 1912 41309 1952
rect 41251 1911 41309 1912
rect 41547 1952 41589 1961
rect 41547 1912 41548 1952
rect 41588 1912 41589 1952
rect 41547 1903 41589 1912
rect 43267 1952 43325 1953
rect 43267 1912 43276 1952
rect 43316 1912 43325 1952
rect 43267 1911 43325 1912
rect 44131 1952 44189 1953
rect 44131 1912 44140 1952
rect 44180 1912 44189 1952
rect 44131 1911 44189 1912
rect 44523 1952 44565 1961
rect 44523 1912 44524 1952
rect 44564 1912 44565 1952
rect 44523 1903 44565 1912
rect 46051 1952 46109 1953
rect 46051 1912 46060 1952
rect 46100 1912 46109 1952
rect 46051 1911 46109 1912
rect 46915 1952 46973 1953
rect 46915 1912 46924 1952
rect 46964 1912 46973 1952
rect 46915 1911 46973 1912
rect 47307 1952 47349 1961
rect 47307 1912 47308 1952
rect 47348 1912 47349 1952
rect 47307 1903 47349 1912
rect 48643 1952 48701 1953
rect 48643 1912 48652 1952
rect 48692 1912 48701 1952
rect 48643 1911 48701 1912
rect 49507 1952 49565 1953
rect 49507 1912 49516 1952
rect 49556 1912 49565 1952
rect 49507 1911 49565 1912
rect 49899 1952 49941 1961
rect 49899 1912 49900 1952
rect 49940 1912 49941 1952
rect 49899 1903 49941 1912
rect 51235 1952 51293 1953
rect 51235 1912 51244 1952
rect 51284 1912 51293 1952
rect 51235 1911 51293 1912
rect 52099 1952 52157 1953
rect 52099 1912 52108 1952
rect 52148 1912 52157 1952
rect 52099 1911 52157 1912
rect 52491 1952 52533 1961
rect 52491 1912 52492 1952
rect 52532 1912 52533 1952
rect 52491 1903 52533 1912
rect 53827 1952 53885 1953
rect 53827 1912 53836 1952
rect 53876 1912 53885 1952
rect 53827 1911 53885 1912
rect 54691 1952 54749 1953
rect 54691 1912 54700 1952
rect 54740 1912 54749 1952
rect 54691 1911 54749 1912
rect 55083 1952 55125 1961
rect 55083 1912 55084 1952
rect 55124 1912 55125 1952
rect 55083 1903 55125 1912
rect 72747 1952 72789 1961
rect 72747 1912 72748 1952
rect 72788 1912 72789 1952
rect 72747 1903 72789 1912
rect 74083 1952 74141 1953
rect 74083 1912 74092 1952
rect 74132 1912 74141 1952
rect 74083 1911 74141 1912
rect 78595 1952 78653 1953
rect 78595 1912 78604 1952
rect 78644 1912 78653 1952
rect 78595 1911 78653 1912
rect 78891 1952 78933 1961
rect 78891 1912 78892 1952
rect 78932 1912 78933 1952
rect 78891 1903 78933 1912
rect 78987 1952 79029 1961
rect 78987 1912 78988 1952
rect 79028 1912 79029 1952
rect 78987 1903 79029 1912
rect 79467 1952 79509 1961
rect 79467 1912 79468 1952
rect 79508 1912 79509 1952
rect 79467 1903 79509 1912
rect 79843 1952 79901 1953
rect 79843 1912 79852 1952
rect 79892 1912 79901 1952
rect 79843 1911 79901 1912
rect 80707 1952 80765 1953
rect 80707 1912 80716 1952
rect 80756 1912 80765 1952
rect 80707 1911 80765 1912
rect 23779 1784 23837 1785
rect 23779 1744 23788 1784
rect 23828 1744 23837 1784
rect 23779 1743 23837 1744
rect 27523 1784 27581 1785
rect 27523 1744 27532 1784
rect 27572 1744 27581 1784
rect 27523 1743 27581 1744
rect 31939 1784 31997 1785
rect 31939 1744 31948 1784
rect 31988 1744 31997 1784
rect 31939 1743 31997 1744
rect 41923 1784 41981 1785
rect 41923 1744 41932 1784
rect 41972 1744 41981 1784
rect 41923 1743 41981 1744
rect 79267 1784 79325 1785
rect 79267 1744 79276 1784
rect 79316 1744 79325 1784
rect 79267 1743 79325 1744
rect 18595 1700 18653 1701
rect 18595 1660 18604 1700
rect 18644 1660 18653 1700
rect 18595 1659 18653 1660
rect 22819 1700 22877 1701
rect 22819 1660 22828 1700
rect 22868 1660 22877 1700
rect 22819 1659 22877 1660
rect 44899 1700 44957 1701
rect 44899 1660 44908 1700
rect 44948 1660 44957 1700
rect 44899 1659 44957 1660
rect 47491 1700 47549 1701
rect 47491 1660 47500 1700
rect 47540 1660 47549 1700
rect 47491 1659 47549 1660
rect 50083 1700 50141 1701
rect 50083 1660 50092 1700
rect 50132 1660 50141 1700
rect 50083 1659 50141 1660
rect 52675 1700 52733 1701
rect 52675 1660 52684 1700
rect 52724 1660 52733 1700
rect 52675 1659 52733 1660
rect 81859 1700 81917 1701
rect 81859 1660 81868 1700
rect 81908 1660 81917 1700
rect 81859 1659 81917 1660
rect 576 1532 81984 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 81984 1532
rect 576 1468 81984 1492
rect 20323 1364 20381 1365
rect 20323 1324 20332 1364
rect 20372 1324 20381 1364
rect 20323 1323 20381 1324
rect 25027 1364 25085 1365
rect 25027 1324 25036 1364
rect 25076 1324 25085 1364
rect 25027 1323 25085 1324
rect 32707 1364 32765 1365
rect 32707 1324 32716 1364
rect 32756 1324 32765 1364
rect 32707 1323 32765 1324
rect 35395 1364 35453 1365
rect 35395 1324 35404 1364
rect 35444 1324 35453 1364
rect 35395 1323 35453 1324
rect 37603 1364 37661 1365
rect 37603 1324 37612 1364
rect 37652 1324 37661 1364
rect 37603 1323 37661 1324
rect 42883 1364 42941 1365
rect 42883 1324 42892 1364
rect 42932 1324 42941 1364
rect 42883 1323 42941 1324
rect 45091 1364 45149 1365
rect 45091 1324 45100 1364
rect 45140 1324 45149 1364
rect 45091 1323 45149 1324
rect 47587 1364 47645 1365
rect 47587 1324 47596 1364
rect 47636 1324 47645 1364
rect 47587 1323 47645 1324
rect 50275 1364 50333 1365
rect 50275 1324 50284 1364
rect 50324 1324 50333 1364
rect 50275 1323 50333 1324
rect 52771 1364 52829 1365
rect 52771 1324 52780 1364
rect 52820 1324 52829 1364
rect 52771 1323 52829 1324
rect 79555 1364 79613 1365
rect 79555 1324 79564 1364
rect 79604 1324 79613 1364
rect 79555 1323 79613 1324
rect 30115 1280 30173 1281
rect 30115 1240 30124 1280
rect 30164 1240 30173 1280
rect 30115 1239 30173 1240
rect 40291 1280 40349 1281
rect 40291 1240 40300 1280
rect 40340 1240 40349 1280
rect 40291 1239 40349 1240
rect 19651 1112 19709 1113
rect 19651 1072 19660 1112
rect 19700 1072 19709 1112
rect 19651 1071 19709 1072
rect 19947 1112 19989 1121
rect 19947 1072 19948 1112
rect 19988 1072 19989 1112
rect 19947 1063 19989 1072
rect 20043 1112 20085 1121
rect 20043 1072 20044 1112
rect 20084 1072 20085 1112
rect 20043 1063 20085 1072
rect 22635 1112 22677 1121
rect 22635 1072 22636 1112
rect 22676 1072 22677 1112
rect 22635 1063 22677 1072
rect 23011 1112 23069 1113
rect 23011 1072 23020 1112
rect 23060 1072 23069 1112
rect 23011 1071 23069 1072
rect 23875 1112 23933 1113
rect 23875 1072 23884 1112
rect 23924 1072 23933 1112
rect 23875 1071 23933 1072
rect 29443 1112 29501 1113
rect 29443 1072 29452 1112
rect 29492 1072 29501 1112
rect 29443 1071 29501 1072
rect 29739 1112 29781 1121
rect 29739 1072 29740 1112
rect 29780 1072 29781 1112
rect 29739 1063 29781 1072
rect 29835 1112 29877 1121
rect 29835 1072 29836 1112
rect 29876 1072 29877 1112
rect 29835 1063 29877 1072
rect 30315 1112 30357 1121
rect 30315 1072 30316 1112
rect 30356 1072 30357 1112
rect 30315 1063 30357 1072
rect 30691 1112 30749 1113
rect 30691 1072 30700 1112
rect 30740 1072 30749 1112
rect 30691 1071 30749 1072
rect 31555 1112 31613 1113
rect 31555 1072 31564 1112
rect 31604 1072 31613 1112
rect 31555 1071 31613 1072
rect 35691 1112 35733 1121
rect 35691 1072 35692 1112
rect 35732 1072 35733 1112
rect 35691 1063 35733 1072
rect 35787 1112 35829 1121
rect 35787 1072 35788 1112
rect 35828 1072 35829 1112
rect 35787 1063 35829 1072
rect 36067 1112 36125 1113
rect 36067 1072 36076 1112
rect 36116 1072 36125 1112
rect 36067 1071 36125 1072
rect 37899 1112 37941 1121
rect 37899 1072 37900 1112
rect 37940 1072 37941 1112
rect 37899 1063 37941 1072
rect 37995 1112 38037 1121
rect 37995 1072 37996 1112
rect 38036 1072 38037 1112
rect 37995 1063 38037 1072
rect 38275 1112 38333 1113
rect 38275 1072 38284 1112
rect 38324 1072 38333 1112
rect 38275 1071 38333 1072
rect 39619 1112 39677 1113
rect 39619 1072 39628 1112
rect 39668 1072 39677 1112
rect 39619 1071 39677 1072
rect 39915 1112 39957 1121
rect 39915 1072 39916 1112
rect 39956 1072 39957 1112
rect 39915 1063 39957 1072
rect 40011 1112 40053 1121
rect 40011 1072 40012 1112
rect 40052 1072 40053 1112
rect 40011 1063 40053 1072
rect 40491 1112 40533 1121
rect 40491 1072 40492 1112
rect 40532 1072 40533 1112
rect 40491 1063 40533 1072
rect 40867 1112 40925 1113
rect 40867 1072 40876 1112
rect 40916 1072 40925 1112
rect 40867 1071 40925 1072
rect 41731 1112 41789 1113
rect 41731 1072 41740 1112
rect 41780 1072 41789 1112
rect 41731 1071 41789 1072
rect 44419 1112 44477 1113
rect 44419 1072 44428 1112
rect 44468 1072 44477 1112
rect 44419 1071 44477 1072
rect 44715 1112 44757 1121
rect 44715 1072 44716 1112
rect 44756 1072 44757 1112
rect 44715 1063 44757 1072
rect 44811 1112 44853 1121
rect 44811 1072 44812 1112
rect 44852 1072 44853 1112
rect 44811 1063 44853 1072
rect 46915 1112 46973 1113
rect 46915 1072 46924 1112
rect 46964 1072 46973 1112
rect 46915 1071 46973 1072
rect 47211 1112 47253 1121
rect 47211 1072 47212 1112
rect 47252 1072 47253 1112
rect 47211 1063 47253 1072
rect 49603 1112 49661 1113
rect 49603 1072 49612 1112
rect 49652 1072 49661 1112
rect 49603 1071 49661 1072
rect 49899 1112 49941 1121
rect 49899 1072 49900 1112
rect 49940 1072 49941 1112
rect 49899 1063 49941 1072
rect 49995 1112 50037 1121
rect 49995 1072 49996 1112
rect 50036 1072 50037 1112
rect 49995 1063 50037 1072
rect 52099 1112 52157 1113
rect 52099 1072 52108 1112
rect 52148 1072 52157 1112
rect 52099 1071 52157 1072
rect 52395 1112 52437 1121
rect 52395 1072 52396 1112
rect 52436 1072 52437 1112
rect 52395 1063 52437 1072
rect 52491 1112 52533 1121
rect 52491 1072 52492 1112
rect 52532 1072 52533 1112
rect 52491 1063 52533 1072
rect 79947 1112 79989 1121
rect 79947 1072 79948 1112
rect 79988 1072 79989 1112
rect 79947 1063 79989 1072
rect 80227 1112 80285 1113
rect 80227 1072 80236 1112
rect 80276 1072 80285 1112
rect 80227 1071 80285 1072
rect 47307 1028 47349 1037
rect 47307 988 47308 1028
rect 47348 988 47349 1028
rect 47307 979 47349 988
rect 79851 1028 79893 1037
rect 79851 988 79852 1028
rect 79892 988 79893 1028
rect 79851 979 79893 988
rect 576 776 81984 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 81984 776
rect 576 712 81984 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 652 38116 692 38156
rect 844 37948 884 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 12172 35848 12212 35888
rect 12460 35848 12500 35888
rect 13324 35848 13364 35888
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 32620 35176 32660 35216
rect 32716 35176 32756 35216
rect 33004 35176 33044 35216
rect 33772 35176 33812 35216
rect 34060 35176 34100 35216
rect 34156 35176 34196 35216
rect 50284 35176 50324 35216
rect 15052 35092 15092 35132
rect 82252 35092 82292 35132
rect 15244 34924 15284 34964
rect 32332 34924 32372 34964
rect 34444 34924 34484 34964
rect 82444 34924 82484 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 22732 34504 22772 34544
rect 28972 34504 29012 34544
rect 34732 34504 34772 34544
rect 38188 34504 38228 34544
rect 49996 34504 50036 34544
rect 50572 34504 50612 34544
rect 52204 34504 52244 34544
rect 83212 34504 83252 34544
rect 20812 34420 20852 34460
rect 21196 34420 21236 34460
rect 21580 34420 21620 34460
rect 22924 34420 22964 34460
rect 45580 34420 45620 34460
rect 15052 34336 15092 34376
rect 15820 34336 15860 34376
rect 16684 34336 16724 34376
rect 18412 34336 18452 34376
rect 19276 34336 19316 34376
rect 22060 34336 22100 34376
rect 22348 34336 22388 34376
rect 29356 34336 29396 34376
rect 29644 34336 29684 34376
rect 32332 34336 32372 34376
rect 32716 34336 32756 34376
rect 33580 34336 33620 34376
rect 36940 34336 36980 34376
rect 37900 34336 37940 34376
rect 38572 34336 38612 34376
rect 38860 34336 38900 34376
rect 49324 34336 49364 34376
rect 49612 34336 49652 34376
rect 50284 34336 50324 34376
rect 51532 34336 51572 34376
rect 51820 34336 51860 34376
rect 81196 34336 81236 34376
rect 82060 34336 82100 34376
rect 15436 34252 15476 34292
rect 18028 34252 18068 34292
rect 22444 34252 22484 34292
rect 29260 34252 29300 34292
rect 38476 34252 38516 34292
rect 49708 34252 49748 34292
rect 51916 34252 51956 34292
rect 80812 34252 80852 34292
rect 14668 34168 14708 34208
rect 17836 34168 17876 34208
rect 20428 34168 20468 34208
rect 21004 34168 21044 34208
rect 21388 34168 21428 34208
rect 21772 34168 21812 34208
rect 23116 34168 23156 34208
rect 45388 34168 45428 34208
rect 50764 34168 50804 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 29548 33832 29588 33872
rect 40300 33832 40340 33872
rect 52492 33832 52532 33872
rect 17356 33748 17396 33788
rect 21100 33748 21140 33788
rect 25324 33748 25364 33788
rect 37900 33748 37940 33788
rect 50092 33748 50132 33788
rect 81868 33748 81908 33788
rect 13996 33664 14036 33704
rect 14380 33664 14420 33704
rect 15244 33664 15284 33704
rect 16972 33664 17012 33704
rect 20716 33664 20756 33704
rect 21004 33664 21044 33704
rect 17260 33622 17300 33662
rect 21772 33664 21812 33704
rect 22636 33664 22676 33704
rect 24076 33664 24116 33704
rect 24940 33664 24980 33704
rect 25612 33664 25652 33704
rect 26572 33664 26612 33704
rect 27148 33664 27188 33704
rect 27532 33664 27572 33704
rect 28396 33664 28436 33704
rect 30220 33664 30260 33704
rect 30508 33664 30548 33704
rect 30604 33664 30644 33704
rect 31084 33664 31124 33704
rect 31468 33664 31508 33704
rect 32332 33664 32372 33704
rect 33772 33664 33812 33704
rect 34060 33664 34100 33704
rect 34156 33664 34196 33704
rect 35308 33664 35348 33704
rect 35692 33664 35732 33704
rect 36556 33664 36596 33704
rect 38284 33664 38324 33704
rect 39148 33664 39188 33704
rect 41644 33664 41684 33704
rect 42028 33664 42068 33704
rect 42892 33664 42932 33704
rect 44908 33664 44948 33704
rect 45292 33664 45332 33704
rect 46156 33664 46196 33704
rect 47500 33664 47540 33704
rect 47884 33664 47924 33704
rect 48748 33664 48788 33704
rect 50476 33664 50516 33704
rect 51340 33664 51380 33704
rect 52684 33664 52724 33704
rect 81964 33664 82004 33704
rect 82252 33664 82292 33704
rect 33484 33580 33524 33620
rect 17644 33496 17684 33536
rect 30892 33496 30932 33536
rect 34444 33496 34484 33536
rect 81580 33496 81620 33536
rect 16396 33412 16436 33452
rect 21388 33412 21428 33452
rect 21964 33412 22004 33452
rect 22924 33412 22964 33452
rect 29548 33412 29588 33452
rect 37708 33412 37748 33452
rect 44044 33412 44084 33452
rect 47308 33412 47348 33452
rect 49900 33412 49940 33452
rect 52492 33412 52532 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 12268 33076 12308 33116
rect 14476 33076 14516 33116
rect 15340 33076 15380 33116
rect 20524 33076 20564 33116
rect 23692 33076 23732 33116
rect 27148 33076 27188 33116
rect 31756 33076 31796 33116
rect 36748 33076 36788 33116
rect 41260 33076 41300 33116
rect 42316 33076 42356 33116
rect 45292 33076 45332 33116
rect 47212 33076 47252 33116
rect 9580 32992 9620 33032
rect 17932 32992 17972 33032
rect 43084 32992 43124 33032
rect 69772 32992 69812 33032
rect 42124 32908 42164 32948
rect 5740 32824 5780 32864
rect 6604 32824 6644 32864
rect 8908 32824 8948 32864
rect 9196 32824 9236 32864
rect 9292 32824 9332 32864
rect 9868 32824 9908 32864
rect 10252 32824 10292 32864
rect 11116 32824 11156 32864
rect 13804 32824 13844 32864
rect 14092 32824 14132 32864
rect 15724 32824 15764 32864
rect 16012 32824 16052 32864
rect 17216 32824 17256 32864
rect 17548 32824 17588 32864
rect 17644 32824 17684 32864
rect 18124 32824 18164 32864
rect 18508 32824 18548 32864
rect 19372 32824 19412 32864
rect 21292 32824 21332 32864
rect 21676 32824 21716 32864
rect 22540 32824 22580 32864
rect 25516 32824 25556 32864
rect 27532 32824 27572 32864
rect 27820 32824 27860 32864
rect 29356 32824 29396 32864
rect 29740 32824 29780 32864
rect 30604 32824 30644 32864
rect 33100 32824 33140 32864
rect 33964 32824 34004 32864
rect 34348 32824 34388 32864
rect 34732 32824 34772 32864
rect 35596 32824 35636 32864
rect 36940 32824 36980 32864
rect 37324 32824 37364 32864
rect 38764 32824 38804 32864
rect 40588 32824 40628 32864
rect 40876 32824 40916 32864
rect 40972 32824 41012 32864
rect 44716 32824 44756 32864
rect 45580 32824 45620 32864
rect 45676 32824 45716 32864
rect 45964 32824 46004 32864
rect 47596 32824 47636 32864
rect 47884 32824 47924 32864
rect 49132 32824 49172 32864
rect 50284 32824 50324 32864
rect 50764 32824 50804 32864
rect 51724 32824 51764 32864
rect 51916 32824 51956 32864
rect 52300 32824 52340 32864
rect 53164 32824 53204 32864
rect 64972 32824 65012 32864
rect 65260 32824 65300 32864
rect 66124 32824 66164 32864
rect 70060 32824 70100 32864
rect 5356 32740 5396 32780
rect 14188 32740 14228 32780
rect 15628 32740 15668 32780
rect 27436 32740 27476 32780
rect 47500 32740 47540 32780
rect 7756 32656 7796 32696
rect 12268 32656 12308 32696
rect 23692 32656 23732 32696
rect 31756 32656 31796 32696
rect 42700 32656 42740 32696
rect 48652 32656 48692 32696
rect 49900 32656 49940 32696
rect 54316 32656 54356 32696
rect 65740 32656 65780 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 80812 32152 80852 32192
rect 81196 32152 81236 32192
rect 82060 32152 82100 32192
rect 1900 32068 1940 32108
rect 83212 31984 83252 32024
rect 2092 31900 2132 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 1516 31564 1556 31604
rect 4972 31564 5012 31604
rect 81388 31564 81428 31604
rect 1900 31480 1940 31520
rect 1324 31396 1364 31436
rect 1708 31396 1748 31436
rect 2764 31312 2804 31352
rect 3628 31312 3668 31352
rect 5260 31312 5300 31352
rect 5356 31308 5396 31348
rect 5680 31312 5720 31352
rect 81676 31312 81716 31352
rect 81772 31312 81812 31352
rect 82060 31312 82100 31352
rect 2380 31228 2420 31268
rect 4780 31144 4820 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 1228 30640 1268 30680
rect 1612 30640 1652 30680
rect 2476 30640 2516 30680
rect 78316 30640 78356 30680
rect 78700 30640 78740 30680
rect 81868 30640 81908 30680
rect 82252 30640 82292 30680
rect 82540 30472 82580 30512
rect 3628 30388 3668 30428
rect 78892 30388 78932 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 1900 30052 1940 30092
rect 2092 29884 2132 29924
rect 1228 29800 1268 29840
rect 1516 29800 1556 29840
rect 2188 29800 2228 29840
rect 2380 29800 2420 29840
rect 2476 29800 2516 29840
rect 2572 29800 2612 29840
rect 2668 29800 2708 29840
rect 3820 29800 3860 29840
rect 4684 29800 4724 29840
rect 1612 29716 1652 29756
rect 3436 29716 3476 29756
rect 5836 29632 5876 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 2668 29296 2708 29336
rect 2764 29296 2804 29336
rect 3532 29296 3572 29336
rect 3820 29296 3860 29336
rect 2860 29212 2900 29252
rect 1516 29128 1556 29168
rect 1708 29128 1748 29168
rect 1900 29128 1940 29168
rect 2092 29128 2132 29168
rect 2188 29128 2228 29168
rect 2956 29128 2996 29168
rect 3052 29128 3092 29168
rect 3340 29128 3380 29168
rect 3436 29128 3476 29168
rect 3628 29128 3668 29168
rect 3916 29128 3956 29168
rect 4588 29128 4628 29168
rect 4780 29128 4820 29168
rect 5644 29128 5684 29168
rect 1900 28960 1940 29000
rect 1516 28876 1556 28916
rect 4108 28876 4148 28916
rect 5068 28876 5108 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 3148 28540 3188 28580
rect 3916 28456 3956 28496
rect 748 28288 788 28328
rect 1132 28288 1172 28328
rect 1996 28288 2036 28328
rect 3436 28288 3476 28328
rect 3532 28288 3572 28328
rect 3628 28288 3668 28328
rect 3724 28288 3764 28328
rect 4108 28288 4148 28328
rect 4300 28288 4340 28328
rect 4588 28288 4628 28328
rect 4780 28288 4820 28328
rect 5644 28288 5684 28328
rect 4204 28120 4244 28160
rect 4492 28120 4532 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 2092 27784 2132 27824
rect 2764 27784 2804 27824
rect 83212 27784 83252 27824
rect 1804 27700 1844 27740
rect 1996 27616 2036 27656
rect 2092 27616 2132 27656
rect 2860 27616 2900 27656
rect 4588 27616 4628 27656
rect 5452 27616 5492 27656
rect 5836 27616 5876 27656
rect 80812 27616 80852 27656
rect 81196 27616 81236 27656
rect 82060 27616 82100 27656
rect 3436 27532 3476 27572
rect 3052 27448 3092 27488
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 4684 27028 4724 27068
rect 81388 27028 81428 27068
rect 4108 26944 4148 26984
rect 1036 26860 1076 26900
rect 1420 26776 1460 26816
rect 1516 26776 1556 26816
rect 1708 26776 1748 26816
rect 2380 26776 2420 26816
rect 2668 26776 2708 26816
rect 3340 26776 3380 26816
rect 3436 26776 3476 26816
rect 3532 26776 3572 26816
rect 3628 26776 3668 26816
rect 4012 26776 4052 26816
rect 4108 26776 4148 26816
rect 4300 26776 4340 26816
rect 4492 26776 4532 26816
rect 4684 26776 4724 26816
rect 81676 26776 81716 26816
rect 81772 26776 81812 26816
rect 82060 26776 82100 26816
rect 1228 26608 1268 26648
rect 1612 26608 1652 26648
rect 2572 26608 2612 26648
rect 3820 26608 3860 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 3052 26272 3092 26312
rect 3340 26272 3380 26312
rect 652 26188 692 26228
rect 3436 26188 3476 26228
rect 1036 26104 1076 26144
rect 1900 26104 1940 26144
rect 3532 26104 3572 26144
rect 3628 26104 3668 26144
rect 3820 26104 3860 26144
rect 3916 26104 3956 26144
rect 4108 26104 4148 26144
rect 4300 26104 4340 26144
rect 4492 26104 4532 26144
rect 4684 26104 4724 26144
rect 4876 26104 4916 26144
rect 3340 25936 3380 25976
rect 3916 25936 3956 25976
rect 4300 25852 4340 25892
rect 4876 25852 4916 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 1708 25516 1748 25556
rect 652 25348 692 25388
rect 1708 25264 1748 25304
rect 1900 25264 1940 25304
rect 1996 25264 2036 25304
rect 3820 25264 3860 25304
rect 4684 25264 4724 25304
rect 3436 25180 3476 25220
rect 844 25096 884 25136
rect 5836 25096 5876 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 844 24760 884 24800
rect 4300 24760 4340 24800
rect 3244 24676 3284 24716
rect 2188 24592 2228 24632
rect 3340 24592 3380 24632
rect 3724 24592 3764 24632
rect 3916 24592 3956 24632
rect 4108 24592 4148 24632
rect 4396 24592 4436 24632
rect 79756 24592 79796 24632
rect 652 24508 692 24548
rect 1036 24508 1076 24548
rect 81772 24508 81812 24548
rect 4108 24424 4148 24464
rect 1228 24340 1268 24380
rect 2092 24340 2132 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 5260 24004 5300 24044
rect 1324 23920 1364 23960
rect 844 23752 884 23792
rect 1036 23752 1076 23792
rect 1132 23745 1172 23785
rect 1612 23752 1652 23792
rect 1708 23752 1748 23792
rect 1996 23752 2036 23792
rect 2092 23752 2132 23792
rect 2860 23794 2900 23834
rect 3244 23752 3284 23792
rect 4108 23752 4148 23792
rect 1804 23580 1844 23620
rect 2284 23584 2324 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 3052 23248 3092 23288
rect 4396 23248 4436 23288
rect 652 23080 692 23120
rect 1036 23080 1076 23120
rect 1900 23080 1940 23120
rect 4204 22996 4244 23036
rect 4588 22996 4628 23036
rect 4780 22828 4820 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 1228 22492 1268 22532
rect 1036 22324 1076 22364
rect 3820 22240 3860 22280
rect 4684 22240 4724 22280
rect 3436 22156 3476 22196
rect 652 22072 692 22112
rect 5836 22072 5876 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 4300 21652 4340 21692
rect 4396 21568 4436 21608
rect 4684 21568 4724 21608
rect 4012 21400 4052 21440
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 5164 20980 5204 21020
rect 3148 20728 3188 20768
rect 4012 20728 4052 20768
rect 2764 20644 2804 20684
rect 652 20560 692 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 652 20224 692 20264
rect 2764 20140 2804 20180
rect 81388 20140 81428 20180
rect 2860 20056 2900 20096
rect 3148 20056 3188 20096
rect 3436 20056 3476 20096
rect 3820 20056 3860 20096
rect 4684 20056 4724 20096
rect 81004 20056 81044 20096
rect 81292 20056 81332 20096
rect 81868 20056 81908 20096
rect 82252 20056 82292 20096
rect 83116 20056 83156 20096
rect 5836 19972 5876 20012
rect 84268 19972 84308 20012
rect 2476 19888 2516 19928
rect 81676 19888 81716 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4300 19468 4340 19508
rect 81484 19468 81524 19508
rect 2092 19300 2132 19340
rect 81292 19300 81332 19340
rect 4588 19216 4628 19256
rect 4684 19216 4724 19256
rect 4972 19216 5012 19256
rect 652 19048 692 19088
rect 1900 19048 1940 19088
rect 81484 19048 81524 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 844 18544 884 18584
rect 1228 18544 1268 18584
rect 2092 18544 2132 18584
rect 3436 18544 3476 18584
rect 3820 18544 3860 18584
rect 4684 18544 4724 18584
rect 3244 18292 3284 18332
rect 5836 18292 5876 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 1612 17956 1652 17996
rect 3916 17956 3956 17996
rect 1420 17788 1460 17828
rect 2668 17788 2708 17828
rect 3244 17788 3284 17828
rect 1900 17704 1940 17744
rect 1996 17704 2036 17744
rect 2284 17704 2324 17744
rect 4300 17704 4340 17744
rect 4588 17704 4628 17744
rect 4204 17620 4244 17660
rect 652 17536 692 17576
rect 1228 17536 1268 17576
rect 2860 17536 2900 17576
rect 3052 17536 3092 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 652 17200 692 17240
rect 1036 17200 1076 17240
rect 1996 17032 2036 17072
rect 2380 17032 2420 17072
rect 3244 17032 3284 17072
rect 74188 17032 74228 17072
rect 75628 16948 75668 16988
rect 4396 16780 4436 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 1612 16444 1652 16484
rect 2572 16444 2612 16484
rect 5836 16444 5876 16484
rect 1228 16276 1268 16316
rect 2764 16276 2804 16316
rect 1900 16192 1940 16232
rect 1996 16192 2036 16232
rect 2284 16192 2324 16232
rect 3820 16192 3860 16232
rect 4684 16192 4724 16232
rect 3436 16108 3476 16148
rect 652 16024 692 16064
rect 1420 16024 1460 16064
rect 2572 16024 2612 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 81868 15688 81908 15728
rect 4492 15604 4532 15644
rect 1420 15520 1460 15560
rect 1516 15520 1556 15560
rect 1612 15520 1652 15560
rect 1996 15520 2036 15560
rect 2188 15520 2228 15560
rect 4588 15520 4628 15560
rect 4876 15520 4916 15560
rect 79468 15520 79508 15560
rect 79852 15520 79892 15560
rect 80716 15520 80756 15560
rect 844 15436 884 15476
rect 2092 15436 2132 15476
rect 1804 15352 1844 15392
rect 4204 15352 4244 15392
rect 652 15268 692 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 3244 14932 3284 14972
rect 80428 14932 80468 14972
rect 1228 14680 1268 14720
rect 2092 14680 2132 14720
rect 3820 14680 3860 14720
rect 4684 14680 4724 14720
rect 80716 14680 80756 14720
rect 80812 14680 80852 14720
rect 81100 14680 81140 14720
rect 844 14596 884 14636
rect 3436 14596 3476 14636
rect 5836 14512 5876 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 1612 14092 1652 14132
rect 3916 14092 3956 14132
rect 1708 14008 1748 14048
rect 1996 14008 2036 14048
rect 4012 14008 4052 14048
rect 4300 14008 4340 14048
rect 844 13924 884 13964
rect 76396 13924 76436 13964
rect 652 13840 692 13880
rect 1324 13840 1364 13880
rect 3628 13840 3668 13880
rect 76204 13756 76244 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 1900 13420 1940 13460
rect 5836 13420 5876 13460
rect 81868 13420 81908 13460
rect 76588 13336 76628 13376
rect 844 13252 884 13292
rect 1516 13168 1556 13208
rect 1708 13168 1748 13208
rect 1996 13157 2036 13197
rect 3820 13168 3860 13208
rect 4684 13168 4724 13208
rect 75916 13168 75956 13208
rect 76204 13168 76244 13208
rect 76780 13168 76820 13208
rect 77164 13168 77204 13208
rect 78028 13168 78068 13208
rect 79852 13168 79892 13208
rect 80716 13168 80756 13208
rect 3436 13084 3476 13124
rect 76300 13084 76340 13124
rect 79468 13084 79508 13124
rect 652 13000 692 13040
rect 1612 13000 1652 13040
rect 75628 13000 75668 13040
rect 79180 13000 79220 13040
rect 81868 13000 81908 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 77260 12664 77300 12704
rect 4204 12580 4244 12620
rect 80236 12580 80276 12620
rect 844 12496 884 12536
rect 1132 12496 1172 12536
rect 1324 12496 1364 12536
rect 1708 12496 1748 12536
rect 2572 12496 2612 12536
rect 4300 12496 4340 12536
rect 4588 12496 4628 12536
rect 79084 12496 79124 12536
rect 79372 12496 79412 12536
rect 79468 12496 79508 12536
rect 80332 12496 80372 12536
rect 80620 12496 80660 12536
rect 940 12412 980 12452
rect 77452 12412 77492 12452
rect 3916 12328 3956 12368
rect 79948 12328 79988 12368
rect 3724 12244 3764 12284
rect 79756 12244 79796 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 652 11908 692 11948
rect 1324 11908 1364 11948
rect 844 11740 884 11780
rect 5836 11740 5876 11780
rect 81868 11740 81908 11780
rect 1612 11656 1652 11696
rect 1708 11656 1748 11696
rect 1996 11656 2036 11696
rect 3820 11656 3860 11696
rect 4684 11656 4724 11696
rect 79468 11656 79508 11696
rect 79852 11656 79892 11696
rect 80716 11656 80756 11696
rect 3436 11572 3476 11612
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 652 11152 692 11192
rect 1708 11152 1748 11192
rect 1420 11068 1460 11108
rect 4012 11068 4052 11108
rect 1612 10984 1652 11024
rect 4108 10984 4148 11024
rect 4396 10984 4436 11024
rect 80140 10984 80180 11024
rect 80236 10984 80276 11024
rect 80524 10984 80564 11024
rect 844 10900 884 10940
rect 1228 10900 1268 10940
rect 3724 10816 3764 10856
rect 1036 10732 1076 10772
rect 79852 10732 79892 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 5836 10396 5876 10436
rect 3244 10228 3284 10268
rect 81868 10228 81908 10268
rect 1228 10144 1268 10184
rect 2092 10144 2132 10184
rect 3820 10144 3860 10184
rect 4684 10144 4724 10184
rect 79468 10144 79508 10184
rect 79852 10144 79892 10184
rect 80716 10144 80756 10184
rect 844 10060 884 10100
rect 3436 10060 3476 10100
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 652 9640 692 9680
rect 1036 9640 1076 9680
rect 1324 9640 1364 9680
rect 1804 9556 1844 9596
rect 4300 9556 4340 9596
rect 1228 9472 1268 9512
rect 1900 9472 1940 9512
rect 2188 9472 2228 9512
rect 4396 9472 4436 9512
rect 4684 9472 4724 9512
rect 844 9388 884 9428
rect 1516 9304 1556 9344
rect 4012 9304 4052 9344
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 652 8884 692 8924
rect 5260 8884 5300 8924
rect 1420 8800 1460 8840
rect 2668 8800 2708 8840
rect 844 8716 884 8756
rect 1612 8632 1652 8672
rect 1996 8632 2036 8672
rect 2284 8632 2324 8672
rect 2380 8632 2420 8672
rect 2860 8632 2900 8672
rect 3244 8632 3284 8672
rect 4108 8632 4148 8672
rect 1036 8464 1076 8504
rect 1708 8464 1748 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 652 8128 692 8168
rect 3436 7960 3476 8000
rect 3820 7960 3860 8000
rect 4684 7960 4724 8000
rect 5836 7708 5876 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 3532 7372 3572 7412
rect 1324 7120 1364 7160
rect 1420 7120 1460 7160
rect 1612 7120 1652 7160
rect 1708 7120 1748 7160
rect 1996 7120 2036 7160
rect 3820 7120 3860 7160
rect 3916 7120 3956 7160
rect 4204 7120 4244 7160
rect 1900 7036 1940 7076
rect 652 6952 692 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 81868 6616 81908 6656
rect 79468 6448 79508 6488
rect 79852 6448 79892 6488
rect 80716 6448 80756 6488
rect 81868 6196 81908 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 80140 5860 80180 5900
rect 5836 5692 5876 5732
rect 3820 5608 3860 5648
rect 4684 5608 4724 5648
rect 80428 5608 80468 5648
rect 80524 5608 80564 5648
rect 80812 5608 80852 5648
rect 3436 5524 3476 5564
rect 652 5440 692 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 652 5104 692 5144
rect 4492 5020 4532 5060
rect 4588 4936 4628 4976
rect 4876 4936 4916 4976
rect 80140 4936 80180 4976
rect 80236 4936 80276 4976
rect 80524 4936 80564 4976
rect 4204 4768 4244 4808
rect 79852 4684 79892 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 81868 4348 81908 4388
rect 79468 4096 79508 4136
rect 79852 4096 79892 4136
rect 80716 4096 80756 4136
rect 652 3928 692 3968
rect 81868 3928 81908 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 652 3592 692 3632
rect 16204 3592 16244 3632
rect 19276 3592 19316 3632
rect 25036 3592 25076 3632
rect 13324 3508 13364 3548
rect 20332 3508 20372 3548
rect 22156 3508 22196 3548
rect 28780 3508 28820 3548
rect 33292 3508 33332 3548
rect 46444 3508 46484 3548
rect 49036 3508 49076 3548
rect 52204 3508 52244 3548
rect 54988 3508 55028 3548
rect 12940 3424 12980 3464
rect 13228 3424 13268 3464
rect 13804 3424 13844 3464
rect 14188 3424 14228 3464
rect 15052 3424 15092 3464
rect 16876 3424 16916 3464
rect 17260 3437 17300 3477
rect 18124 3424 18164 3464
rect 20428 3424 20468 3464
rect 20716 3424 20756 3464
rect 21772 3424 21812 3464
rect 22060 3424 22100 3464
rect 22636 3424 22676 3464
rect 23020 3424 23060 3464
rect 23884 3424 23924 3464
rect 28396 3424 28436 3464
rect 28684 3424 28724 3464
rect 30796 3424 30836 3464
rect 31180 3424 31220 3464
rect 33388 3424 33428 3464
rect 33676 3424 33716 3464
rect 33964 3424 34004 3464
rect 34348 3424 34388 3464
rect 34636 3424 34676 3464
rect 34924 3424 34964 3464
rect 35020 3424 35060 3464
rect 36652 3424 36692 3464
rect 37036 3424 37076 3464
rect 37228 3424 37268 3464
rect 37612 3424 37652 3464
rect 37804 3424 37844 3464
rect 38188 3424 38228 3464
rect 39244 3424 39284 3464
rect 39340 3424 39380 3464
rect 39628 3424 39668 3464
rect 42700 3424 42740 3464
rect 46060 3424 46100 3464
rect 46348 3424 46388 3464
rect 48652 3424 48692 3464
rect 48940 3424 48980 3464
rect 51820 3424 51860 3464
rect 52108 3424 52148 3464
rect 54604 3424 54644 3464
rect 54892 3424 54932 3464
rect 21292 3340 21332 3380
rect 30892 3340 30932 3380
rect 31084 3340 31124 3380
rect 32812 3340 32852 3380
rect 34060 3340 34100 3380
rect 34252 3340 34292 3380
rect 36748 3340 36788 3380
rect 36940 3340 36980 3380
rect 37324 3340 37364 3380
rect 37516 3340 37556 3380
rect 37900 3340 37940 3380
rect 38092 3340 38132 3380
rect 42412 3340 42452 3380
rect 44524 3340 44564 3380
rect 45196 3340 45236 3380
rect 13612 3256 13652 3296
rect 22444 3256 22484 3296
rect 30988 3256 31028 3296
rect 34156 3256 34196 3296
rect 36844 3256 36884 3296
rect 37420 3256 37460 3296
rect 37996 3256 38036 3296
rect 20044 3172 20084 3212
rect 21484 3172 21524 3212
rect 29068 3172 29108 3212
rect 32620 3172 32660 3212
rect 33004 3172 33044 3212
rect 35308 3172 35348 3212
rect 38956 3172 38996 3212
rect 42220 3172 42260 3212
rect 45004 3172 45044 3212
rect 46732 3172 46772 3212
rect 49324 3172 49364 3212
rect 52492 3172 52532 3212
rect 55276 3172 55316 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 16876 2836 16916 2876
rect 22540 2836 22580 2876
rect 23212 2836 23252 2876
rect 32044 2836 32084 2876
rect 35212 2836 35252 2876
rect 38188 2836 38228 2876
rect 41356 2836 41396 2876
rect 49132 2836 49172 2876
rect 52012 2836 52052 2876
rect 55180 2836 55220 2876
rect 57772 2836 57812 2876
rect 25804 2752 25844 2792
rect 31180 2752 31220 2792
rect 43084 2752 43124 2792
rect 23404 2668 23444 2708
rect 32236 2668 32276 2708
rect 43276 2668 43316 2708
rect 17164 2584 17204 2624
rect 17260 2584 17300 2624
rect 17548 2584 17588 2624
rect 20140 2584 20180 2624
rect 20524 2584 20564 2624
rect 21388 2584 21428 2624
rect 25132 2584 25172 2624
rect 25420 2584 25460 2624
rect 25996 2584 26036 2624
rect 26380 2584 26420 2624
rect 27244 2584 27284 2624
rect 28780 2584 28820 2624
rect 29164 2584 29204 2624
rect 30028 2584 30068 2624
rect 32812 2584 32852 2624
rect 33196 2584 33236 2624
rect 34060 2584 34100 2624
rect 35788 2584 35828 2624
rect 36172 2584 36212 2624
rect 37036 2584 37076 2624
rect 38956 2584 38996 2624
rect 39340 2584 39380 2624
rect 40204 2584 40244 2624
rect 42412 2584 42452 2624
rect 42700 2584 42740 2624
rect 42796 2584 42836 2624
rect 44428 2584 44468 2624
rect 45292 2584 45332 2624
rect 45676 2584 45716 2624
rect 46732 2584 46772 2624
rect 47116 2584 47156 2624
rect 47980 2584 48020 2624
rect 49612 2584 49652 2624
rect 49996 2584 50036 2624
rect 50860 2584 50900 2624
rect 52780 2584 52820 2624
rect 53164 2584 53204 2624
rect 54053 2584 54093 2624
rect 55372 2584 55412 2624
rect 55756 2584 55796 2624
rect 56620 2584 56660 2624
rect 79852 2584 79892 2624
rect 80716 2584 80756 2624
rect 25516 2500 25556 2540
rect 79468 2500 79508 2540
rect 652 2416 692 2456
rect 23212 2416 23252 2456
rect 28396 2416 28436 2456
rect 81868 2416 81908 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 26476 2080 26516 2120
rect 30124 2080 30164 2120
rect 34540 2080 34580 2120
rect 34828 2080 34868 2120
rect 40108 2080 40148 2120
rect 42124 2080 42164 2120
rect 44908 2080 44948 2120
rect 22540 1996 22580 2036
rect 23500 1996 23540 2036
rect 31660 1996 31700 2036
rect 41644 1996 41684 2036
rect 19756 1912 19796 1952
rect 20620 1912 20660 1952
rect 21004 1912 21044 1952
rect 22156 1912 22196 1952
rect 22444 1912 22484 1952
rect 23116 1912 23156 1952
rect 23404 1912 23444 1952
rect 24076 1912 24116 1952
rect 24460 1912 24500 1952
rect 25324 1912 25364 1952
rect 26860 1912 26900 1952
rect 27148 1912 27188 1952
rect 27244 1912 27284 1952
rect 27724 1912 27764 1952
rect 28108 1912 28148 1952
rect 28972 1912 29012 1952
rect 31276 1912 31316 1952
rect 31564 1912 31604 1952
rect 32140 1912 32180 1952
rect 32524 1912 32564 1952
rect 33388 1912 33428 1952
rect 35980 1912 36020 1952
rect 36844 1912 36884 1952
rect 37228 1912 37268 1952
rect 37708 1912 37748 1952
rect 38092 1912 38132 1952
rect 38956 1912 38996 1952
rect 41260 1912 41300 1952
rect 41548 1912 41588 1952
rect 43276 1912 43316 1952
rect 44140 1912 44180 1952
rect 44524 1912 44564 1952
rect 46060 1912 46100 1952
rect 46924 1912 46964 1952
rect 47308 1912 47348 1952
rect 48652 1912 48692 1952
rect 49516 1912 49556 1952
rect 49900 1912 49940 1952
rect 51244 1912 51284 1952
rect 52108 1912 52148 1952
rect 52492 1912 52532 1952
rect 53836 1912 53876 1952
rect 54700 1912 54740 1952
rect 55084 1912 55124 1952
rect 72748 1912 72788 1952
rect 74092 1912 74132 1952
rect 78604 1912 78644 1952
rect 78892 1912 78932 1952
rect 78988 1912 79028 1952
rect 79468 1912 79508 1952
rect 79852 1912 79892 1952
rect 80716 1912 80756 1952
rect 23788 1744 23828 1784
rect 27532 1744 27572 1784
rect 31948 1744 31988 1784
rect 41932 1744 41972 1784
rect 79276 1744 79316 1784
rect 18604 1660 18644 1700
rect 22828 1660 22868 1700
rect 44908 1660 44948 1700
rect 47500 1660 47540 1700
rect 50092 1660 50132 1700
rect 52684 1660 52724 1700
rect 81868 1660 81908 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 20332 1324 20372 1364
rect 25036 1324 25076 1364
rect 32716 1324 32756 1364
rect 35404 1324 35444 1364
rect 37612 1324 37652 1364
rect 42892 1324 42932 1364
rect 45100 1324 45140 1364
rect 47596 1324 47636 1364
rect 50284 1324 50324 1364
rect 52780 1324 52820 1364
rect 79564 1324 79604 1364
rect 30124 1240 30164 1280
rect 40300 1240 40340 1280
rect 19660 1072 19700 1112
rect 19948 1072 19988 1112
rect 20044 1072 20084 1112
rect 22636 1072 22676 1112
rect 23020 1072 23060 1112
rect 23884 1072 23924 1112
rect 29452 1072 29492 1112
rect 29740 1072 29780 1112
rect 29836 1072 29876 1112
rect 30316 1072 30356 1112
rect 30700 1072 30740 1112
rect 31564 1072 31604 1112
rect 35692 1072 35732 1112
rect 35788 1072 35828 1112
rect 36076 1072 36116 1112
rect 37900 1072 37940 1112
rect 37996 1072 38036 1112
rect 38284 1072 38324 1112
rect 39628 1072 39668 1112
rect 39916 1072 39956 1112
rect 40012 1072 40052 1112
rect 40492 1072 40532 1112
rect 40876 1072 40916 1112
rect 41740 1072 41780 1112
rect 44428 1072 44468 1112
rect 44716 1072 44756 1112
rect 44812 1072 44852 1112
rect 46924 1072 46964 1112
rect 47212 1072 47252 1112
rect 49612 1072 49652 1112
rect 49900 1072 49940 1112
rect 49996 1072 50036 1112
rect 52108 1072 52148 1112
rect 52396 1072 52436 1112
rect 52492 1072 52532 1112
rect 79948 1072 79988 1112
rect 80236 1072 80276 1112
rect 47308 988 47348 1028
rect 79852 988 79892 1028
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 652 38156 692 38165
rect 652 37577 692 38116
rect 844 37988 884 37997
rect 651 37568 693 37577
rect 651 37528 652 37568
rect 692 37528 693 37568
rect 651 37519 693 37528
rect 267 35888 309 35897
rect 267 35848 268 35888
rect 308 35848 309 35888
rect 267 35839 309 35848
rect 268 5573 308 35839
rect 844 32117 884 37948
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 5739 36728 5781 36737
rect 5739 36688 5740 36728
rect 5780 36688 5781 36728
rect 5739 36679 5781 36688
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 5547 33872 5589 33881
rect 5547 33832 5548 33872
rect 5588 33832 5589 33872
rect 5547 33823 5589 33832
rect 3531 33704 3573 33713
rect 3531 33664 3532 33704
rect 3572 33664 3573 33704
rect 3531 33655 3573 33664
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 1707 33200 1749 33209
rect 1707 33160 1708 33200
rect 1748 33160 1749 33200
rect 1707 33151 1749 33160
rect 843 32108 885 32117
rect 843 32068 844 32108
rect 884 32068 885 32108
rect 843 32059 885 32068
rect 1419 31940 1461 31949
rect 1419 31900 1420 31940
rect 1460 31900 1461 31940
rect 1419 31891 1461 31900
rect 1324 31436 1364 31445
rect 1420 31436 1460 31891
rect 1516 31604 1556 31613
rect 1708 31604 1748 33151
rect 1899 32108 1941 32117
rect 1899 32068 1900 32108
rect 1940 32068 1941 32108
rect 1899 32059 1941 32068
rect 1900 31974 1940 32059
rect 2091 31940 2133 31949
rect 2091 31900 2092 31940
rect 2132 31900 2133 31940
rect 2091 31891 2133 31900
rect 2955 31940 2997 31949
rect 2955 31900 2956 31940
rect 2996 31900 2997 31940
rect 2955 31891 2997 31900
rect 2092 31806 2132 31891
rect 1556 31564 1748 31604
rect 1516 31555 1556 31564
rect 1364 31396 1460 31436
rect 1611 31436 1653 31445
rect 1611 31396 1612 31436
rect 1652 31396 1653 31436
rect 1324 31387 1364 31396
rect 1611 31387 1653 31396
rect 1708 31436 1748 31564
rect 1900 31520 1940 31531
rect 1900 31445 1940 31480
rect 1708 31387 1748 31396
rect 1899 31436 1941 31445
rect 1899 31396 1900 31436
rect 1940 31396 1941 31436
rect 1899 31387 1941 31396
rect 2763 31436 2805 31445
rect 2763 31396 2764 31436
rect 2804 31396 2805 31436
rect 2763 31387 2805 31396
rect 1515 30764 1557 30773
rect 1515 30724 1516 30764
rect 1556 30724 1557 30764
rect 1515 30715 1557 30724
rect 1228 30680 1268 30689
rect 1131 30260 1173 30269
rect 1131 30220 1132 30260
rect 1172 30220 1173 30260
rect 1131 30211 1173 30220
rect 939 29756 981 29765
rect 939 29716 940 29756
rect 980 29716 981 29756
rect 939 29707 981 29716
rect 747 28916 789 28925
rect 747 28876 748 28916
rect 788 28876 789 28916
rect 747 28867 789 28876
rect 748 28328 788 28867
rect 748 28279 788 28288
rect 651 26228 693 26237
rect 651 26188 652 26228
rect 692 26188 693 26228
rect 651 26179 693 26188
rect 652 26094 692 26179
rect 652 25388 692 25397
rect 652 24977 692 25348
rect 844 25136 884 25145
rect 748 25096 844 25136
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 748 24716 788 25096
rect 844 25087 884 25096
rect 844 24800 884 24809
rect 940 24800 980 29707
rect 1132 28328 1172 30211
rect 1228 30017 1268 30640
rect 1227 30008 1269 30017
rect 1227 29968 1228 30008
rect 1268 29968 1269 30008
rect 1227 29959 1269 29968
rect 1228 29840 1268 29849
rect 1228 29177 1268 29800
rect 1516 29840 1556 30715
rect 1612 30680 1652 31387
rect 2764 31352 2804 31387
rect 2764 31301 2804 31312
rect 1612 30269 1652 30640
rect 2380 31268 2420 31277
rect 1611 30260 1653 30269
rect 1611 30220 1612 30260
rect 1652 30220 1653 30260
rect 1611 30211 1653 30220
rect 1900 30092 1940 30101
rect 2380 30092 2420 31228
rect 2475 30932 2517 30941
rect 2475 30892 2476 30932
rect 2516 30892 2517 30932
rect 2475 30883 2517 30892
rect 2476 30680 2516 30883
rect 2476 30631 2516 30640
rect 1940 30052 2420 30092
rect 1900 30043 1940 30052
rect 2091 29924 2133 29933
rect 2956 29924 2996 31891
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 2091 29884 2092 29924
rect 2132 29884 2133 29924
rect 2091 29875 2133 29884
rect 2860 29884 2996 29924
rect 1516 29791 1556 29800
rect 1803 29840 1845 29849
rect 1803 29800 1804 29840
rect 1844 29800 1845 29840
rect 1803 29791 1845 29800
rect 1611 29756 1653 29765
rect 1611 29716 1612 29756
rect 1652 29716 1653 29756
rect 1611 29707 1653 29716
rect 1612 29622 1652 29707
rect 1227 29168 1269 29177
rect 1227 29128 1228 29168
rect 1268 29128 1269 29168
rect 1227 29119 1269 29128
rect 1419 29168 1461 29177
rect 1419 29128 1420 29168
rect 1460 29128 1461 29168
rect 1419 29119 1461 29128
rect 1516 29168 1556 29177
rect 1708 29168 1748 29177
rect 1804 29168 1844 29791
rect 2092 29790 2132 29875
rect 2188 29840 2228 29849
rect 2380 29840 2420 29849
rect 2228 29800 2380 29840
rect 2188 29791 2228 29800
rect 2380 29791 2420 29800
rect 2476 29840 2516 29849
rect 2091 29336 2133 29345
rect 2091 29296 2092 29336
rect 2132 29296 2133 29336
rect 2091 29287 2133 29296
rect 1556 29128 1652 29168
rect 1516 29119 1556 29128
rect 1036 26900 1076 26909
rect 1132 26900 1172 28288
rect 1420 27497 1460 29119
rect 1612 29009 1652 29128
rect 1748 29128 1844 29168
rect 1708 29119 1748 29128
rect 1611 29000 1653 29009
rect 1611 28960 1612 29000
rect 1652 28960 1653 29000
rect 1611 28951 1653 28960
rect 1515 28916 1557 28925
rect 1515 28876 1516 28916
rect 1556 28876 1557 28916
rect 1515 28867 1557 28876
rect 1516 28782 1556 28867
rect 1804 27740 1844 29128
rect 1900 29168 1940 29177
rect 2092 29168 2132 29287
rect 2188 29177 2228 29262
rect 2476 29261 2516 29800
rect 2571 29840 2613 29849
rect 2571 29800 2572 29840
rect 2612 29800 2613 29840
rect 2571 29791 2613 29800
rect 2668 29840 2708 29851
rect 2572 29706 2612 29791
rect 2668 29765 2708 29800
rect 2667 29756 2709 29765
rect 2667 29716 2668 29756
rect 2708 29716 2709 29756
rect 2667 29707 2709 29716
rect 2860 29504 2900 29884
rect 2955 29756 2997 29765
rect 2955 29716 2956 29756
rect 2996 29716 2997 29756
rect 2955 29707 2997 29716
rect 3436 29756 3476 29765
rect 2572 29464 2900 29504
rect 2475 29252 2517 29261
rect 2475 29212 2476 29252
rect 2516 29212 2517 29252
rect 2475 29203 2517 29212
rect 1940 29128 2036 29168
rect 1900 29119 1940 29128
rect 1899 29000 1941 29009
rect 1899 28960 1900 29000
rect 1940 28960 1941 29000
rect 1899 28951 1941 28960
rect 1900 28866 1940 28951
rect 1996 28757 2036 29128
rect 1995 28748 2037 28757
rect 1995 28708 1996 28748
rect 2036 28708 2037 28748
rect 1995 28699 2037 28708
rect 2092 28496 2132 29128
rect 2187 29168 2229 29177
rect 2187 29128 2188 29168
rect 2228 29128 2229 29168
rect 2187 29119 2229 29128
rect 2379 28748 2421 28757
rect 2379 28708 2380 28748
rect 2420 28708 2421 28748
rect 2379 28699 2421 28708
rect 1804 27691 1844 27700
rect 1900 28456 2132 28496
rect 1900 27824 1940 28456
rect 1996 28328 2036 28337
rect 2036 28288 2228 28328
rect 1996 28279 2036 28288
rect 2092 27824 2132 27833
rect 1900 27784 2092 27824
rect 1419 27488 1461 27497
rect 1419 27448 1420 27488
rect 1460 27448 1461 27488
rect 1419 27439 1461 27448
rect 1076 26860 1172 26900
rect 1036 26851 1076 26860
rect 1035 26144 1077 26153
rect 1035 26104 1036 26144
rect 1076 26104 1077 26144
rect 1035 26095 1077 26104
rect 1036 26010 1076 26095
rect 884 24760 980 24800
rect 844 24751 884 24760
rect 1132 24716 1172 26860
rect 1420 26816 1460 27439
rect 1900 26825 1940 27784
rect 2092 27775 2132 27784
rect 1996 27656 2036 27665
rect 1996 27497 2036 27616
rect 2091 27656 2133 27665
rect 2091 27616 2092 27656
rect 2132 27616 2133 27656
rect 2091 27607 2133 27616
rect 2092 27522 2132 27607
rect 1995 27488 2037 27497
rect 1995 27448 1996 27488
rect 2036 27448 2037 27488
rect 1995 27439 2037 27448
rect 1996 27329 2036 27439
rect 1995 27320 2037 27329
rect 1995 27280 1996 27320
rect 2036 27280 2037 27320
rect 1995 27271 2037 27280
rect 1228 26648 1268 26657
rect 1228 26153 1268 26608
rect 1227 26144 1269 26153
rect 1227 26104 1228 26144
rect 1268 26104 1269 26144
rect 1227 26095 1269 26104
rect 460 24676 788 24716
rect 940 24676 1172 24716
rect 460 15569 500 24676
rect 652 24548 692 24557
rect 652 23297 692 24508
rect 844 23792 884 23803
rect 844 23717 884 23752
rect 843 23708 885 23717
rect 843 23668 844 23708
rect 884 23668 885 23708
rect 843 23659 885 23668
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 651 23120 693 23129
rect 651 23080 652 23120
rect 692 23080 693 23120
rect 940 23120 980 24676
rect 1420 24557 1460 26776
rect 1515 26816 1557 26825
rect 1515 26776 1516 26816
rect 1556 26776 1557 26816
rect 1515 26767 1557 26776
rect 1708 26816 1748 26825
rect 1516 25304 1556 26767
rect 1612 26648 1652 26657
rect 1612 26237 1652 26608
rect 1611 26228 1653 26237
rect 1611 26188 1612 26228
rect 1652 26188 1653 26228
rect 1611 26179 1653 26188
rect 1708 25556 1748 26776
rect 1899 26816 1941 26825
rect 1899 26776 1900 26816
rect 1940 26776 1941 26816
rect 1899 26767 1941 26776
rect 1900 26144 1940 26153
rect 2188 26144 2228 28288
rect 2380 27665 2420 28699
rect 2379 27656 2421 27665
rect 2379 27616 2380 27656
rect 2420 27616 2421 27656
rect 2379 27607 2421 27616
rect 2380 26816 2420 27607
rect 2572 27380 2612 29464
rect 2668 29336 2708 29347
rect 2956 29345 2996 29707
rect 2668 29261 2708 29296
rect 2763 29336 2805 29345
rect 2763 29296 2764 29336
rect 2804 29296 2805 29336
rect 2763 29287 2805 29296
rect 2955 29336 2997 29345
rect 2955 29296 2956 29336
rect 2996 29296 2997 29336
rect 3436 29336 3476 29716
rect 3532 29513 3572 33655
rect 5356 32780 5396 32789
rect 5164 32740 5356 32780
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4972 31604 5012 31613
rect 5164 31604 5204 32740
rect 5356 32731 5396 32740
rect 5259 32444 5301 32453
rect 5259 32404 5260 32444
rect 5300 32404 5301 32444
rect 5259 32395 5301 32404
rect 5012 31564 5204 31604
rect 4972 31555 5012 31564
rect 3819 31436 3861 31445
rect 3819 31396 3820 31436
rect 3860 31396 3861 31436
rect 3819 31387 3861 31396
rect 3627 31352 3669 31361
rect 3627 31312 3628 31352
rect 3668 31312 3669 31352
rect 3627 31303 3669 31312
rect 3628 30941 3668 31303
rect 3627 30932 3669 30941
rect 3627 30892 3628 30932
rect 3668 30892 3669 30932
rect 3627 30883 3669 30892
rect 3628 30428 3668 30437
rect 3668 30388 3764 30428
rect 3628 30379 3668 30388
rect 3531 29504 3573 29513
rect 3531 29464 3532 29504
rect 3572 29464 3573 29504
rect 3531 29455 3573 29464
rect 3724 29345 3764 30388
rect 3820 30269 3860 31387
rect 4875 31352 4917 31361
rect 4875 31312 4876 31352
rect 4916 31312 4917 31352
rect 4875 31303 4917 31312
rect 5260 31352 5300 32395
rect 5260 31303 5300 31312
rect 5356 31348 5396 31357
rect 4779 31184 4821 31193
rect 4779 31144 4780 31184
rect 4820 31144 4821 31184
rect 4779 31135 4821 31144
rect 4780 31050 4820 31135
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 4876 30848 4916 31303
rect 4684 30808 4916 30848
rect 3819 30260 3861 30269
rect 3819 30220 3820 30260
rect 3860 30220 3861 30260
rect 3819 30211 3861 30220
rect 3820 29840 3860 30211
rect 3820 29791 3860 29800
rect 4684 29840 4724 30808
rect 4684 29791 4724 29800
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3532 29336 3572 29345
rect 3436 29296 3532 29336
rect 2955 29287 2997 29296
rect 3532 29287 3572 29296
rect 3723 29336 3765 29345
rect 3820 29336 3860 29345
rect 3723 29296 3724 29336
rect 3764 29296 3820 29336
rect 3723 29287 3765 29296
rect 3820 29287 3860 29296
rect 2667 29252 2709 29261
rect 2667 29212 2668 29252
rect 2708 29212 2709 29252
rect 2667 29203 2709 29212
rect 2764 29202 2804 29287
rect 2860 29252 2900 29261
rect 2860 28757 2900 29212
rect 2956 29168 2996 29287
rect 3724 29202 3764 29287
rect 2956 29119 2996 29128
rect 3051 29168 3093 29177
rect 3051 29128 3052 29168
rect 3092 29128 3093 29168
rect 3051 29119 3093 29128
rect 3339 29168 3381 29177
rect 3339 29128 3340 29168
rect 3380 29128 3381 29168
rect 3339 29119 3381 29128
rect 3436 29168 3476 29177
rect 3052 29034 3092 29119
rect 3340 29034 3380 29119
rect 3436 28925 3476 29128
rect 3628 29168 3668 29177
rect 3435 28916 3477 28925
rect 3435 28876 3436 28916
rect 3476 28876 3477 28916
rect 3435 28867 3477 28876
rect 2859 28748 2901 28757
rect 3112 28748 3480 28757
rect 2859 28708 2860 28748
rect 2900 28708 2996 28748
rect 2859 28699 2901 28708
rect 2860 28614 2900 28699
rect 2956 28580 2996 28708
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3147 28580 3189 28589
rect 2956 28540 3148 28580
rect 3188 28540 3189 28580
rect 3147 28531 3189 28540
rect 3531 28580 3573 28589
rect 3531 28540 3532 28580
rect 3572 28540 3573 28580
rect 3531 28531 3573 28540
rect 3148 28446 3188 28531
rect 3436 28328 3476 28337
rect 2764 28288 3436 28328
rect 2764 27824 2804 28288
rect 3436 28279 3476 28288
rect 3532 28328 3572 28531
rect 3628 28505 3668 29128
rect 3915 29168 3957 29177
rect 3915 29128 3916 29168
rect 3956 29128 3957 29168
rect 3915 29119 3957 29128
rect 4491 29168 4533 29177
rect 4491 29128 4492 29168
rect 4532 29128 4533 29168
rect 4491 29119 4533 29128
rect 4588 29168 4628 29177
rect 4780 29168 4820 29177
rect 4628 29128 4780 29168
rect 4588 29119 4628 29128
rect 4780 29119 4820 29128
rect 3916 29034 3956 29119
rect 4108 28916 4148 28925
rect 3724 28876 4108 28916
rect 3627 28496 3669 28505
rect 3627 28456 3628 28496
rect 3668 28456 3669 28496
rect 3627 28447 3669 28456
rect 3532 28279 3572 28288
rect 3628 28328 3668 28337
rect 2764 27380 2804 27784
rect 2859 27656 2901 27665
rect 3628 27656 3668 28288
rect 2859 27616 2860 27656
rect 2900 27616 2901 27656
rect 2859 27607 2901 27616
rect 3532 27616 3668 27656
rect 3724 28328 3764 28876
rect 4108 28867 4148 28876
rect 4395 28916 4437 28925
rect 4395 28876 4396 28916
rect 4436 28876 4437 28916
rect 4395 28867 4437 28876
rect 3915 28496 3957 28505
rect 3915 28456 3916 28496
rect 3956 28456 4148 28496
rect 3915 28447 3957 28456
rect 3916 28362 3956 28447
rect 2860 27522 2900 27607
rect 3052 27497 3092 27582
rect 3435 27572 3477 27581
rect 3435 27532 3436 27572
rect 3476 27532 3477 27572
rect 3435 27523 3477 27532
rect 3051 27488 3093 27497
rect 3051 27448 3052 27488
rect 3092 27448 3093 27488
rect 3051 27439 3093 27448
rect 3436 27438 3476 27523
rect 3532 27413 3572 27616
rect 3627 27488 3669 27497
rect 3627 27448 3628 27488
rect 3668 27448 3669 27488
rect 3627 27439 3669 27448
rect 3531 27404 3573 27413
rect 2572 27340 2708 27380
rect 2764 27340 2996 27380
rect 3531 27364 3532 27404
rect 3572 27364 3573 27404
rect 3531 27355 3573 27364
rect 2668 26984 2708 27340
rect 2668 26944 2804 26984
rect 2380 26767 2420 26776
rect 2667 26816 2709 26825
rect 2667 26776 2668 26816
rect 2708 26776 2709 26816
rect 2667 26767 2709 26776
rect 2668 26682 2708 26767
rect 2572 26648 2612 26657
rect 2572 26153 2612 26608
rect 2764 26480 2804 26944
rect 2956 26816 2996 27340
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3532 27068 3572 27355
rect 3436 27028 3572 27068
rect 3051 26816 3093 26825
rect 2956 26776 3052 26816
rect 3092 26776 3093 26816
rect 3051 26767 3093 26776
rect 3340 26816 3380 26827
rect 2668 26440 2804 26480
rect 1940 26104 2228 26144
rect 1900 26095 1940 26104
rect 1995 25976 2037 25985
rect 1995 25936 1996 25976
rect 2036 25936 2037 25976
rect 1995 25927 2037 25936
rect 1708 25507 1748 25516
rect 1708 25304 1748 25313
rect 1516 25264 1708 25304
rect 1708 25255 1748 25264
rect 1900 25304 1940 25313
rect 1900 24557 1940 25264
rect 1996 25304 2036 25927
rect 2188 25313 2228 26104
rect 2571 26144 2613 26153
rect 2571 26104 2572 26144
rect 2612 26104 2613 26144
rect 2571 26095 2613 26104
rect 2187 25304 2229 25313
rect 2036 25264 2132 25304
rect 1996 25255 2036 25264
rect 2092 24632 2132 25264
rect 2187 25264 2188 25304
rect 2228 25264 2229 25304
rect 2187 25255 2229 25264
rect 2188 24632 2228 24641
rect 2092 24592 2188 24632
rect 2188 24583 2228 24592
rect 1036 24548 1076 24557
rect 1036 24137 1076 24508
rect 1131 24548 1173 24557
rect 1131 24508 1132 24548
rect 1172 24508 1173 24548
rect 1131 24499 1173 24508
rect 1419 24548 1461 24557
rect 1419 24508 1420 24548
rect 1460 24508 1461 24548
rect 1419 24499 1461 24508
rect 1899 24548 1941 24557
rect 1899 24508 1900 24548
rect 1940 24508 1941 24548
rect 1899 24499 1941 24508
rect 1035 24128 1077 24137
rect 1035 24088 1036 24128
rect 1076 24088 1077 24128
rect 1035 24079 1077 24088
rect 1132 23876 1172 24499
rect 1228 24380 1268 24389
rect 2092 24380 2132 24389
rect 1268 24340 1460 24380
rect 1228 24331 1268 24340
rect 1036 23836 1172 23876
rect 1324 23960 1364 23969
rect 1036 23792 1076 23836
rect 1036 23743 1076 23752
rect 1132 23785 1172 23794
rect 1132 23633 1172 23745
rect 1227 23708 1269 23717
rect 1227 23668 1228 23708
rect 1268 23668 1269 23708
rect 1227 23659 1269 23668
rect 1131 23624 1173 23633
rect 1131 23584 1132 23624
rect 1172 23584 1173 23624
rect 1131 23575 1173 23584
rect 1036 23120 1076 23129
rect 940 23080 1036 23120
rect 651 23071 693 23080
rect 1036 23071 1076 23080
rect 652 22986 692 23071
rect 1228 22532 1268 23659
rect 1324 23129 1364 23920
rect 1323 23120 1365 23129
rect 1323 23080 1324 23120
rect 1364 23080 1365 23120
rect 1323 23071 1365 23080
rect 1228 22483 1268 22492
rect 1035 22364 1077 22373
rect 1035 22324 1036 22364
rect 1076 22324 1077 22364
rect 1035 22315 1077 22324
rect 1036 22230 1076 22315
rect 652 22112 692 22121
rect 652 21617 692 22072
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 1420 20852 1460 24340
rect 1804 24340 2092 24380
rect 1611 23792 1653 23801
rect 1611 23752 1612 23792
rect 1652 23752 1653 23792
rect 1611 23743 1653 23752
rect 1708 23792 1748 23803
rect 1612 23633 1652 23743
rect 1708 23717 1748 23752
rect 1707 23708 1749 23717
rect 1707 23668 1708 23708
rect 1748 23668 1749 23708
rect 1707 23659 1749 23668
rect 1611 23624 1653 23633
rect 1611 23584 1612 23624
rect 1652 23584 1653 23624
rect 1611 23575 1653 23584
rect 1804 23620 1844 24340
rect 2092 24331 2132 24340
rect 1995 23792 2037 23801
rect 1995 23752 1996 23792
rect 2036 23752 2037 23792
rect 1995 23743 2037 23752
rect 2092 23792 2132 23803
rect 1804 23571 1844 23580
rect 1996 23297 2036 23743
rect 2092 23717 2132 23752
rect 2091 23708 2133 23717
rect 2091 23668 2092 23708
rect 2132 23668 2133 23708
rect 2091 23659 2133 23668
rect 2284 23624 2324 23633
rect 1995 23288 2037 23297
rect 1995 23248 1996 23288
rect 2036 23248 2037 23288
rect 1995 23239 2037 23248
rect 2284 23213 2324 23584
rect 2283 23204 2325 23213
rect 2283 23164 2284 23204
rect 2324 23164 2325 23204
rect 2283 23155 2325 23164
rect 1899 23120 1941 23129
rect 1899 23080 1900 23120
rect 1940 23080 2036 23120
rect 1899 23071 1941 23080
rect 1900 22986 1940 23071
rect 1515 21524 1557 21533
rect 1515 21484 1516 21524
rect 1556 21484 1557 21524
rect 1515 21475 1557 21484
rect 1324 20812 1460 20852
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 652 20600 692 20719
rect 652 20551 692 20560
rect 652 20264 692 20273
rect 652 19937 692 20224
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18954 692 19039
rect 1227 18668 1269 18677
rect 1227 18628 1228 18668
rect 1268 18628 1269 18668
rect 1227 18619 1269 18628
rect 843 18584 885 18593
rect 843 18544 844 18584
rect 884 18544 885 18584
rect 843 18535 885 18544
rect 1228 18584 1268 18619
rect 844 18450 884 18535
rect 1228 18533 1268 18544
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17576 692 18199
rect 1227 17744 1269 17753
rect 1227 17704 1228 17744
rect 1268 17704 1269 17744
rect 1227 17695 1269 17704
rect 652 17527 692 17536
rect 1228 17576 1268 17695
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 17240 692 17359
rect 652 17191 692 17200
rect 1036 17240 1076 17249
rect 1036 16577 1076 17200
rect 1035 16568 1077 16577
rect 1035 16528 1036 16568
rect 1076 16528 1077 16568
rect 1035 16519 1077 16528
rect 1228 16316 1268 17536
rect 652 16064 692 16073
rect 652 15737 692 16024
rect 1228 15905 1268 16276
rect 1227 15896 1269 15905
rect 1227 15856 1228 15896
rect 1268 15856 1269 15896
rect 1227 15847 1269 15856
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 459 15560 501 15569
rect 459 15520 460 15560
rect 500 15520 501 15560
rect 1324 15560 1364 20812
rect 1420 17828 1460 17837
rect 1420 17669 1460 17788
rect 1419 17660 1461 17669
rect 1419 17620 1420 17660
rect 1460 17620 1461 17660
rect 1419 17611 1461 17620
rect 1516 16316 1556 21475
rect 1900 19088 1940 19097
rect 1804 19048 1900 19088
rect 1611 18584 1653 18593
rect 1611 18544 1612 18584
rect 1652 18544 1653 18584
rect 1611 18535 1653 18544
rect 1612 17996 1652 18535
rect 1612 17947 1652 17956
rect 1804 17669 1844 19048
rect 1900 19039 1940 19048
rect 1996 18584 2036 23080
rect 2091 20936 2133 20945
rect 2091 20896 2092 20936
rect 2132 20896 2133 20936
rect 2091 20887 2133 20896
rect 2092 19340 2132 20887
rect 2475 20684 2517 20693
rect 2475 20644 2476 20684
rect 2516 20644 2517 20684
rect 2475 20635 2517 20644
rect 2476 19928 2516 20635
rect 2476 19879 2516 19888
rect 2092 19291 2132 19300
rect 2092 18584 2132 18593
rect 1996 18544 2092 18584
rect 2092 18535 2132 18544
rect 1899 18332 1941 18341
rect 1899 18292 1900 18332
rect 1940 18292 1941 18332
rect 1899 18283 1941 18292
rect 1900 17744 1940 18283
rect 2668 17828 2708 26440
rect 3052 26312 3092 26767
rect 3340 26741 3380 26776
rect 3436 26816 3476 27028
rect 3628 26825 3668 27439
rect 3436 26767 3476 26776
rect 3532 26816 3572 26825
rect 3339 26732 3381 26741
rect 3339 26692 3340 26732
rect 3380 26692 3381 26732
rect 3339 26683 3381 26692
rect 3532 26564 3572 26776
rect 3627 26816 3669 26825
rect 3627 26776 3628 26816
rect 3668 26776 3669 26816
rect 3627 26767 3669 26776
rect 3628 26682 3668 26767
rect 3724 26573 3764 28288
rect 4108 28328 4148 28456
rect 4108 28279 4148 28288
rect 4300 28328 4340 28337
rect 4300 28169 4340 28288
rect 4107 28160 4149 28169
rect 4107 28120 4108 28160
rect 4148 28120 4149 28160
rect 4107 28111 4149 28120
rect 4204 28160 4244 28169
rect 4108 27329 4148 28111
rect 4204 27413 4244 28120
rect 4299 28160 4341 28169
rect 4299 28120 4300 28160
rect 4340 28120 4341 28160
rect 4396 28160 4436 28867
rect 4492 28328 4532 29119
rect 5068 28916 5108 28925
rect 4588 28328 4628 28337
rect 4492 28288 4588 28328
rect 4588 28279 4628 28288
rect 4780 28328 4820 28337
rect 4492 28160 4532 28169
rect 4396 28120 4492 28160
rect 4299 28111 4341 28120
rect 4492 28111 4532 28120
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 4587 27656 4629 27665
rect 4587 27616 4588 27656
rect 4628 27616 4629 27656
rect 4587 27607 4629 27616
rect 4588 27522 4628 27607
rect 4203 27404 4245 27413
rect 4203 27364 4204 27404
rect 4244 27364 4245 27404
rect 4203 27355 4245 27364
rect 4587 27404 4629 27413
rect 4587 27364 4588 27404
rect 4628 27364 4629 27404
rect 4587 27355 4629 27364
rect 4107 27320 4149 27329
rect 4107 27280 4108 27320
rect 4148 27280 4149 27320
rect 4107 27271 4149 27280
rect 4299 27320 4341 27329
rect 4299 27280 4300 27320
rect 4340 27280 4341 27320
rect 4299 27271 4341 27280
rect 4108 26984 4148 26993
rect 3916 26944 4108 26984
rect 3819 26648 3861 26657
rect 3819 26608 3820 26648
rect 3860 26608 3861 26648
rect 3819 26599 3861 26608
rect 3723 26564 3765 26573
rect 3532 26524 3724 26564
rect 3764 26524 3765 26564
rect 3340 26312 3380 26321
rect 3052 26263 3092 26272
rect 3244 26272 3340 26312
rect 3244 26144 3284 26272
rect 3340 26263 3380 26272
rect 2956 26104 3284 26144
rect 3436 26228 3476 26237
rect 2956 25145 2996 26104
rect 3340 25985 3380 26070
rect 3436 26069 3476 26188
rect 3531 26144 3573 26153
rect 3531 26104 3532 26144
rect 3572 26104 3573 26144
rect 3531 26095 3573 26104
rect 3628 26144 3668 26524
rect 3723 26515 3765 26524
rect 3724 26430 3764 26515
rect 3820 26514 3860 26599
rect 3916 26396 3956 26944
rect 4108 26935 4148 26944
rect 4011 26816 4053 26825
rect 4011 26776 4012 26816
rect 4052 26776 4053 26816
rect 4011 26767 4053 26776
rect 4108 26816 4148 26825
rect 4012 26682 4052 26767
rect 4108 26573 4148 26776
rect 4300 26816 4340 27271
rect 4300 26741 4340 26776
rect 4492 26816 4532 26825
rect 4588 26816 4628 27355
rect 4684 27077 4724 27162
rect 4683 27068 4725 27077
rect 4683 27028 4684 27068
rect 4724 27028 4725 27068
rect 4683 27019 4725 27028
rect 4684 26816 4724 26825
rect 4588 26776 4684 26816
rect 4299 26732 4341 26741
rect 4299 26692 4300 26732
rect 4340 26692 4341 26732
rect 4299 26683 4341 26692
rect 4492 26657 4532 26776
rect 4684 26767 4724 26776
rect 4203 26648 4245 26657
rect 4203 26608 4204 26648
rect 4244 26608 4245 26648
rect 4203 26599 4245 26608
rect 4491 26648 4533 26657
rect 4491 26608 4492 26648
rect 4532 26608 4533 26648
rect 4491 26599 4533 26608
rect 4107 26564 4149 26573
rect 4107 26524 4108 26564
rect 4148 26524 4149 26564
rect 4107 26515 4149 26524
rect 3820 26356 3956 26396
rect 3723 26228 3765 26237
rect 3723 26188 3724 26228
rect 3764 26188 3765 26228
rect 3723 26179 3765 26188
rect 3628 26095 3668 26104
rect 3435 26060 3477 26069
rect 3435 26020 3436 26060
rect 3476 26020 3477 26060
rect 3435 26011 3477 26020
rect 3532 26010 3572 26095
rect 3339 25976 3381 25985
rect 3339 25936 3340 25976
rect 3380 25936 3381 25976
rect 3339 25927 3381 25936
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3724 25304 3764 26179
rect 3820 26144 3860 26356
rect 4204 26312 4244 26599
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 4683 26312 4725 26321
rect 4204 26272 4340 26312
rect 3915 26228 3957 26237
rect 3915 26188 3916 26228
rect 3956 26188 3957 26228
rect 3915 26179 3957 26188
rect 3820 26095 3860 26104
rect 3916 26144 3956 26179
rect 3916 26093 3956 26104
rect 4108 26144 4148 26153
rect 4300 26144 4340 26272
rect 4683 26272 4684 26312
rect 4724 26272 4725 26312
rect 4683 26263 4725 26272
rect 4148 26104 4244 26144
rect 4108 26095 4148 26104
rect 3916 25976 3956 25985
rect 3820 25304 3860 25313
rect 3532 25264 3820 25304
rect 3436 25220 3476 25229
rect 2955 25136 2997 25145
rect 2955 25096 2956 25136
rect 2996 25096 2997 25136
rect 2955 25087 2997 25096
rect 3244 24716 3284 24725
rect 2956 24676 3244 24716
rect 2956 24212 2996 24676
rect 3244 24667 3284 24676
rect 3339 24632 3381 24641
rect 3339 24592 3340 24632
rect 3380 24592 3381 24632
rect 3339 24583 3381 24592
rect 3340 24498 3380 24583
rect 3436 24473 3476 25180
rect 3435 24464 3477 24473
rect 3435 24424 3436 24464
rect 3476 24424 3477 24464
rect 3435 24415 3477 24424
rect 2860 24172 2996 24212
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 2860 23834 2900 24172
rect 3112 24163 3480 24172
rect 2860 23785 2900 23794
rect 3244 23792 3284 23801
rect 3532 23792 3572 25264
rect 3820 25255 3860 25264
rect 3723 25136 3765 25145
rect 3723 25096 3724 25136
rect 3764 25096 3765 25136
rect 3723 25087 3765 25096
rect 3724 24632 3764 25087
rect 3916 24641 3956 25936
rect 4107 25892 4149 25901
rect 4107 25852 4108 25892
rect 4148 25852 4149 25892
rect 4107 25843 4149 25852
rect 4011 25304 4053 25313
rect 4011 25264 4012 25304
rect 4052 25264 4053 25304
rect 4011 25255 4053 25264
rect 3724 24557 3764 24592
rect 3915 24632 3957 24641
rect 3915 24592 3916 24632
rect 3956 24592 3957 24632
rect 3915 24583 3957 24592
rect 3723 24548 3765 24557
rect 3723 24508 3724 24548
rect 3764 24508 3765 24548
rect 3723 24499 3765 24508
rect 3916 24498 3956 24583
rect 3284 23752 3572 23792
rect 4012 23792 4052 25255
rect 4108 24632 4148 25843
rect 4204 24800 4244 26104
rect 4300 26095 4340 26104
rect 4491 26144 4533 26153
rect 4491 26104 4492 26144
rect 4532 26104 4533 26144
rect 4491 26095 4533 26104
rect 4684 26144 4724 26263
rect 4684 26095 4724 26104
rect 4299 25892 4341 25901
rect 4299 25852 4300 25892
rect 4340 25852 4341 25892
rect 4299 25843 4341 25852
rect 4300 25758 4340 25843
rect 4492 25145 4532 26095
rect 4683 25304 4725 25313
rect 4683 25264 4684 25304
rect 4724 25264 4725 25304
rect 4683 25255 4725 25264
rect 4684 25170 4724 25255
rect 4491 25136 4533 25145
rect 4491 25096 4492 25136
rect 4532 25096 4533 25136
rect 4491 25087 4533 25096
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 4300 24800 4340 24809
rect 4204 24760 4300 24800
rect 4300 24751 4340 24760
rect 4395 24800 4437 24809
rect 4395 24760 4396 24800
rect 4436 24760 4437 24800
rect 4395 24751 4437 24760
rect 4108 24583 4148 24592
rect 4396 24632 4436 24751
rect 4396 24583 4436 24592
rect 4107 24464 4149 24473
rect 4107 24424 4108 24464
rect 4148 24424 4149 24464
rect 4107 24415 4149 24424
rect 4108 24330 4148 24415
rect 4203 24380 4245 24389
rect 4203 24340 4204 24380
rect 4244 24340 4245 24380
rect 4203 24331 4245 24340
rect 4108 23792 4148 23801
rect 4012 23752 4108 23792
rect 3244 23743 3284 23752
rect 3051 23288 3093 23297
rect 3051 23248 3052 23288
rect 3092 23248 3093 23288
rect 3051 23239 3093 23248
rect 3052 23154 3092 23239
rect 3532 23060 3572 23752
rect 4108 23743 4148 23752
rect 4204 23060 4244 24331
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 4395 23288 4437 23297
rect 4395 23248 4396 23288
rect 4436 23248 4437 23288
rect 4395 23239 4437 23248
rect 4396 23154 4436 23239
rect 4587 23204 4629 23213
rect 4587 23164 4588 23204
rect 4628 23164 4629 23204
rect 4587 23155 4629 23164
rect 3532 23020 3860 23060
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 3820 22280 3860 23020
rect 3436 22196 3476 22205
rect 3476 22156 3764 22196
rect 3436 22147 3476 22156
rect 3531 21608 3573 21617
rect 3531 21568 3532 21608
rect 3572 21568 3573 21608
rect 3531 21559 3573 21568
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 3532 21020 3572 21559
rect 3724 21440 3764 22156
rect 3820 21617 3860 22240
rect 4108 23036 4244 23060
rect 4588 23045 4628 23155
rect 4683 23120 4725 23129
rect 4683 23080 4684 23120
rect 4724 23080 4725 23120
rect 4683 23071 4725 23080
rect 4108 23020 4204 23036
rect 3819 21608 3861 21617
rect 3819 21568 3820 21608
rect 3860 21568 3861 21608
rect 3819 21559 3861 21568
rect 4012 21440 4052 21449
rect 3724 21400 4012 21440
rect 4012 21391 4052 21400
rect 3148 20980 3860 21020
rect 3148 20768 3188 20980
rect 3148 20719 3188 20728
rect 2763 20684 2805 20693
rect 2763 20644 2764 20684
rect 2804 20644 2805 20684
rect 2763 20635 2805 20644
rect 2764 20550 2804 20635
rect 2859 20600 2901 20609
rect 2859 20560 2860 20600
rect 2900 20560 2901 20600
rect 2859 20551 2901 20560
rect 2860 20264 2900 20551
rect 2764 20224 2900 20264
rect 2764 20180 2804 20224
rect 2764 20131 2804 20140
rect 2860 20096 2900 20105
rect 2860 18341 2900 20056
rect 3147 20096 3189 20105
rect 3147 20056 3148 20096
rect 3188 20056 3189 20096
rect 3147 20047 3189 20056
rect 3436 20096 3476 20107
rect 3148 19962 3188 20047
rect 3436 20021 3476 20056
rect 3820 20096 3860 20980
rect 4108 20945 4148 23020
rect 4204 22877 4244 22996
rect 4587 23036 4629 23045
rect 4587 22996 4588 23036
rect 4628 22996 4629 23036
rect 4587 22987 4629 22996
rect 4588 22902 4628 22987
rect 4203 22868 4245 22877
rect 4203 22828 4204 22868
rect 4244 22828 4245 22868
rect 4203 22819 4245 22828
rect 4684 22280 4724 23071
rect 4780 23036 4820 28288
rect 4971 27656 5013 27665
rect 4971 27616 4972 27656
rect 5012 27616 5013 27656
rect 4971 27607 5013 27616
rect 4875 26144 4917 26153
rect 4875 26104 4876 26144
rect 4916 26104 4917 26144
rect 4875 26095 4917 26104
rect 4876 26010 4916 26095
rect 4875 25892 4917 25901
rect 4875 25852 4876 25892
rect 4916 25852 4917 25892
rect 4875 25843 4917 25852
rect 4876 25758 4916 25843
rect 4972 25313 5012 27607
rect 4971 25304 5013 25313
rect 4971 25264 4972 25304
rect 5012 25264 5013 25304
rect 4971 25255 5013 25264
rect 4971 24464 5013 24473
rect 4971 24424 4972 24464
rect 5012 24424 5013 24464
rect 4971 24415 5013 24424
rect 4780 22996 4916 23036
rect 4779 22868 4821 22877
rect 4779 22828 4780 22868
rect 4820 22828 4821 22868
rect 4779 22819 4821 22828
rect 4780 22734 4820 22819
rect 4204 22240 4684 22280
rect 4107 20936 4149 20945
rect 4107 20896 4108 20936
rect 4148 20896 4149 20936
rect 4107 20887 4149 20896
rect 4012 20768 4052 20777
rect 4204 20768 4244 22240
rect 4684 22231 4724 22240
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 4683 21776 4725 21785
rect 4683 21736 4684 21776
rect 4724 21736 4725 21776
rect 4683 21727 4725 21736
rect 4299 21692 4341 21701
rect 4299 21652 4300 21692
rect 4340 21652 4341 21692
rect 4299 21643 4341 21652
rect 4300 21558 4340 21643
rect 4395 21608 4437 21617
rect 4395 21568 4396 21608
rect 4436 21568 4437 21608
rect 4395 21559 4437 21568
rect 4684 21608 4724 21727
rect 4724 21568 4820 21608
rect 4684 21559 4724 21568
rect 4396 21474 4436 21559
rect 4052 20728 4244 20768
rect 4012 20719 4052 20728
rect 4204 20264 4244 20728
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4204 20224 4724 20264
rect 3435 20012 3477 20021
rect 3435 19972 3436 20012
rect 3476 19972 3477 20012
rect 3435 19963 3477 19972
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3820 18677 3860 20056
rect 4684 20096 4724 20224
rect 4780 20105 4820 21568
rect 4684 20047 4724 20056
rect 4779 20096 4821 20105
rect 4779 20056 4780 20096
rect 4820 20056 4821 20096
rect 4779 20047 4821 20056
rect 4299 20012 4341 20021
rect 4299 19972 4300 20012
rect 4340 19972 4341 20012
rect 4299 19963 4341 19972
rect 4300 19508 4340 19963
rect 4587 19592 4629 19601
rect 4587 19552 4588 19592
rect 4628 19552 4629 19592
rect 4587 19543 4629 19552
rect 4300 19459 4340 19468
rect 4588 19256 4628 19543
rect 4588 19207 4628 19216
rect 4684 19256 4724 19265
rect 4684 19097 4724 19216
rect 4683 19088 4725 19097
rect 4683 19048 4684 19088
rect 4724 19048 4725 19088
rect 4683 19039 4725 19048
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4587 18752 4629 18761
rect 4876 18752 4916 22996
rect 4972 21617 5012 24415
rect 5068 23129 5108 28876
rect 5259 24548 5301 24557
rect 5259 24508 5260 24548
rect 5300 24508 5301 24548
rect 5259 24499 5301 24508
rect 5260 24044 5300 24499
rect 5260 23995 5300 24004
rect 5067 23120 5109 23129
rect 5067 23080 5068 23120
rect 5108 23080 5109 23120
rect 5067 23071 5109 23080
rect 5356 22028 5396 31308
rect 5548 30428 5588 33823
rect 5740 33041 5780 36679
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 83211 36224 83253 36233
rect 83211 36184 83212 36224
rect 83252 36184 83253 36224
rect 83211 36175 83253 36184
rect 91600 36182 91642 36191
rect 12171 35888 12213 35897
rect 12171 35848 12172 35888
rect 12212 35848 12213 35888
rect 12171 35839 12213 35848
rect 12459 35888 12501 35897
rect 12459 35848 12460 35888
rect 12500 35848 12501 35888
rect 12459 35839 12501 35848
rect 13324 35888 13364 35897
rect 12172 35754 12212 35839
rect 12460 35754 12500 35839
rect 13324 34385 13364 35848
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 32620 35216 32660 35225
rect 15052 35132 15092 35141
rect 14860 35092 15052 35132
rect 13323 34376 13365 34385
rect 13323 34336 13324 34376
rect 13364 34336 13365 34376
rect 13323 34327 13365 34336
rect 5931 34208 5973 34217
rect 5931 34168 5932 34208
rect 5972 34168 5973 34208
rect 5931 34159 5973 34168
rect 5932 33209 5972 34159
rect 13324 33881 13364 34327
rect 14379 34208 14421 34217
rect 14379 34168 14380 34208
rect 14420 34168 14421 34208
rect 14379 34159 14421 34168
rect 14668 34208 14708 34217
rect 13323 33872 13365 33881
rect 13323 33832 13324 33872
rect 13364 33832 13365 33872
rect 13323 33823 13365 33832
rect 11115 33704 11157 33713
rect 11115 33664 11116 33704
rect 11156 33664 11157 33704
rect 11115 33655 11157 33664
rect 13996 33704 14036 33713
rect 5931 33200 5973 33209
rect 5931 33160 5932 33200
rect 5972 33160 5973 33200
rect 5931 33151 5973 33160
rect 5739 33032 5781 33041
rect 5739 32992 5740 33032
rect 5780 32992 5781 33032
rect 5739 32983 5781 32992
rect 5740 32864 5780 32873
rect 5932 32864 5972 33151
rect 9291 33116 9333 33125
rect 9291 33076 9292 33116
rect 9332 33076 9333 33116
rect 9291 33067 9333 33076
rect 7083 33032 7125 33041
rect 7083 32992 7084 33032
rect 7124 32992 7125 33032
rect 7083 32983 7125 32992
rect 7275 33032 7317 33041
rect 7275 32992 7276 33032
rect 7316 32992 7317 33032
rect 7275 32983 7317 32992
rect 7084 32873 7124 32983
rect 5780 32824 5972 32864
rect 6604 32864 6644 32873
rect 5740 32815 5780 32824
rect 6604 32705 6644 32824
rect 7083 32864 7125 32873
rect 7083 32824 7084 32864
rect 7124 32824 7125 32864
rect 7083 32815 7125 32824
rect 6603 32696 6645 32705
rect 6603 32656 6604 32696
rect 6644 32656 6645 32696
rect 6603 32647 6645 32656
rect 5739 32528 5781 32537
rect 5739 32488 5740 32528
rect 5780 32488 5781 32528
rect 5739 32479 5781 32488
rect 5740 31700 5780 32479
rect 6027 31856 6069 31865
rect 6027 31816 6028 31856
rect 6068 31816 6069 31856
rect 6027 31807 6069 31816
rect 5740 31660 5876 31700
rect 5680 31352 5720 31361
rect 5720 31312 5732 31348
rect 5680 31303 5732 31312
rect 5692 31268 5732 31303
rect 5836 31268 5876 31660
rect 5692 31228 5972 31268
rect 5548 30388 5684 30428
rect 5451 30260 5493 30269
rect 5451 30220 5452 30260
rect 5492 30220 5493 30260
rect 5451 30211 5493 30220
rect 5452 27656 5492 30211
rect 5644 29168 5684 30388
rect 5836 29672 5876 29681
rect 5836 29177 5876 29632
rect 5644 28328 5684 29128
rect 5835 29168 5877 29177
rect 5835 29128 5836 29168
rect 5876 29128 5877 29168
rect 5835 29119 5877 29128
rect 5644 28279 5684 28288
rect 5452 27607 5492 27616
rect 5836 27656 5876 27665
rect 5836 27077 5876 27616
rect 5835 27068 5877 27077
rect 5835 27028 5836 27068
rect 5876 27028 5877 27068
rect 5835 27019 5877 27028
rect 5932 26237 5972 31228
rect 5931 26228 5973 26237
rect 5931 26188 5932 26228
rect 5972 26188 5973 26228
rect 5931 26179 5973 26188
rect 5835 25136 5877 25145
rect 5835 25096 5836 25136
rect 5876 25096 5877 25136
rect 5835 25087 5877 25096
rect 5836 25002 5876 25087
rect 5739 24548 5781 24557
rect 5739 24508 5740 24548
rect 5780 24508 5781 24548
rect 5739 24499 5781 24508
rect 5260 21988 5396 22028
rect 4971 21608 5013 21617
rect 4971 21568 4972 21608
rect 5012 21568 5013 21608
rect 4971 21559 5013 21568
rect 5164 21020 5204 21029
rect 5260 21020 5300 21988
rect 5204 20980 5300 21020
rect 5164 20971 5204 20980
rect 5260 20609 5300 20980
rect 5259 20600 5301 20609
rect 5259 20560 5260 20600
rect 5300 20560 5301 20600
rect 5259 20551 5301 20560
rect 4971 20096 5013 20105
rect 4971 20056 4972 20096
rect 5012 20056 5013 20096
rect 4971 20047 5013 20056
rect 4972 19256 5012 20047
rect 5012 19216 5108 19256
rect 4972 19207 5012 19216
rect 4971 19088 5013 19097
rect 4971 19048 4972 19088
rect 5012 19048 5013 19088
rect 4971 19039 5013 19048
rect 4587 18712 4588 18752
rect 4628 18712 4629 18752
rect 4587 18703 4629 18712
rect 4684 18712 4916 18752
rect 3819 18668 3861 18677
rect 3819 18628 3820 18668
rect 3860 18628 3861 18668
rect 3819 18619 3861 18628
rect 3436 18584 3476 18593
rect 3820 18584 3860 18619
rect 3476 18544 3572 18584
rect 3436 18535 3476 18544
rect 3244 18341 3284 18426
rect 2859 18332 2901 18341
rect 2859 18292 2860 18332
rect 2900 18292 2901 18332
rect 2859 18283 2901 18292
rect 3243 18332 3285 18341
rect 3243 18292 3244 18332
rect 3284 18292 3285 18332
rect 3243 18283 3285 18292
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3532 17996 3572 18544
rect 3820 18534 3860 18544
rect 4011 18332 4053 18341
rect 4011 18292 4012 18332
rect 4052 18292 4053 18332
rect 4011 18283 4053 18292
rect 3916 17996 3956 18005
rect 3532 17956 3916 17996
rect 3916 17947 3956 17956
rect 2668 17779 2708 17788
rect 3244 17828 3284 17837
rect 1900 17695 1940 17704
rect 1996 17744 2036 17753
rect 1803 17660 1845 17669
rect 1803 17620 1804 17660
rect 1844 17620 1845 17660
rect 1803 17611 1845 17620
rect 1996 17300 2036 17704
rect 2283 17744 2325 17753
rect 3244 17744 3284 17788
rect 2283 17704 2284 17744
rect 2324 17704 2325 17744
rect 2283 17695 2325 17704
rect 2956 17704 3284 17744
rect 2284 17610 2324 17695
rect 2667 17660 2709 17669
rect 2667 17620 2668 17660
rect 2708 17620 2709 17660
rect 2667 17611 2709 17620
rect 1996 17260 2132 17300
rect 1996 17072 2036 17081
rect 1612 16484 1652 16493
rect 1996 16484 2036 17032
rect 1652 16444 2036 16484
rect 1612 16435 1652 16444
rect 1516 16276 1652 16316
rect 1419 16064 1461 16073
rect 1419 16024 1420 16064
rect 1460 16024 1461 16064
rect 1419 16015 1461 16024
rect 1420 15930 1460 16015
rect 1420 15560 1460 15569
rect 1324 15520 1420 15560
rect 459 15511 501 15520
rect 843 15476 885 15485
rect 843 15436 844 15476
rect 884 15436 885 15476
rect 843 15427 885 15436
rect 844 15342 884 15427
rect 652 15308 692 15317
rect 652 14897 692 15268
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 1228 14720 1268 14729
rect 844 14636 884 14645
rect 884 14596 1076 14636
rect 844 14587 884 14596
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 652 13880 692 13999
rect 652 13831 692 13840
rect 844 13964 884 13973
rect 844 13637 884 13924
rect 1036 13880 1076 14596
rect 1228 14561 1268 14680
rect 1227 14552 1269 14561
rect 1227 14512 1228 14552
rect 1268 14512 1269 14552
rect 1227 14503 1269 14512
rect 1324 13880 1364 13889
rect 1036 13840 1324 13880
rect 1324 13831 1364 13840
rect 1420 13721 1460 15520
rect 1515 15560 1557 15569
rect 1515 15520 1516 15560
rect 1556 15520 1557 15560
rect 1515 15511 1557 15520
rect 1612 15560 1652 16276
rect 2092 16241 2132 17260
rect 2380 17072 2420 17081
rect 2380 16484 2420 17032
rect 2572 16484 2612 16493
rect 2380 16444 2572 16484
rect 2572 16435 2612 16444
rect 1899 16232 1941 16241
rect 1899 16192 1900 16232
rect 1940 16192 1941 16232
rect 1899 16183 1941 16192
rect 1996 16232 2036 16241
rect 1900 16098 1940 16183
rect 1899 15980 1941 15989
rect 1899 15940 1900 15980
rect 1940 15940 1941 15980
rect 1899 15931 1941 15940
rect 1707 15644 1749 15653
rect 1707 15604 1708 15644
rect 1748 15604 1749 15644
rect 1707 15595 1749 15604
rect 1612 15511 1652 15520
rect 1131 13712 1173 13721
rect 1131 13672 1132 13712
rect 1172 13672 1173 13712
rect 1131 13663 1173 13672
rect 1419 13712 1461 13721
rect 1419 13672 1420 13712
rect 1460 13672 1461 13712
rect 1419 13663 1461 13672
rect 843 13628 885 13637
rect 843 13588 844 13628
rect 884 13588 885 13628
rect 843 13579 885 13588
rect 844 13292 884 13301
rect 748 13252 844 13292
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 748 12536 788 13252
rect 844 13243 884 13252
rect 843 13040 885 13049
rect 843 13000 844 13040
rect 884 13000 885 13040
rect 843 12991 885 13000
rect 460 12496 788 12536
rect 844 12536 884 12991
rect 460 7220 500 12496
rect 844 12487 884 12496
rect 1132 12536 1172 13663
rect 1419 13544 1461 13553
rect 1419 13504 1420 13544
rect 1460 13504 1461 13544
rect 1419 13495 1461 13504
rect 1132 12487 1172 12496
rect 1324 12536 1364 12545
rect 940 12452 980 12461
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 652 11948 692 12319
rect 652 11899 692 11908
rect 844 11780 884 11789
rect 748 11740 844 11780
rect 555 11528 597 11537
rect 555 11488 556 11528
rect 596 11488 597 11528
rect 555 11479 597 11488
rect 556 11192 596 11479
rect 652 11192 692 11201
rect 556 11152 652 11192
rect 652 11143 692 11152
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9680 692 9799
rect 652 9631 692 9640
rect 748 9260 788 11740
rect 844 11731 884 11740
rect 940 11285 980 12412
rect 1324 11948 1364 12496
rect 1324 11899 1364 11908
rect 1420 11696 1460 13495
rect 1516 13208 1556 15511
rect 1708 15056 1748 15595
rect 1803 15560 1845 15569
rect 1803 15520 1804 15560
rect 1844 15520 1845 15560
rect 1803 15511 1845 15520
rect 1804 15392 1844 15511
rect 1804 15343 1844 15352
rect 1612 15016 1748 15056
rect 1612 14132 1652 15016
rect 1612 14083 1652 14092
rect 1708 14048 1748 14057
rect 1900 14048 1940 15931
rect 1996 15812 2036 16192
rect 2091 16232 2133 16241
rect 2091 16192 2092 16232
rect 2132 16192 2133 16232
rect 2091 16183 2133 16192
rect 2284 16232 2324 16241
rect 2284 16073 2324 16192
rect 2283 16064 2325 16073
rect 2283 16024 2284 16064
rect 2324 16024 2325 16064
rect 2283 16015 2325 16024
rect 2572 16064 2612 16073
rect 2283 15896 2325 15905
rect 2283 15856 2284 15896
rect 2324 15856 2325 15896
rect 2283 15847 2325 15856
rect 1996 15772 2132 15812
rect 2092 15653 2132 15772
rect 2091 15644 2133 15653
rect 2091 15604 2092 15644
rect 2132 15604 2133 15644
rect 2091 15595 2133 15604
rect 1995 15560 2037 15569
rect 1995 15520 1996 15560
rect 2036 15520 2037 15560
rect 1995 15511 2037 15520
rect 2188 15560 2228 15569
rect 1996 15426 2036 15511
rect 2091 15476 2133 15485
rect 2091 15436 2092 15476
rect 2132 15436 2133 15476
rect 2091 15427 2133 15436
rect 2092 15342 2132 15427
rect 2091 14720 2133 14729
rect 2091 14680 2092 14720
rect 2132 14680 2133 14720
rect 2091 14671 2133 14680
rect 1996 14048 2036 14057
rect 1748 14008 1844 14048
rect 1900 14008 1996 14048
rect 1708 13999 1748 14008
rect 1707 13712 1749 13721
rect 1707 13672 1708 13712
rect 1748 13672 1749 13712
rect 1707 13663 1749 13672
rect 1516 13049 1556 13168
rect 1708 13208 1748 13663
rect 1804 13553 1844 14008
rect 1899 13628 1941 13637
rect 1899 13588 1900 13628
rect 1940 13588 1941 13628
rect 1899 13579 1941 13588
rect 1803 13544 1845 13553
rect 1803 13504 1804 13544
rect 1844 13504 1845 13544
rect 1803 13495 1845 13504
rect 1900 13460 1940 13579
rect 1900 13411 1940 13420
rect 1996 13292 2036 14008
rect 1708 13159 1748 13168
rect 1900 13252 2036 13292
rect 1515 13040 1557 13049
rect 1515 13000 1516 13040
rect 1556 13000 1557 13040
rect 1515 12991 1557 13000
rect 1612 13040 1652 13049
rect 1612 11873 1652 13000
rect 1900 12872 1940 13252
rect 1996 13197 2036 13206
rect 1996 13049 2036 13157
rect 1995 13040 2037 13049
rect 1995 13000 1996 13040
rect 2036 13000 2037 13040
rect 1995 12991 2037 13000
rect 1900 12832 2036 12872
rect 1707 12536 1749 12545
rect 1707 12496 1708 12536
rect 1748 12496 1749 12536
rect 1707 12487 1749 12496
rect 1708 12402 1748 12487
rect 1611 11864 1653 11873
rect 1611 11824 1612 11864
rect 1652 11824 1653 11864
rect 1611 11815 1653 11824
rect 1612 11696 1652 11705
rect 1420 11656 1612 11696
rect 1612 11647 1652 11656
rect 1708 11696 1748 11705
rect 1996 11696 2036 12832
rect 1748 11656 1844 11696
rect 1708 11647 1748 11656
rect 939 11276 981 11285
rect 939 11236 940 11276
rect 980 11236 981 11276
rect 939 11227 981 11236
rect 1611 11276 1653 11285
rect 1611 11236 1612 11276
rect 1652 11236 1653 11276
rect 1611 11227 1653 11236
rect 1420 11108 1460 11117
rect 940 11068 1420 11108
rect 843 10940 885 10949
rect 843 10900 844 10940
rect 884 10900 885 10940
rect 843 10891 885 10900
rect 844 10806 884 10891
rect 843 10100 885 10109
rect 843 10060 844 10100
rect 884 10060 885 10100
rect 843 10051 885 10060
rect 844 9966 884 10051
rect 844 9428 884 9437
rect 940 9428 980 11068
rect 1420 11059 1460 11068
rect 1612 11024 1652 11227
rect 1707 11192 1749 11201
rect 1707 11152 1708 11192
rect 1748 11152 1749 11192
rect 1707 11143 1749 11152
rect 1708 11058 1748 11143
rect 1228 10940 1268 10949
rect 1132 10900 1228 10940
rect 1035 10772 1077 10781
rect 1035 10732 1036 10772
rect 1076 10732 1077 10772
rect 1035 10723 1077 10732
rect 1036 10638 1076 10723
rect 1036 9680 1076 9689
rect 1132 9680 1172 10900
rect 1228 10891 1268 10900
rect 1419 10940 1461 10949
rect 1419 10900 1420 10940
rect 1460 10900 1461 10940
rect 1419 10891 1461 10900
rect 1227 10352 1269 10361
rect 1227 10312 1228 10352
rect 1268 10312 1269 10352
rect 1227 10303 1269 10312
rect 1228 10184 1268 10303
rect 1228 10135 1268 10144
rect 1323 10184 1365 10193
rect 1323 10144 1324 10184
rect 1364 10144 1365 10184
rect 1323 10135 1365 10144
rect 1324 9848 1364 10135
rect 1076 9640 1172 9680
rect 1228 9808 1364 9848
rect 1036 9631 1076 9640
rect 1228 9512 1268 9808
rect 1228 9463 1268 9472
rect 1324 9680 1364 9689
rect 884 9388 980 9428
rect 844 9379 884 9388
rect 748 9220 980 9260
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 652 8924 692 8959
rect 652 8873 692 8884
rect 843 8840 885 8849
rect 843 8800 844 8840
rect 884 8800 885 8840
rect 843 8791 885 8800
rect 844 8756 884 8791
rect 844 8705 884 8716
rect 652 8168 692 8177
rect 652 7337 692 8128
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 460 7180 596 7220
rect 556 7085 596 7180
rect 940 7169 980 9220
rect 1036 8504 1076 8513
rect 1036 8177 1076 8464
rect 1324 8420 1364 9640
rect 1420 9176 1460 10891
rect 1612 10193 1652 10984
rect 1804 10193 1844 11656
rect 1996 11033 2036 11656
rect 1995 11024 2037 11033
rect 1995 10984 1996 11024
rect 2036 10984 2037 11024
rect 1995 10975 2037 10984
rect 1611 10184 1653 10193
rect 1611 10144 1612 10184
rect 1652 10144 1653 10184
rect 1611 10135 1653 10144
rect 1803 10184 1845 10193
rect 1803 10144 1804 10184
rect 1844 10144 1845 10184
rect 1803 10135 1845 10144
rect 1515 10100 1557 10109
rect 1515 10060 1516 10100
rect 1556 10060 1557 10100
rect 1515 10051 1557 10060
rect 1516 9344 1556 10051
rect 1516 9295 1556 9304
rect 1420 9136 1556 9176
rect 1516 9092 1556 9136
rect 1516 9052 1559 9092
rect 1519 9008 1559 9052
rect 1516 8968 1559 9008
rect 1420 8849 1460 8934
rect 1419 8840 1461 8849
rect 1419 8800 1420 8840
rect 1460 8800 1461 8840
rect 1419 8791 1461 8800
rect 1516 8672 1556 8968
rect 1228 8380 1364 8420
rect 1420 8632 1556 8672
rect 1612 8672 1652 10135
rect 1804 9596 1844 10135
rect 1804 9547 1844 9556
rect 1900 9512 1940 9521
rect 1996 9512 2036 10975
rect 2092 10184 2132 14671
rect 2188 14477 2228 15520
rect 2187 14468 2229 14477
rect 2187 14428 2188 14468
rect 2228 14428 2229 14468
rect 2187 14419 2229 14428
rect 2284 13973 2324 15847
rect 2572 15821 2612 16024
rect 2571 15812 2613 15821
rect 2571 15772 2572 15812
rect 2612 15772 2613 15812
rect 2571 15763 2613 15772
rect 2572 14561 2612 15763
rect 2571 14552 2613 14561
rect 2571 14512 2572 14552
rect 2612 14512 2613 14552
rect 2571 14503 2613 14512
rect 2283 13964 2325 13973
rect 2283 13924 2284 13964
rect 2324 13924 2325 13964
rect 2283 13915 2325 13924
rect 2187 12536 2229 12545
rect 2187 12496 2188 12536
rect 2228 12496 2229 12536
rect 2187 12487 2229 12496
rect 2188 10361 2228 12487
rect 2187 10352 2229 10361
rect 2187 10312 2188 10352
rect 2228 10312 2229 10352
rect 2187 10303 2229 10312
rect 2092 10135 2132 10144
rect 2188 9512 2228 9521
rect 1996 9472 2188 9512
rect 1900 8933 1940 9472
rect 2188 9463 2228 9472
rect 2284 9344 2324 13915
rect 2571 13208 2613 13217
rect 2571 13168 2572 13208
rect 2612 13168 2613 13208
rect 2571 13159 2613 13168
rect 2572 12536 2612 13159
rect 2572 12487 2612 12496
rect 2668 12284 2708 17611
rect 2860 17576 2900 17585
rect 2956 17576 2996 17704
rect 4012 17669 4052 18283
rect 4300 17753 4340 17838
rect 4299 17744 4341 17753
rect 4299 17704 4300 17744
rect 4340 17704 4341 17744
rect 4299 17695 4341 17704
rect 4588 17744 4628 18703
rect 4684 18584 4724 18712
rect 4684 18535 4724 18544
rect 4588 17695 4628 17704
rect 4011 17660 4053 17669
rect 4011 17620 4012 17660
rect 4052 17620 4053 17660
rect 4011 17611 4053 17620
rect 4204 17660 4244 17669
rect 2900 17536 2996 17576
rect 3052 17576 3092 17585
rect 4204 17576 4244 17620
rect 4299 17576 4341 17585
rect 4204 17536 4300 17576
rect 4340 17536 4341 17576
rect 2860 17300 2900 17536
rect 2860 17260 2996 17300
rect 2763 16820 2805 16829
rect 2763 16780 2764 16820
rect 2804 16780 2805 16820
rect 2763 16771 2805 16780
rect 2764 16316 2804 16771
rect 2764 15905 2804 16276
rect 2763 15896 2805 15905
rect 2763 15856 2764 15896
rect 2804 15856 2805 15896
rect 2763 15847 2805 15856
rect 2572 12244 2708 12284
rect 2475 11864 2517 11873
rect 2475 11824 2476 11864
rect 2516 11824 2517 11864
rect 2475 11815 2517 11824
rect 2188 9304 2324 9344
rect 1899 8924 1941 8933
rect 1899 8884 1900 8924
rect 1940 8884 1941 8924
rect 1899 8875 1941 8884
rect 1035 8168 1077 8177
rect 1035 8128 1036 8168
rect 1076 8128 1077 8168
rect 1035 8119 1077 8128
rect 939 7160 981 7169
rect 939 7120 940 7160
rect 980 7120 981 7160
rect 939 7111 981 7120
rect 555 7076 597 7085
rect 555 7036 556 7076
rect 596 7036 597 7076
rect 555 7027 597 7036
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 1228 5657 1268 8380
rect 1420 8336 1460 8632
rect 1612 8588 1652 8632
rect 1996 8672 2036 8681
rect 2188 8672 2228 9304
rect 2379 8924 2421 8933
rect 2379 8884 2380 8924
rect 2420 8884 2421 8924
rect 2379 8875 2421 8884
rect 2036 8632 2228 8672
rect 2284 8672 2324 8681
rect 1996 8623 2036 8632
rect 1324 8296 1460 8336
rect 1516 8548 1652 8588
rect 1324 7160 1364 8296
rect 1324 7111 1364 7120
rect 1420 7160 1460 7169
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 1227 5648 1269 5657
rect 1227 5608 1228 5648
rect 1268 5608 1269 5648
rect 1227 5599 1269 5608
rect 267 5564 309 5573
rect 267 5524 268 5564
rect 308 5524 309 5564
rect 267 5515 309 5524
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 652 5144 692 5153
rect 652 4817 692 5104
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 1420 3641 1460 7120
rect 1516 5153 1556 8548
rect 1707 8504 1749 8513
rect 1707 8464 1708 8504
rect 1748 8464 1749 8504
rect 1707 8455 1749 8464
rect 1708 8370 1748 8455
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 1708 7160 1748 7169
rect 1612 7026 1652 7111
rect 1515 5144 1557 5153
rect 1515 5104 1516 5144
rect 1556 5104 1557 5144
rect 1515 5095 1557 5104
rect 1708 3725 1748 7120
rect 1996 7160 2036 7169
rect 1899 7076 1941 7085
rect 1899 7036 1900 7076
rect 1940 7036 1941 7076
rect 1899 7027 1941 7036
rect 1900 6942 1940 7027
rect 1707 3716 1749 3725
rect 1707 3676 1708 3716
rect 1748 3676 1749 3716
rect 1707 3667 1749 3676
rect 652 3632 692 3641
rect 652 3137 692 3592
rect 1419 3632 1461 3641
rect 1419 3592 1420 3632
rect 1460 3592 1461 3632
rect 1419 3583 1461 3592
rect 1996 3305 2036 7120
rect 2092 7085 2132 8632
rect 2284 7169 2324 8632
rect 2380 8672 2420 8875
rect 2380 8623 2420 8632
rect 2283 7160 2325 7169
rect 2283 7120 2284 7160
rect 2324 7120 2325 7160
rect 2283 7111 2325 7120
rect 2091 7076 2133 7085
rect 2091 7036 2092 7076
rect 2132 7036 2133 7076
rect 2091 7027 2133 7036
rect 2476 3893 2516 11815
rect 2572 4061 2612 12244
rect 2668 8840 2708 8849
rect 2708 8800 2900 8840
rect 2668 8791 2708 8800
rect 2860 8672 2900 8800
rect 2860 8623 2900 8632
rect 2956 4229 2996 17260
rect 3052 16829 3092 17536
rect 4299 17527 4341 17536
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4780 17081 4820 18712
rect 4875 17744 4917 17753
rect 4875 17704 4876 17744
rect 4916 17704 4917 17744
rect 4875 17695 4917 17704
rect 4876 17324 4916 17695
rect 4972 17585 5012 19039
rect 5068 18761 5108 19216
rect 5067 18752 5109 18761
rect 5067 18712 5068 18752
rect 5108 18712 5109 18752
rect 5067 18703 5109 18712
rect 4971 17576 5013 17585
rect 4971 17536 4972 17576
rect 5012 17536 5013 17576
rect 4971 17527 5013 17536
rect 5740 17333 5780 24499
rect 5836 22112 5876 22121
rect 5876 22072 5972 22112
rect 5836 22063 5876 22072
rect 5932 21701 5972 22072
rect 5931 21692 5973 21701
rect 5931 21652 5932 21692
rect 5972 21652 5973 21692
rect 5931 21643 5973 21652
rect 5835 20012 5877 20021
rect 5835 19972 5836 20012
rect 5876 19972 5877 20012
rect 5835 19963 5877 19972
rect 5836 19878 5876 19963
rect 5836 18332 5876 18341
rect 5836 17585 5876 18292
rect 5835 17576 5877 17585
rect 5835 17536 5836 17576
rect 5876 17536 5877 17576
rect 5835 17527 5877 17536
rect 4971 17324 5013 17333
rect 4876 17284 4972 17324
rect 5012 17284 5013 17324
rect 4971 17275 5013 17284
rect 5739 17324 5781 17333
rect 5739 17284 5740 17324
rect 5780 17300 5781 17324
rect 5932 17300 5972 21643
rect 6028 20021 6068 31807
rect 6411 31100 6453 31109
rect 6411 31060 6412 31100
rect 6452 31060 6453 31100
rect 6411 31051 6453 31060
rect 6412 23045 6452 31051
rect 6604 27665 6644 32647
rect 6891 31268 6933 31277
rect 6891 31228 6892 31268
rect 6932 31228 6933 31268
rect 6891 31219 6933 31228
rect 6603 27656 6645 27665
rect 6603 27616 6604 27656
rect 6644 27616 6645 27656
rect 6603 27607 6645 27616
rect 6411 23036 6453 23045
rect 6411 22996 6412 23036
rect 6452 22996 6453 23036
rect 6411 22987 6453 22996
rect 6027 20012 6069 20021
rect 6027 19972 6028 20012
rect 6068 19972 6069 20012
rect 6027 19963 6069 19972
rect 6028 19601 6068 19963
rect 6027 19592 6069 19601
rect 6027 19552 6028 19592
rect 6068 19552 6069 19592
rect 6027 19543 6069 19552
rect 5780 17284 5876 17300
rect 5739 17275 5876 17284
rect 3243 17072 3285 17081
rect 3243 17032 3244 17072
rect 3284 17032 3285 17072
rect 3243 17023 3285 17032
rect 4779 17072 4821 17081
rect 4779 17032 4780 17072
rect 4820 17032 4821 17072
rect 4779 17023 4821 17032
rect 3244 16938 3284 17023
rect 3051 16820 3093 16829
rect 3051 16780 3052 16820
rect 3092 16780 3093 16820
rect 3051 16771 3093 16780
rect 4396 16820 4436 16829
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 4396 16577 4436 16780
rect 4395 16568 4437 16577
rect 4395 16528 4396 16568
rect 4436 16528 4437 16568
rect 4395 16519 4437 16528
rect 4396 16241 4436 16519
rect 3820 16232 3860 16241
rect 3436 16148 3476 16157
rect 3476 16108 3764 16148
rect 3436 16099 3476 16108
rect 3627 15896 3669 15905
rect 3627 15856 3628 15896
rect 3668 15856 3669 15896
rect 3627 15847 3669 15856
rect 3531 15476 3573 15485
rect 3531 15436 3532 15476
rect 3572 15436 3573 15476
rect 3531 15427 3573 15436
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 3244 14972 3284 14981
rect 3532 14972 3572 15427
rect 3284 14932 3572 14972
rect 3244 14923 3284 14932
rect 3628 14720 3668 15847
rect 3724 15812 3764 16108
rect 3820 15989 3860 16192
rect 4395 16232 4437 16241
rect 4395 16192 4396 16232
rect 4436 16192 4437 16232
rect 4395 16183 4437 16192
rect 4684 16232 4724 16241
rect 4780 16232 4820 17023
rect 4724 16192 4820 16232
rect 4684 16183 4724 16192
rect 3819 15980 3861 15989
rect 3819 15940 3820 15980
rect 3860 15940 3861 15980
rect 3819 15931 3861 15940
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 3724 15772 4244 15812
rect 4204 15392 4244 15772
rect 4491 15644 4533 15653
rect 4491 15604 4492 15644
rect 4532 15604 4533 15644
rect 4491 15595 4533 15604
rect 4492 15510 4532 15595
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 4588 15426 4628 15511
rect 4204 15343 4244 15352
rect 3820 14720 3860 14729
rect 3628 14680 3820 14720
rect 3436 14636 3476 14645
rect 3476 14596 3668 14636
rect 3436 14587 3476 14596
rect 3628 13880 3668 14596
rect 3628 13831 3668 13840
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 3724 13292 3764 14680
rect 3820 14671 3860 14680
rect 4683 14720 4725 14729
rect 4780 14720 4820 16192
rect 4972 15653 5012 17275
rect 5740 17260 5876 17275
rect 5932 17260 6068 17300
rect 5836 16484 5876 17260
rect 5836 16435 5876 16444
rect 4971 15644 5013 15653
rect 4971 15604 4972 15644
rect 5012 15604 5013 15644
rect 4971 15595 5013 15604
rect 4683 14680 4684 14720
rect 4724 14680 4820 14720
rect 4876 15560 4916 15569
rect 4683 14671 4725 14680
rect 4684 14586 4724 14671
rect 3819 14552 3861 14561
rect 3819 14512 3820 14552
rect 3860 14512 3861 14552
rect 3819 14503 3861 14512
rect 3532 13252 3764 13292
rect 3436 13124 3476 13133
rect 3436 12377 3476 13084
rect 3435 12368 3477 12377
rect 3435 12328 3436 12368
rect 3476 12328 3477 12368
rect 3435 12319 3477 12328
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3436 11612 3476 11621
rect 3436 10865 3476 11572
rect 3435 10856 3477 10865
rect 3435 10816 3436 10856
rect 3476 10816 3477 10856
rect 3435 10807 3477 10816
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3244 10268 3284 10279
rect 3532 10268 3572 13252
rect 3820 13208 3860 14503
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3915 14132 3957 14141
rect 3915 14092 3916 14132
rect 3956 14092 3957 14132
rect 3915 14083 3957 14092
rect 3916 13998 3956 14083
rect 4011 14048 4053 14057
rect 4011 14008 4012 14048
rect 4052 14008 4053 14048
rect 4011 13999 4053 14008
rect 4203 14048 4245 14057
rect 4203 14008 4204 14048
rect 4244 14008 4245 14048
rect 4203 13999 4245 14008
rect 4300 14048 4340 14059
rect 4012 13914 4052 13999
rect 4011 13460 4053 13469
rect 4011 13420 4012 13460
rect 4052 13420 4053 13460
rect 4011 13411 4053 13420
rect 3820 12965 3860 13168
rect 3627 12956 3669 12965
rect 3627 12916 3628 12956
rect 3668 12916 3669 12956
rect 3627 12907 3669 12916
rect 3819 12956 3861 12965
rect 3819 12916 3820 12956
rect 3860 12916 3861 12956
rect 3819 12907 3861 12916
rect 3628 11696 3668 12907
rect 3916 12377 3956 12462
rect 3915 12368 3957 12377
rect 3915 12328 3916 12368
rect 3956 12328 3957 12368
rect 3915 12319 3957 12328
rect 3724 12284 3764 12293
rect 3724 12200 3764 12244
rect 4012 12200 4052 13411
rect 4204 12620 4244 13999
rect 4300 13973 4340 14008
rect 4299 13964 4341 13973
rect 4299 13924 4300 13964
rect 4340 13924 4341 13964
rect 4299 13915 4341 13924
rect 4683 13208 4725 13217
rect 4683 13168 4684 13208
rect 4724 13168 4820 13208
rect 4683 13159 4725 13168
rect 4684 13074 4724 13159
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4204 12571 4244 12580
rect 3724 12160 4052 12200
rect 4300 12536 4340 12545
rect 3820 11696 3860 11705
rect 3628 11656 3820 11696
rect 3723 10856 3765 10865
rect 3723 10816 3724 10856
rect 3764 10816 3765 10856
rect 3723 10807 3765 10816
rect 3724 10722 3764 10807
rect 3820 10361 3860 11656
rect 4300 11528 4340 12496
rect 4588 12536 4628 12545
rect 4588 11537 4628 12496
rect 4684 11696 4724 11705
rect 4780 11696 4820 13168
rect 4724 11656 4820 11696
rect 4684 11647 4724 11656
rect 4204 11488 4340 11528
rect 4587 11528 4629 11537
rect 4587 11488 4588 11528
rect 4628 11488 4629 11528
rect 4204 11285 4244 11488
rect 4587 11479 4629 11488
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4011 11276 4053 11285
rect 4011 11236 4012 11276
rect 4052 11236 4053 11276
rect 4011 11227 4053 11236
rect 4203 11276 4245 11285
rect 4203 11236 4204 11276
rect 4244 11236 4245 11276
rect 4203 11227 4245 11236
rect 4012 11108 4052 11227
rect 4012 11059 4052 11068
rect 4108 11024 4148 11035
rect 4108 10949 4148 10984
rect 4395 11024 4437 11033
rect 4395 10984 4396 11024
rect 4436 10984 4437 11024
rect 4395 10975 4437 10984
rect 4587 11024 4629 11033
rect 4587 10984 4588 11024
rect 4628 10984 4629 11024
rect 4587 10975 4629 10984
rect 4107 10940 4149 10949
rect 4107 10900 4108 10940
rect 4148 10900 4244 10940
rect 4107 10891 4149 10900
rect 4107 10604 4149 10613
rect 4107 10564 4108 10604
rect 4148 10564 4149 10604
rect 4107 10555 4149 10564
rect 3819 10352 3861 10361
rect 3819 10312 3820 10352
rect 3860 10312 3861 10352
rect 3819 10303 3861 10312
rect 3244 10193 3284 10228
rect 3340 10228 3572 10268
rect 3243 10184 3285 10193
rect 3243 10144 3244 10184
rect 3284 10144 3285 10184
rect 3243 10135 3285 10144
rect 3340 9260 3380 10228
rect 3820 10184 3860 10303
rect 3820 10135 3860 10144
rect 3436 10100 3476 10109
rect 3476 10060 3764 10100
rect 3436 10051 3476 10060
rect 3724 9512 3764 10060
rect 3724 9472 4052 9512
rect 4012 9344 4052 9472
rect 4012 9295 4052 9304
rect 3340 9220 3572 9260
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3244 8672 3284 8681
rect 3532 8672 3572 9220
rect 4108 9176 4148 10555
rect 4204 9680 4244 10900
rect 4396 10890 4436 10975
rect 4588 10016 4628 10975
rect 4684 10184 4724 10193
rect 4780 10184 4820 11656
rect 4876 11537 4916 15520
rect 5931 15140 5973 15149
rect 5931 15100 5932 15140
rect 5972 15100 5973 15140
rect 5931 15091 5973 15100
rect 5835 14552 5877 14561
rect 5835 14512 5836 14552
rect 5876 14512 5877 14552
rect 5835 14503 5877 14512
rect 5836 14141 5876 14503
rect 5835 14132 5877 14141
rect 5835 14092 5836 14132
rect 5876 14092 5877 14132
rect 5835 14083 5877 14092
rect 5932 14057 5972 15091
rect 5931 14048 5973 14057
rect 5931 14008 5932 14048
rect 5972 14008 5973 14048
rect 5931 13999 5973 14008
rect 5836 13460 5876 13469
rect 5932 13460 5972 13999
rect 5876 13420 5972 13460
rect 5836 13411 5876 13420
rect 5836 11780 5876 11789
rect 4875 11528 4917 11537
rect 4875 11488 4876 11528
rect 4916 11488 4917 11528
rect 4875 11479 4917 11488
rect 4876 11033 4916 11479
rect 4971 11444 5013 11453
rect 4971 11404 4972 11444
rect 5012 11404 5013 11444
rect 4971 11395 5013 11404
rect 4875 11024 4917 11033
rect 4875 10984 4876 11024
rect 4916 10984 4917 11024
rect 4875 10975 4917 10984
rect 4724 10144 4916 10184
rect 4684 10135 4724 10144
rect 4588 9976 4820 10016
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4204 9640 4340 9680
rect 4300 9596 4340 9640
rect 4300 9547 4340 9556
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4684 9512 4724 9521
rect 4780 9512 4820 9976
rect 4724 9472 4820 9512
rect 4684 9463 4724 9472
rect 4396 9378 4436 9463
rect 4012 9136 4148 9176
rect 3284 8632 3860 8672
rect 3244 8623 3284 8632
rect 3436 8000 3476 8009
rect 3820 8000 3860 8632
rect 3476 7960 3572 8000
rect 3436 7951 3476 7960
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 3532 7412 3572 7960
rect 3532 7363 3572 7372
rect 3724 7960 3820 8000
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 3724 5648 3764 7960
rect 3820 7951 3860 7960
rect 4012 7220 4052 9136
rect 4107 8672 4149 8681
rect 4107 8632 4108 8672
rect 4148 8632 4149 8672
rect 4107 8623 4149 8632
rect 4779 8672 4821 8681
rect 4779 8632 4780 8672
rect 4820 8632 4821 8672
rect 4779 8623 4821 8632
rect 4108 8538 4148 8623
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4684 7866 4724 7951
rect 3916 7180 4052 7220
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 3916 7160 3956 7180
rect 3916 7111 3956 7120
rect 4204 7160 4244 7171
rect 3820 7026 3860 7111
rect 4204 7085 4244 7120
rect 4203 7076 4245 7085
rect 4203 7036 4204 7076
rect 4244 7036 4245 7076
rect 4203 7027 4245 7036
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3820 5648 3860 5657
rect 3724 5608 3820 5648
rect 3820 5599 3860 5608
rect 4684 5648 4724 5657
rect 4780 5648 4820 8623
rect 4876 8009 4916 10144
rect 4972 9521 5012 11395
rect 5836 11369 5876 11740
rect 5835 11360 5877 11369
rect 5835 11320 5836 11360
rect 5876 11320 5877 11360
rect 5835 11311 5877 11320
rect 5259 11108 5301 11117
rect 5259 11068 5260 11108
rect 5300 11068 5301 11108
rect 5259 11059 5301 11068
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 4875 8000 4917 8009
rect 4875 7960 4876 8000
rect 4916 7960 4917 8000
rect 4875 7951 4917 7960
rect 4875 7076 4917 7085
rect 4875 7036 4876 7076
rect 4916 7036 4917 7076
rect 4875 7027 4917 7036
rect 4724 5608 4820 5648
rect 4684 5599 4724 5608
rect 3436 5564 3476 5573
rect 3476 5524 3764 5564
rect 3436 5515 3476 5524
rect 3724 4976 3764 5524
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 4491 5060 4533 5069
rect 4491 5020 4492 5060
rect 4532 5020 4533 5060
rect 4491 5011 4533 5020
rect 3724 4936 4244 4976
rect 4204 4808 4244 4936
rect 4492 4926 4532 5011
rect 4588 4976 4628 4985
rect 4204 4759 4244 4768
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 2955 4220 2997 4229
rect 2955 4180 2956 4220
rect 2996 4180 2997 4220
rect 2955 4171 2997 4180
rect 4588 4145 4628 4936
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 2571 4052 2613 4061
rect 2571 4012 2572 4052
rect 2612 4012 2613 4052
rect 2571 4003 2613 4012
rect 2475 3884 2517 3893
rect 2475 3844 2476 3884
rect 2516 3844 2517 3884
rect 2475 3835 2517 3844
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 1995 3296 2037 3305
rect 1995 3256 1996 3296
rect 2036 3256 2037 3296
rect 1995 3247 2037 3256
rect 651 3128 693 3137
rect 651 3088 652 3128
rect 692 3088 693 3128
rect 651 3079 693 3088
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 4780 2885 4820 5608
rect 4876 4976 4916 7027
rect 4972 5741 5012 9463
rect 5260 8933 5300 11059
rect 5835 10940 5877 10949
rect 5835 10900 5836 10940
rect 5876 10900 5877 10940
rect 5835 10891 5877 10900
rect 5836 10436 5876 10891
rect 6028 10613 6068 17260
rect 6603 15560 6645 15569
rect 6603 15520 6604 15560
rect 6644 15520 6645 15560
rect 6603 15511 6645 15520
rect 6027 10604 6069 10613
rect 6027 10564 6028 10604
rect 6068 10564 6069 10604
rect 6027 10555 6069 10564
rect 5836 10387 5876 10396
rect 5259 8924 5301 8933
rect 5259 8884 5260 8924
rect 5300 8884 5301 8924
rect 5259 8875 5301 8884
rect 5260 8790 5300 8875
rect 5836 7748 5876 7757
rect 5876 7708 5972 7748
rect 5836 7699 5876 7708
rect 5932 7169 5972 7708
rect 5931 7160 5973 7169
rect 5931 7120 5932 7160
rect 5972 7120 5973 7160
rect 5931 7111 5973 7120
rect 4971 5732 5013 5741
rect 4971 5692 4972 5732
rect 5012 5692 5013 5732
rect 4971 5683 5013 5692
rect 5835 5732 5877 5741
rect 5835 5692 5836 5732
rect 5876 5692 5877 5732
rect 5835 5683 5877 5692
rect 4972 5069 5012 5683
rect 5836 5598 5876 5683
rect 5932 5405 5972 7111
rect 6604 5909 6644 15511
rect 6603 5900 6645 5909
rect 6603 5860 6604 5900
rect 6644 5860 6645 5900
rect 6603 5851 6645 5860
rect 5931 5396 5973 5405
rect 5931 5356 5932 5396
rect 5972 5356 5973 5396
rect 5931 5347 5973 5356
rect 4971 5060 5013 5069
rect 4971 5020 4972 5060
rect 5012 5020 5013 5060
rect 4971 5011 5013 5020
rect 4876 4927 4916 4936
rect 4779 2876 4821 2885
rect 4779 2836 4780 2876
rect 4820 2836 4821 2876
rect 4779 2827 4821 2836
rect 6892 2717 6932 31219
rect 7084 3473 7124 32815
rect 7276 32705 7316 32983
rect 8908 32864 8948 32873
rect 7275 32696 7317 32705
rect 7275 32656 7276 32696
rect 7316 32656 7317 32696
rect 7275 32647 7317 32656
rect 7756 32696 7796 32705
rect 7756 32453 7796 32656
rect 8908 32537 8948 32824
rect 9196 32864 9236 32873
rect 8907 32528 8949 32537
rect 8907 32488 8908 32528
rect 8948 32488 8949 32528
rect 8907 32479 8949 32488
rect 7755 32444 7797 32453
rect 7755 32404 7756 32444
rect 7796 32404 7797 32444
rect 7755 32395 7797 32404
rect 7947 32360 7989 32369
rect 7947 32320 7948 32360
rect 7988 32320 7989 32360
rect 7947 32311 7989 32320
rect 7851 31772 7893 31781
rect 7851 31732 7852 31772
rect 7892 31732 7893 31772
rect 7851 31723 7893 31732
rect 7659 15325 7701 15334
rect 7659 15285 7660 15325
rect 7700 15285 7701 15325
rect 7659 15276 7701 15285
rect 7660 14561 7700 15276
rect 7659 14552 7701 14561
rect 7659 14512 7660 14552
rect 7700 14512 7701 14552
rect 7659 14503 7701 14512
rect 7563 10772 7605 10781
rect 7563 10732 7564 10772
rect 7604 10732 7605 10772
rect 7563 10723 7605 10732
rect 7564 10193 7604 10723
rect 7563 10184 7605 10193
rect 7563 10144 7564 10184
rect 7604 10144 7605 10184
rect 7563 10135 7605 10144
rect 7660 5657 7700 14503
rect 7852 8681 7892 31723
rect 7851 8672 7893 8681
rect 7851 8632 7852 8672
rect 7892 8632 7893 8672
rect 7851 8623 7893 8632
rect 7659 5648 7701 5657
rect 7659 5608 7660 5648
rect 7700 5608 7701 5648
rect 7659 5599 7701 5608
rect 7948 5489 7988 32311
rect 9196 31865 9236 32824
rect 9292 32864 9332 33067
rect 9580 33032 9620 33041
rect 9620 32992 9908 33032
rect 9580 32983 9620 32992
rect 9292 32815 9332 32824
rect 9868 32864 9908 32992
rect 9868 32815 9908 32824
rect 10252 32864 10292 32873
rect 9195 31856 9237 31865
rect 9195 31816 9196 31856
rect 9236 31816 9237 31856
rect 9195 31807 9237 31816
rect 8235 31016 8277 31025
rect 8235 30976 8236 31016
rect 8276 30976 8277 31016
rect 8235 30967 8277 30976
rect 7947 5480 7989 5489
rect 7947 5440 7948 5480
rect 7988 5440 7989 5480
rect 7947 5431 7989 5440
rect 8236 3977 8276 30967
rect 10252 30269 10292 32824
rect 11116 32864 11156 33655
rect 13996 33125 14036 33664
rect 14380 33704 14420 34159
rect 14380 33655 14420 33664
rect 12267 33116 12309 33125
rect 12267 33076 12268 33116
rect 12308 33076 12309 33116
rect 12267 33067 12309 33076
rect 13995 33116 14037 33125
rect 13995 33076 13996 33116
rect 14036 33076 14037 33116
rect 13995 33067 14037 33076
rect 14475 33116 14517 33125
rect 14475 33076 14476 33116
rect 14516 33076 14517 33116
rect 14475 33067 14517 33076
rect 12268 32982 12308 33067
rect 14476 32982 14516 33067
rect 11116 31361 11156 32824
rect 13804 32864 13844 32873
rect 12267 32696 12309 32705
rect 12267 32656 12268 32696
rect 12308 32656 12309 32696
rect 12267 32647 12309 32656
rect 12268 32562 12308 32647
rect 13804 32537 13844 32824
rect 14092 32864 14132 32873
rect 14092 32705 14132 32824
rect 14188 32780 14228 32789
rect 14091 32696 14133 32705
rect 14091 32656 14092 32696
rect 14132 32656 14133 32696
rect 14091 32647 14133 32656
rect 14188 32621 14228 32740
rect 14187 32612 14229 32621
rect 14187 32572 14188 32612
rect 14228 32572 14229 32612
rect 14187 32563 14229 32572
rect 13803 32528 13845 32537
rect 13803 32488 13804 32528
rect 13844 32488 13845 32528
rect 13803 32479 13845 32488
rect 14668 31781 14708 34168
rect 14860 33629 14900 35092
rect 15052 35083 15092 35092
rect 32620 35057 32660 35176
rect 32716 35216 32756 35225
rect 33004 35216 33044 35225
rect 33772 35216 33812 35225
rect 32756 35176 32852 35216
rect 32716 35167 32756 35176
rect 32619 35048 32661 35057
rect 32619 35008 32620 35048
rect 32660 35008 32661 35048
rect 32619 34999 32661 35008
rect 15244 34964 15284 34973
rect 15051 34376 15093 34385
rect 15051 34336 15052 34376
rect 15092 34336 15093 34376
rect 15051 34327 15093 34336
rect 15052 34242 15092 34327
rect 15244 33881 15284 34924
rect 32332 34964 32372 34973
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 20811 34544 20853 34553
rect 20811 34504 20812 34544
rect 20852 34504 20853 34544
rect 20811 34495 20853 34504
rect 21579 34544 21621 34553
rect 21579 34504 21580 34544
rect 21620 34504 21621 34544
rect 21579 34495 21621 34504
rect 22731 34544 22773 34553
rect 22731 34504 22732 34544
rect 22772 34504 22773 34544
rect 22731 34495 22773 34504
rect 25323 34544 25365 34553
rect 25323 34504 25324 34544
rect 25364 34504 25365 34544
rect 25323 34495 25365 34504
rect 28972 34544 29012 34553
rect 29012 34504 29204 34544
rect 28972 34495 29012 34504
rect 20812 34460 20852 34495
rect 15820 34376 15860 34385
rect 15436 34292 15476 34301
rect 15340 34252 15436 34292
rect 15243 33872 15285 33881
rect 15243 33832 15244 33872
rect 15284 33832 15285 33872
rect 15243 33823 15285 33832
rect 15243 33704 15285 33713
rect 15243 33664 15244 33704
rect 15284 33664 15285 33704
rect 15243 33655 15285 33664
rect 14859 33620 14901 33629
rect 14859 33580 14860 33620
rect 14900 33580 14901 33620
rect 14859 33571 14901 33580
rect 14860 33377 14900 33571
rect 15244 33570 15284 33655
rect 14859 33368 14901 33377
rect 14859 33328 14860 33368
rect 14900 33328 14901 33368
rect 14859 33319 14901 33328
rect 15340 33116 15380 34252
rect 15436 34243 15476 34252
rect 15820 34217 15860 34336
rect 16684 34376 16724 34385
rect 16684 34217 16724 34336
rect 18412 34376 18452 34385
rect 19276 34376 19316 34385
rect 18452 34336 18740 34376
rect 18028 34292 18068 34301
rect 17932 34252 18028 34292
rect 15819 34208 15861 34217
rect 15819 34168 15820 34208
rect 15860 34168 15861 34208
rect 15819 34159 15861 34168
rect 16683 34208 16725 34217
rect 17836 34208 17876 34217
rect 16683 34168 16684 34208
rect 16724 34168 16725 34208
rect 16683 34159 16725 34168
rect 17452 34168 17836 34208
rect 16011 33872 16053 33881
rect 16011 33832 16012 33872
rect 16052 33832 16053 33872
rect 16011 33823 16053 33832
rect 16971 33872 17013 33881
rect 16971 33832 16972 33872
rect 17012 33832 17013 33872
rect 16971 33823 17013 33832
rect 15723 33788 15765 33797
rect 15723 33748 15724 33788
rect 15764 33748 15765 33788
rect 15723 33739 15765 33748
rect 15340 33067 15380 33076
rect 15724 32864 15764 33739
rect 15724 32815 15764 32824
rect 16012 32864 16052 33823
rect 16972 33704 17012 33823
rect 17355 33788 17397 33797
rect 17355 33748 17356 33788
rect 17396 33748 17397 33788
rect 17355 33739 17397 33748
rect 16972 33629 17012 33664
rect 17260 33662 17300 33671
rect 16971 33620 17013 33629
rect 16971 33580 16972 33620
rect 17012 33580 17013 33620
rect 16971 33571 17013 33580
rect 17356 33654 17396 33739
rect 16396 33452 16436 33461
rect 16396 33125 16436 33412
rect 16395 33116 16437 33125
rect 16395 33076 16396 33116
rect 16436 33076 16437 33116
rect 16395 33067 16437 33076
rect 16012 32815 16052 32824
rect 15628 32780 15668 32789
rect 15147 32696 15189 32705
rect 15147 32656 15148 32696
rect 15188 32656 15189 32696
rect 15147 32647 15189 32656
rect 14667 31772 14709 31781
rect 14667 31732 14668 31772
rect 14708 31732 14709 31772
rect 14667 31723 14709 31732
rect 11115 31352 11157 31361
rect 11115 31312 11116 31352
rect 11156 31312 11157 31352
rect 11115 31303 11157 31312
rect 15148 30344 15188 32647
rect 15628 32285 15668 32740
rect 16396 32621 16436 33067
rect 16972 32948 17012 33571
rect 17260 33125 17300 33622
rect 17259 33116 17301 33125
rect 17259 33076 17260 33116
rect 17300 33076 17301 33116
rect 17259 33067 17301 33076
rect 16972 32908 17256 32948
rect 17216 32864 17256 32908
rect 17216 32815 17256 32824
rect 16395 32612 16437 32621
rect 16395 32572 16396 32612
rect 16436 32572 16437 32612
rect 16395 32563 16437 32572
rect 16299 32528 16341 32537
rect 16299 32488 16300 32528
rect 16340 32488 16341 32528
rect 16299 32479 16341 32488
rect 15627 32276 15669 32285
rect 15627 32236 15628 32276
rect 15668 32236 15669 32276
rect 15627 32227 15669 32236
rect 16300 30344 16340 32479
rect 17452 32285 17492 34168
rect 17836 34159 17876 34168
rect 17932 33704 17972 34252
rect 18028 34243 18068 34252
rect 18412 34133 18452 34336
rect 18411 34124 18453 34133
rect 18411 34084 18412 34124
rect 18452 34084 18453 34124
rect 18411 34075 18453 34084
rect 17740 33664 17972 33704
rect 17644 33536 17684 33545
rect 17740 33536 17780 33664
rect 17684 33496 17780 33536
rect 17644 33487 17684 33496
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 17643 33116 17685 33125
rect 17643 33076 17644 33116
rect 17684 33076 17685 33116
rect 17643 33067 17685 33076
rect 17548 32864 17588 32873
rect 17548 32537 17588 32824
rect 17644 32864 17684 33067
rect 17932 33032 17972 33041
rect 17972 32992 18164 33032
rect 17932 32983 17972 32992
rect 17644 32815 17684 32824
rect 18124 32864 18164 32992
rect 18124 32815 18164 32824
rect 18508 32864 18548 32873
rect 18700 32864 18740 34336
rect 19276 34217 19316 34336
rect 19275 34208 19317 34217
rect 19275 34168 19276 34208
rect 19316 34168 19317 34208
rect 19275 34159 19317 34168
rect 20428 34208 20468 34217
rect 19276 33452 19316 34159
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 20428 33797 20468 34168
rect 20427 33788 20469 33797
rect 20427 33748 20428 33788
rect 20468 33748 20469 33788
rect 20427 33739 20469 33748
rect 20428 33545 20468 33739
rect 20716 33704 20756 33713
rect 20619 33620 20661 33629
rect 20716 33620 20756 33664
rect 20619 33580 20620 33620
rect 20660 33580 20756 33620
rect 20619 33571 20661 33580
rect 20427 33536 20469 33545
rect 20427 33496 20428 33536
rect 20468 33496 20469 33536
rect 20427 33487 20469 33496
rect 19371 33452 19413 33461
rect 19276 33412 19372 33452
rect 19412 33412 19413 33452
rect 19371 33403 19413 33412
rect 19275 33116 19317 33125
rect 19275 33076 19276 33116
rect 19316 33076 19317 33116
rect 19275 33067 19317 33076
rect 18548 32824 18740 32864
rect 18508 32815 18548 32824
rect 18795 32696 18837 32705
rect 18795 32656 18796 32696
rect 18836 32656 18837 32696
rect 18795 32647 18837 32656
rect 17547 32528 17589 32537
rect 17547 32488 17548 32528
rect 17588 32488 17589 32528
rect 17547 32479 17589 32488
rect 17451 32276 17493 32285
rect 17451 32236 17452 32276
rect 17492 32236 17493 32276
rect 17451 32227 17493 32236
rect 18027 32276 18069 32285
rect 18027 32236 18028 32276
rect 18068 32236 18069 32276
rect 18027 32227 18069 32236
rect 18028 30344 18068 32227
rect 18796 30344 18836 32647
rect 19276 30344 19316 33067
rect 19372 32864 19412 33403
rect 20523 33116 20565 33125
rect 20523 33076 20524 33116
rect 20564 33076 20565 33116
rect 20523 33067 20565 33076
rect 20524 32982 20564 33067
rect 19372 32815 19412 32824
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 20812 31949 20852 34420
rect 21196 34460 21236 34469
rect 21004 34208 21044 34217
rect 21196 34208 21236 34420
rect 21580 34460 21620 34495
rect 21580 34409 21620 34420
rect 22732 34410 22772 34495
rect 22924 34460 22964 34469
rect 22828 34420 22924 34460
rect 22060 34376 22100 34385
rect 22060 34217 22100 34336
rect 22347 34376 22389 34385
rect 22347 34336 22348 34376
rect 22388 34336 22389 34376
rect 22347 34327 22389 34336
rect 21044 34168 21236 34208
rect 21004 34159 21044 34168
rect 21099 33788 21141 33797
rect 21099 33748 21100 33788
rect 21140 33748 21141 33788
rect 21099 33739 21141 33748
rect 21004 33704 21044 33713
rect 21004 33125 21044 33664
rect 21100 33654 21140 33739
rect 21196 33629 21236 34168
rect 21388 34208 21428 34217
rect 21388 33881 21428 34168
rect 21772 34208 21812 34217
rect 22059 34208 22101 34217
rect 21812 34168 22060 34208
rect 22100 34168 22101 34208
rect 21772 34159 21812 34168
rect 22059 34159 22101 34168
rect 21771 34040 21813 34049
rect 21771 34000 21772 34040
rect 21812 34000 21813 34040
rect 21771 33991 21813 34000
rect 21387 33872 21429 33881
rect 21387 33832 21388 33872
rect 21428 33832 21429 33872
rect 21387 33823 21429 33832
rect 21579 33872 21621 33881
rect 21579 33832 21580 33872
rect 21620 33832 21621 33872
rect 21579 33823 21621 33832
rect 21195 33620 21237 33629
rect 21195 33580 21196 33620
rect 21236 33580 21237 33620
rect 21195 33571 21237 33580
rect 21003 33116 21045 33125
rect 21003 33076 21004 33116
rect 21044 33076 21045 33116
rect 21003 33067 21045 33076
rect 20811 31940 20853 31949
rect 20811 31900 20812 31940
rect 20852 31900 20853 31940
rect 20811 31891 20853 31900
rect 21196 31277 21236 33571
rect 21388 33452 21428 33461
rect 21292 32864 21332 32873
rect 21388 32864 21428 33412
rect 21332 32824 21428 32864
rect 21580 32864 21620 33823
rect 21772 33704 21812 33991
rect 22348 33797 22388 34327
rect 22444 34292 22484 34301
rect 22347 33788 22389 33797
rect 22347 33748 22348 33788
rect 22388 33748 22389 33788
rect 22347 33739 22389 33748
rect 21772 33655 21812 33664
rect 22444 33461 22484 34252
rect 22635 33788 22677 33797
rect 22635 33748 22636 33788
rect 22676 33748 22677 33788
rect 22635 33739 22677 33748
rect 22636 33704 22676 33739
rect 21963 33452 22005 33461
rect 21963 33412 21964 33452
rect 22004 33412 22005 33452
rect 21963 33403 22005 33412
rect 22443 33452 22485 33461
rect 22443 33412 22444 33452
rect 22484 33412 22485 33452
rect 22443 33403 22485 33412
rect 21964 33318 22004 33403
rect 21676 32864 21716 32873
rect 21580 32824 21676 32864
rect 21292 32815 21332 32824
rect 21676 32815 21716 32824
rect 22540 32864 22580 32873
rect 22636 32864 22676 33664
rect 22828 33377 22868 34420
rect 22924 34411 22964 34420
rect 23115 34460 23157 34469
rect 23115 34420 23116 34460
rect 23156 34420 23157 34460
rect 23115 34411 23157 34420
rect 23116 34208 23156 34411
rect 23691 34376 23733 34385
rect 23691 34336 23692 34376
rect 23732 34336 23733 34376
rect 23691 34327 23733 34336
rect 23019 33620 23061 33629
rect 23019 33580 23020 33620
rect 23060 33580 23061 33620
rect 23019 33571 23061 33580
rect 22923 33452 22965 33461
rect 22923 33412 22924 33452
rect 22964 33412 22965 33452
rect 22923 33403 22965 33412
rect 22827 33368 22869 33377
rect 22827 33328 22828 33368
rect 22868 33328 22869 33368
rect 22827 33319 22869 33328
rect 22924 33318 22964 33403
rect 22580 32824 22676 32864
rect 22540 32815 22580 32824
rect 23020 32453 23060 33571
rect 23019 32444 23061 32453
rect 23019 32404 23020 32444
rect 23060 32404 23061 32444
rect 23019 32395 23061 32404
rect 21195 31268 21237 31277
rect 21195 31228 21196 31268
rect 21236 31228 21237 31268
rect 21195 31219 21237 31228
rect 23116 31025 23156 34168
rect 23692 33116 23732 34327
rect 24939 33872 24981 33881
rect 24939 33832 24940 33872
rect 24980 33832 24981 33872
rect 24939 33823 24981 33832
rect 24075 33788 24117 33797
rect 24075 33748 24076 33788
rect 24116 33748 24117 33788
rect 24075 33739 24117 33748
rect 24076 33704 24116 33739
rect 24076 33653 24116 33664
rect 24940 33704 24980 33823
rect 25324 33788 25364 34495
rect 25803 34460 25845 34469
rect 25803 34420 25804 34460
rect 25844 34420 25845 34460
rect 25803 34411 25845 34420
rect 25804 34133 25844 34411
rect 27819 34208 27861 34217
rect 27819 34168 27820 34208
rect 27860 34168 27861 34208
rect 27819 34159 27861 34168
rect 25803 34124 25845 34133
rect 25803 34084 25804 34124
rect 25844 34084 25845 34124
rect 25803 34075 25845 34084
rect 25611 34040 25653 34049
rect 25611 34000 25612 34040
rect 25652 34000 25653 34040
rect 25611 33991 25653 34000
rect 25324 33739 25364 33748
rect 24940 33655 24980 33664
rect 25612 33704 25652 33991
rect 27531 33872 27573 33881
rect 27531 33832 27532 33872
rect 27572 33832 27573 33872
rect 27531 33823 27573 33832
rect 26572 33704 26612 33713
rect 25652 33664 25748 33704
rect 25612 33655 25652 33664
rect 23979 33536 24021 33545
rect 23979 33496 23980 33536
rect 24020 33496 24021 33536
rect 23979 33487 24021 33496
rect 23692 33067 23732 33076
rect 23692 32696 23732 32705
rect 23115 31016 23157 31025
rect 23115 30976 23116 31016
rect 23156 30976 23157 31016
rect 23115 30967 23157 30976
rect 23692 30344 23732 32656
rect 23980 30344 24020 33487
rect 25515 33452 25557 33461
rect 25515 33412 25516 33452
rect 25556 33412 25557 33452
rect 25515 33403 25557 33412
rect 25516 32864 25556 33403
rect 25516 32815 25556 32824
rect 25708 32705 25748 33664
rect 26572 33461 26612 33664
rect 27148 33704 27188 33713
rect 26571 33452 26613 33461
rect 26571 33412 26572 33452
rect 26612 33412 26613 33452
rect 26571 33403 26613 33412
rect 27148 33116 27188 33664
rect 27532 33704 27572 33823
rect 27532 33209 27572 33664
rect 27531 33200 27573 33209
rect 27531 33160 27532 33200
rect 27572 33160 27573 33200
rect 27531 33151 27573 33160
rect 27148 33067 27188 33076
rect 27532 32864 27572 32873
rect 27436 32780 27476 32789
rect 25707 32696 25749 32705
rect 25707 32656 25708 32696
rect 25748 32656 25749 32696
rect 25707 32647 25749 32656
rect 27436 32537 27476 32740
rect 27435 32528 27477 32537
rect 27435 32488 27436 32528
rect 27476 32488 27477 32528
rect 27435 32479 27477 32488
rect 27532 31193 27572 32824
rect 27820 32864 27860 34159
rect 28395 33704 28437 33713
rect 28395 33664 28396 33704
rect 28436 33664 28437 33704
rect 28395 33655 28437 33664
rect 28396 33570 28436 33655
rect 29164 32864 29204 34504
rect 29356 34376 29396 34385
rect 29260 34292 29300 34301
rect 29260 33545 29300 34252
rect 29356 33872 29396 34336
rect 29644 34376 29684 34385
rect 29644 34217 29684 34336
rect 31467 34376 31509 34385
rect 31467 34336 31468 34376
rect 31508 34336 31509 34376
rect 31467 34327 31509 34336
rect 32332 34376 32372 34924
rect 32332 34327 32372 34336
rect 32715 34376 32757 34385
rect 32715 34336 32716 34376
rect 32756 34336 32757 34376
rect 32715 34327 32757 34336
rect 29643 34208 29685 34217
rect 29643 34168 29644 34208
rect 29684 34168 29685 34208
rect 29643 34159 29685 34168
rect 29644 33965 29684 34159
rect 29643 33956 29685 33965
rect 29643 33916 29644 33956
rect 29684 33916 29685 33956
rect 29643 33907 29685 33916
rect 30219 33956 30261 33965
rect 30219 33916 30220 33956
rect 30260 33916 30261 33956
rect 30219 33907 30261 33916
rect 29548 33872 29588 33881
rect 29356 33832 29548 33872
rect 29548 33823 29588 33832
rect 30220 33704 30260 33907
rect 30220 33655 30260 33664
rect 30508 33704 30548 33713
rect 30508 33545 30548 33664
rect 30603 33704 30645 33713
rect 30603 33664 30604 33704
rect 30644 33664 30645 33704
rect 30603 33655 30645 33664
rect 31084 33704 31124 33713
rect 30604 33570 30644 33655
rect 29259 33536 29301 33545
rect 29259 33496 29260 33536
rect 29300 33496 29301 33536
rect 29259 33487 29301 33496
rect 30507 33536 30549 33545
rect 30507 33496 30508 33536
rect 30548 33496 30549 33536
rect 30507 33487 30549 33496
rect 30892 33536 30932 33545
rect 31084 33536 31124 33664
rect 30932 33496 31124 33536
rect 31468 33704 31508 34327
rect 32716 34242 32756 34327
rect 32812 34217 32852 35176
rect 33044 35176 33140 35216
rect 33004 35167 33044 35176
rect 33003 35048 33045 35057
rect 33003 35008 33004 35048
rect 33044 35008 33045 35048
rect 33003 34999 33045 35008
rect 32811 34208 32853 34217
rect 32811 34168 32812 34208
rect 32852 34168 32853 34208
rect 32811 34159 32853 34168
rect 30892 33487 30932 33496
rect 29548 33452 29588 33461
rect 30603 33452 30645 33461
rect 29588 33412 29684 33452
rect 29548 33403 29588 33412
rect 29356 32864 29396 32873
rect 29164 32824 29356 32864
rect 27820 32815 27860 32824
rect 29356 32815 29396 32824
rect 29644 32537 29684 33412
rect 30603 33412 30604 33452
rect 30644 33412 30645 33452
rect 30603 33403 30645 33412
rect 30219 33368 30261 33377
rect 30219 33328 30220 33368
rect 30260 33328 30261 33368
rect 30219 33319 30261 33328
rect 29739 33200 29781 33209
rect 29739 33160 29740 33200
rect 29780 33160 29781 33200
rect 29739 33151 29781 33160
rect 29740 32864 29780 33151
rect 29740 32815 29780 32824
rect 29643 32528 29685 32537
rect 29643 32488 29644 32528
rect 29684 32488 29685 32528
rect 29643 32479 29685 32488
rect 27531 31184 27573 31193
rect 27531 31144 27532 31184
rect 27572 31144 27573 31184
rect 27531 31135 27573 31144
rect 29547 31184 29589 31193
rect 29547 31144 29548 31184
rect 29588 31144 29589 31184
rect 29547 31135 29589 31144
rect 29548 30344 29588 31135
rect 29644 30344 29684 32479
rect 30220 30344 30260 33319
rect 30604 32864 30644 33403
rect 31468 33209 31508 33664
rect 31563 33704 31605 33713
rect 31563 33664 31564 33704
rect 31604 33664 31605 33704
rect 31563 33655 31605 33664
rect 32332 33704 32372 33713
rect 31467 33200 31509 33209
rect 31467 33160 31468 33200
rect 31508 33160 31509 33200
rect 31467 33151 31509 33160
rect 30604 32815 30644 32824
rect 31564 30344 31604 33655
rect 31755 33536 31797 33545
rect 31755 33496 31756 33536
rect 31796 33496 31797 33536
rect 31755 33487 31797 33496
rect 31756 33116 31796 33487
rect 32332 33461 32372 33664
rect 32331 33452 32373 33461
rect 32331 33412 32332 33452
rect 32372 33412 32373 33452
rect 32331 33403 32373 33412
rect 31756 33067 31796 33076
rect 15148 30304 15201 30344
rect 16300 30304 16353 30344
rect 18028 30304 18081 30344
rect 18796 30304 18849 30344
rect 19276 30304 19617 30344
rect 23692 30304 23841 30344
rect 23980 30304 24033 30344
rect 29548 30304 29601 30344
rect 29644 30304 29793 30344
rect 10251 30260 10293 30269
rect 10251 30220 10252 30260
rect 10292 30220 10293 30260
rect 10251 30211 10293 30220
rect 15161 29960 15201 30304
rect 16313 29960 16353 30304
rect 18041 29960 18081 30304
rect 18232 30092 18274 30101
rect 18232 30052 18233 30092
rect 18273 30052 18274 30092
rect 18232 30043 18274 30052
rect 18233 29960 18273 30043
rect 18809 29960 18849 30304
rect 19577 29960 19617 30304
rect 23801 29960 23841 30304
rect 23993 29960 24033 30304
rect 29561 29960 29601 30304
rect 29753 29960 29793 30304
rect 30172 30304 30260 30344
rect 31516 30304 31604 30344
rect 31756 32696 31796 32705
rect 31756 30344 31796 32656
rect 32812 30344 32852 34159
rect 33004 30344 33044 34999
rect 33100 33965 33140 35176
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 33580 34376 33620 34385
rect 33099 33956 33141 33965
rect 33099 33916 33100 33956
rect 33140 33916 33141 33956
rect 33099 33907 33141 33916
rect 33483 33704 33525 33713
rect 33483 33664 33484 33704
rect 33524 33664 33525 33704
rect 33483 33655 33525 33664
rect 33484 33620 33524 33655
rect 33484 33569 33524 33580
rect 33580 33461 33620 34336
rect 33772 34133 33812 35176
rect 34060 35216 34100 35225
rect 34060 35057 34100 35176
rect 34156 35216 34196 35225
rect 50284 35216 50324 35225
rect 34196 35176 34292 35216
rect 34156 35167 34196 35176
rect 34059 35048 34101 35057
rect 34059 35008 34060 35048
rect 34100 35008 34101 35048
rect 34059 34999 34101 35008
rect 33771 34124 33813 34133
rect 33771 34084 33772 34124
rect 33812 34084 33813 34124
rect 33771 34075 33813 34084
rect 33771 33956 33813 33965
rect 33771 33916 33772 33956
rect 33812 33916 33813 33956
rect 33771 33907 33813 33916
rect 33772 33704 33812 33907
rect 34156 33797 34196 33828
rect 34155 33788 34197 33797
rect 34155 33748 34156 33788
rect 34196 33748 34197 33788
rect 34155 33739 34197 33748
rect 33772 33655 33812 33664
rect 34059 33704 34101 33713
rect 34059 33664 34060 33704
rect 34100 33664 34101 33704
rect 34059 33655 34101 33664
rect 34156 33704 34196 33739
rect 34060 33570 34100 33655
rect 33579 33452 33621 33461
rect 33579 33412 33580 33452
rect 33620 33412 33621 33452
rect 33579 33403 33621 33412
rect 34156 33377 34196 33664
rect 34155 33368 34197 33377
rect 34155 33328 34156 33368
rect 34196 33328 34197 33368
rect 34155 33319 34197 33328
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 34252 33125 34292 35176
rect 34731 35048 34773 35057
rect 34731 35008 34732 35048
rect 34772 35008 34773 35048
rect 34731 34999 34773 35008
rect 34444 34964 34484 34973
rect 34348 34924 34444 34964
rect 34251 33116 34293 33125
rect 34251 33076 34252 33116
rect 34292 33076 34293 33116
rect 34251 33067 34293 33076
rect 33099 33032 33141 33041
rect 33099 32992 33100 33032
rect 33140 32992 33141 33032
rect 33099 32983 33141 32992
rect 33100 32864 33140 32983
rect 33100 32815 33140 32824
rect 33964 32864 34004 32873
rect 33964 32705 34004 32824
rect 33963 32696 34005 32705
rect 33963 32656 33964 32696
rect 34004 32656 34005 32696
rect 33963 32647 34005 32656
rect 34252 32369 34292 33067
rect 34348 32864 34388 34924
rect 34444 34915 34484 34924
rect 34732 34544 34772 34999
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 34732 34495 34772 34504
rect 38188 34544 38228 34553
rect 35691 34376 35733 34385
rect 35691 34336 35692 34376
rect 35732 34336 35733 34376
rect 35691 34327 35733 34336
rect 36940 34376 36980 34385
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 35692 33713 35732 34327
rect 34443 33704 34485 33713
rect 34443 33664 34444 33704
rect 34484 33664 34485 33704
rect 34443 33655 34485 33664
rect 35307 33704 35349 33713
rect 35307 33664 35308 33704
rect 35348 33664 35349 33704
rect 35307 33655 35349 33664
rect 35691 33704 35733 33713
rect 35691 33664 35692 33704
rect 35732 33664 35733 33704
rect 35691 33655 35733 33664
rect 36556 33704 36596 33713
rect 34444 33536 34484 33655
rect 35308 33570 35348 33655
rect 35692 33570 35732 33655
rect 34444 33487 34484 33496
rect 36556 33461 36596 33664
rect 36940 33629 36980 34336
rect 37900 34376 37940 34385
rect 37940 34336 38132 34376
rect 37900 34327 37940 34336
rect 37899 34208 37941 34217
rect 37899 34168 37900 34208
rect 37940 34168 37941 34208
rect 37899 34159 37941 34168
rect 37707 33788 37749 33797
rect 37707 33748 37708 33788
rect 37748 33748 37749 33788
rect 37707 33739 37749 33748
rect 37900 33788 37940 34159
rect 37900 33739 37940 33748
rect 36939 33620 36981 33629
rect 36939 33580 36940 33620
rect 36980 33580 36981 33620
rect 36939 33571 36981 33580
rect 35595 33452 35637 33461
rect 35595 33412 35596 33452
rect 35636 33412 35637 33452
rect 35595 33403 35637 33412
rect 36555 33452 36597 33461
rect 36555 33412 36556 33452
rect 36596 33412 36597 33452
rect 36555 33403 36597 33412
rect 34348 32815 34388 32824
rect 34732 32864 34772 32873
rect 34732 32696 34772 32824
rect 35596 32864 35636 33403
rect 36747 33116 36789 33125
rect 36747 33076 36748 33116
rect 36788 33076 36789 33116
rect 36747 33067 36789 33076
rect 36748 32982 36788 33067
rect 35596 32815 35636 32824
rect 36940 32864 36980 33571
rect 37708 33461 37748 33739
rect 37707 33452 37749 33461
rect 37707 33412 37708 33452
rect 37748 33412 37749 33452
rect 37707 33403 37749 33412
rect 37708 33318 37748 33403
rect 36940 32815 36980 32824
rect 37323 32864 37365 32873
rect 37323 32824 37324 32864
rect 37364 32824 37365 32864
rect 37323 32815 37365 32824
rect 37324 32730 37364 32815
rect 38092 32705 38132 34336
rect 38188 34217 38228 34504
rect 49995 34544 50037 34553
rect 49995 34504 49996 34544
rect 50036 34504 50037 34544
rect 50284 34544 50324 35176
rect 82252 35132 82292 35141
rect 81195 34964 81237 34973
rect 81195 34924 81196 34964
rect 81236 34924 81237 34964
rect 81195 34915 81237 34924
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 50572 34544 50612 34553
rect 50284 34504 50572 34544
rect 49995 34495 50037 34504
rect 50572 34495 50612 34504
rect 52204 34544 52244 34553
rect 42123 34460 42165 34469
rect 45580 34460 45620 34469
rect 42123 34420 42124 34460
rect 42164 34420 42165 34460
rect 42123 34411 42165 34420
rect 45484 34420 45580 34460
rect 38572 34376 38612 34385
rect 38476 34292 38516 34301
rect 38187 34208 38229 34217
rect 38187 34168 38188 34208
rect 38228 34168 38229 34208
rect 38187 34159 38229 34168
rect 38476 34133 38516 34252
rect 38475 34124 38517 34133
rect 38475 34084 38476 34124
rect 38516 34084 38517 34124
rect 38475 34075 38517 34084
rect 38476 33881 38516 34075
rect 38475 33872 38517 33881
rect 38475 33832 38476 33872
rect 38516 33832 38517 33872
rect 38475 33823 38517 33832
rect 38283 33704 38325 33713
rect 38283 33664 38284 33704
rect 38324 33664 38325 33704
rect 38283 33655 38325 33664
rect 38284 33570 38324 33655
rect 38572 33209 38612 34336
rect 38859 34376 38901 34385
rect 38859 34336 38860 34376
rect 38900 34336 38901 34376
rect 38859 34327 38901 34336
rect 40587 34376 40629 34385
rect 40587 34336 40588 34376
rect 40628 34336 40629 34376
rect 40587 34327 40629 34336
rect 38860 33965 38900 34327
rect 38859 33956 38901 33965
rect 38859 33916 38860 33956
rect 38900 33916 38901 33956
rect 38859 33907 38901 33916
rect 40299 33872 40341 33881
rect 40299 33832 40300 33872
rect 40340 33832 40341 33872
rect 40299 33823 40341 33832
rect 40300 33738 40340 33823
rect 39147 33704 39189 33713
rect 39147 33664 39148 33704
rect 39188 33664 39189 33704
rect 39147 33655 39189 33664
rect 39148 33570 39188 33655
rect 38571 33200 38613 33209
rect 38571 33160 38572 33200
rect 38612 33160 38613 33200
rect 38571 33151 38613 33160
rect 38764 32864 38804 32873
rect 34444 32656 34772 32696
rect 38091 32696 38133 32705
rect 38091 32656 38092 32696
rect 38132 32656 38133 32696
rect 34444 32453 34484 32656
rect 38091 32647 38133 32656
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 34443 32444 34485 32453
rect 34443 32404 34444 32444
rect 34484 32404 34485 32444
rect 34443 32395 34485 32404
rect 34251 32360 34293 32369
rect 34251 32320 34252 32360
rect 34292 32320 34293 32360
rect 34251 32311 34293 32320
rect 38764 30941 38804 32824
rect 40588 32864 40628 34327
rect 42124 33881 42164 34411
rect 45388 34208 45428 34217
rect 42123 33872 42165 33881
rect 42123 33832 42124 33872
rect 42164 33832 42165 33872
rect 42123 33823 42165 33832
rect 41644 33704 41684 33713
rect 40875 33452 40917 33461
rect 40875 33412 40876 33452
rect 40916 33412 40917 33452
rect 40875 33403 40917 33412
rect 40588 32815 40628 32824
rect 40876 32864 40916 33403
rect 41260 33116 41300 33125
rect 41644 33116 41684 33664
rect 42028 33704 42068 33715
rect 42028 33629 42068 33664
rect 42027 33620 42069 33629
rect 42027 33580 42028 33620
rect 42068 33580 42069 33620
rect 42027 33571 42069 33580
rect 41300 33076 41684 33116
rect 41260 33067 41300 33076
rect 42124 32948 42164 33823
rect 42891 33704 42933 33713
rect 42891 33664 42892 33704
rect 42932 33664 42933 33704
rect 42891 33655 42933 33664
rect 44908 33704 44948 33713
rect 42315 33620 42357 33629
rect 42315 33580 42316 33620
rect 42356 33580 42357 33620
rect 42315 33571 42357 33580
rect 42316 33116 42356 33571
rect 42892 33570 42932 33655
rect 42316 33067 42356 33076
rect 44044 33452 44084 33461
rect 43083 33032 43125 33041
rect 43083 32992 43084 33032
rect 43124 32992 43125 33032
rect 43083 32983 43125 32992
rect 42124 32899 42164 32908
rect 43084 32898 43124 32983
rect 44044 32873 44084 33412
rect 44908 33140 44948 33664
rect 45292 33704 45332 33715
rect 45292 33629 45332 33664
rect 45291 33620 45333 33629
rect 45291 33580 45292 33620
rect 45332 33580 45333 33620
rect 45291 33571 45333 33580
rect 44908 33116 45332 33140
rect 44908 33100 45292 33116
rect 45292 33067 45332 33076
rect 40876 32815 40916 32824
rect 40971 32864 41013 32873
rect 40971 32824 40972 32864
rect 41012 32824 41013 32864
rect 40971 32815 41013 32824
rect 44043 32864 44085 32873
rect 44043 32824 44044 32864
rect 44084 32824 44085 32864
rect 44043 32815 44085 32824
rect 44715 32864 44757 32873
rect 44715 32824 44716 32864
rect 44756 32824 44757 32864
rect 44715 32815 44757 32824
rect 40972 32730 41012 32815
rect 42699 32696 42741 32705
rect 42699 32656 42700 32696
rect 42740 32656 42741 32696
rect 42699 32647 42741 32656
rect 42700 32562 42740 32647
rect 44044 32537 44084 32815
rect 44716 32730 44756 32815
rect 45388 32705 45428 34168
rect 45387 32696 45429 32705
rect 45387 32656 45388 32696
rect 45428 32656 45429 32696
rect 45387 32647 45429 32656
rect 44043 32528 44085 32537
rect 44043 32488 44044 32528
rect 44084 32488 44085 32528
rect 44043 32479 44085 32488
rect 45484 31277 45524 34420
rect 45580 34411 45620 34420
rect 49996 34410 50036 34495
rect 51820 34385 51860 34470
rect 49323 34376 49365 34385
rect 49323 34336 49324 34376
rect 49364 34336 49365 34376
rect 49323 34327 49365 34336
rect 49612 34376 49652 34385
rect 49324 34242 49364 34327
rect 46156 33704 46196 33713
rect 45579 33200 45621 33209
rect 45579 33160 45580 33200
rect 45620 33160 45621 33200
rect 45579 33151 45621 33160
rect 45580 32864 45620 33151
rect 45580 32815 45620 32824
rect 45676 32864 45716 32873
rect 45676 32621 45716 32824
rect 45964 32864 46004 32873
rect 45964 32705 46004 32824
rect 46156 32705 46196 33664
rect 47500 33704 47540 33713
rect 47308 33452 47348 33461
rect 47308 33293 47348 33412
rect 47307 33284 47349 33293
rect 47307 33244 47308 33284
rect 47348 33244 47349 33284
rect 47307 33235 47349 33244
rect 47500 33140 47540 33664
rect 47884 33704 47924 33715
rect 47884 33629 47924 33664
rect 48747 33704 48789 33713
rect 48747 33664 48748 33704
rect 48788 33664 48789 33704
rect 48747 33655 48789 33664
rect 47883 33620 47925 33629
rect 47883 33580 47884 33620
rect 47924 33580 47925 33620
rect 47883 33571 47925 33580
rect 48748 33570 48788 33655
rect 49612 33536 49652 34336
rect 50284 34376 50324 34385
rect 49707 34292 49749 34301
rect 49707 34252 49708 34292
rect 49748 34252 49749 34292
rect 49707 34243 49749 34252
rect 49708 34158 49748 34243
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 50091 33788 50133 33797
rect 50091 33748 50092 33788
rect 50132 33748 50133 33788
rect 50091 33739 50133 33748
rect 50092 33654 50132 33739
rect 48940 33496 49652 33536
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 47979 33200 48021 33209
rect 47979 33160 47980 33200
rect 48020 33160 48021 33200
rect 47979 33151 48021 33160
rect 47212 33116 47540 33140
rect 47252 33100 47540 33116
rect 47212 33067 47252 33076
rect 47596 32864 47636 32873
rect 47500 32780 47540 32789
rect 45963 32696 46005 32705
rect 45963 32656 45964 32696
rect 46004 32656 46005 32696
rect 45963 32647 46005 32656
rect 46155 32696 46197 32705
rect 46155 32656 46156 32696
rect 46196 32656 46197 32696
rect 46155 32647 46197 32656
rect 45675 32612 45717 32621
rect 45675 32572 45676 32612
rect 45716 32572 45717 32612
rect 45675 32563 45717 32572
rect 45964 32285 46004 32647
rect 47500 32621 47540 32740
rect 47499 32612 47541 32621
rect 47499 32572 47500 32612
rect 47540 32572 47541 32612
rect 47499 32563 47541 32572
rect 47596 32453 47636 32824
rect 47884 32864 47924 32873
rect 47595 32444 47637 32453
rect 47595 32404 47596 32444
rect 47636 32404 47637 32444
rect 47595 32395 47637 32404
rect 47884 32285 47924 32824
rect 45963 32276 46005 32285
rect 45963 32236 45964 32276
rect 46004 32236 46005 32276
rect 45963 32227 46005 32236
rect 47883 32276 47925 32285
rect 47883 32236 47884 32276
rect 47924 32236 47925 32276
rect 47883 32227 47925 32236
rect 45483 31268 45525 31277
rect 45483 31228 45484 31268
rect 45524 31228 45525 31268
rect 45483 31219 45525 31228
rect 38763 30932 38805 30941
rect 38763 30892 38764 30932
rect 38804 30892 38805 30932
rect 38763 30883 38805 30892
rect 47980 30344 48020 33151
rect 48652 32696 48692 32705
rect 48652 31109 48692 32656
rect 48940 32537 48980 33496
rect 49900 33452 49940 33461
rect 49324 33412 49900 33452
rect 49131 33032 49173 33041
rect 49131 32992 49132 33032
rect 49172 32992 49173 33032
rect 49131 32983 49173 32992
rect 49132 32864 49172 32983
rect 49132 32815 49172 32824
rect 49324 32621 49364 33412
rect 49900 33403 49940 33412
rect 50284 33041 50324 34336
rect 51531 34376 51573 34385
rect 51531 34336 51532 34376
rect 51572 34336 51573 34376
rect 51531 34327 51573 34336
rect 51819 34376 51861 34385
rect 51819 34336 51820 34376
rect 51860 34336 51861 34376
rect 51819 34327 51861 34336
rect 50764 34208 50804 34217
rect 50476 33704 50516 33715
rect 50764 33713 50804 34168
rect 50476 33629 50516 33664
rect 50763 33704 50805 33713
rect 50763 33664 50764 33704
rect 50804 33664 50805 33704
rect 50763 33655 50805 33664
rect 51339 33704 51381 33713
rect 51339 33664 51340 33704
rect 51380 33664 51381 33704
rect 51339 33655 51381 33664
rect 50475 33620 50517 33629
rect 50475 33580 50476 33620
rect 50516 33580 50612 33620
rect 50475 33571 50517 33580
rect 50283 33032 50325 33041
rect 50283 32992 50284 33032
rect 50324 32992 50325 33032
rect 50283 32983 50325 32992
rect 50284 32864 50324 32983
rect 50284 32815 50324 32824
rect 49900 32705 49940 32790
rect 49899 32696 49941 32705
rect 49899 32656 49900 32696
rect 49940 32656 49941 32696
rect 49899 32647 49941 32656
rect 50572 32621 50612 33580
rect 51340 33570 51380 33655
rect 50763 33032 50805 33041
rect 50763 32992 50764 33032
rect 50804 32992 50805 33032
rect 50763 32983 50805 32992
rect 50764 32864 50804 32983
rect 50764 32815 50804 32824
rect 49323 32612 49365 32621
rect 49323 32572 49324 32612
rect 49364 32572 49365 32612
rect 49323 32563 49365 32572
rect 50571 32612 50613 32621
rect 50571 32572 50572 32612
rect 50612 32572 50613 32612
rect 50571 32563 50613 32572
rect 48939 32528 48981 32537
rect 48939 32488 48940 32528
rect 48980 32488 48981 32528
rect 48939 32479 48981 32488
rect 48651 31100 48693 31109
rect 48651 31060 48652 31100
rect 48692 31060 48693 31100
rect 48651 31051 48693 31060
rect 48940 30344 48980 32479
rect 49324 30344 49364 32563
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 51532 32285 51572 34327
rect 51916 34292 51956 34301
rect 51916 34208 51956 34252
rect 51628 34168 51956 34208
rect 51628 32453 51668 34168
rect 51819 33704 51861 33713
rect 51819 33664 51820 33704
rect 51860 33664 51861 33704
rect 51819 33655 51861 33664
rect 51820 33140 51860 33655
rect 52204 33140 52244 34504
rect 81196 34376 81236 34915
rect 52491 34292 52533 34301
rect 52491 34252 52492 34292
rect 52532 34252 52533 34292
rect 52491 34243 52533 34252
rect 80812 34292 80852 34301
rect 52492 33872 52532 34243
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 52492 33823 52532 33832
rect 52683 33704 52725 33713
rect 52683 33664 52684 33704
rect 52724 33664 52725 33704
rect 52683 33655 52725 33664
rect 71979 33704 72021 33713
rect 71979 33664 71980 33704
rect 72020 33664 72021 33704
rect 71979 33655 72021 33664
rect 52684 33570 52724 33655
rect 53163 33620 53205 33629
rect 53163 33580 53164 33620
rect 53204 33580 53205 33620
rect 53163 33571 53205 33580
rect 52491 33452 52533 33461
rect 52491 33412 52492 33452
rect 52532 33412 52533 33452
rect 52491 33403 52533 33412
rect 52971 33452 53013 33461
rect 52971 33412 52972 33452
rect 53012 33412 53013 33452
rect 52971 33403 53013 33412
rect 52492 33318 52532 33403
rect 51724 33100 51860 33140
rect 51916 33100 52244 33140
rect 51724 32864 51764 33100
rect 51724 32815 51764 32824
rect 51916 32864 51956 33100
rect 51916 32815 51956 32824
rect 52300 32864 52340 32873
rect 52300 32621 52340 32824
rect 52299 32612 52341 32621
rect 52299 32572 52300 32612
rect 52340 32572 52341 32612
rect 52299 32563 52341 32572
rect 51627 32444 51669 32453
rect 51627 32404 51628 32444
rect 51668 32404 51669 32444
rect 51627 32395 51669 32404
rect 51531 32276 51573 32285
rect 51531 32236 51532 32276
rect 51572 32236 51573 32276
rect 51531 32227 51573 32236
rect 31756 30304 32097 30344
rect 32812 30304 32865 30344
rect 33004 30304 33057 30344
rect 47980 30304 48033 30344
rect 48940 30304 48993 30344
rect 30172 29979 30212 30304
rect 31516 29979 31556 30304
rect 32057 29960 32097 30304
rect 32825 29960 32865 30304
rect 33017 29960 33057 30304
rect 47993 29960 48033 30304
rect 48953 29960 48993 30304
rect 49180 30304 49364 30344
rect 52972 30344 53012 33403
rect 53164 32864 53204 33571
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 65931 33200 65973 33209
rect 65931 33160 65932 33200
rect 65972 33160 65973 33200
rect 65931 33151 65973 33160
rect 65547 33032 65589 33041
rect 65547 32992 65548 33032
rect 65588 32992 65589 33032
rect 65547 32983 65589 32992
rect 53164 32815 53204 32824
rect 64972 32864 65012 32873
rect 65260 32864 65300 32873
rect 65012 32824 65260 32864
rect 64972 32815 65012 32824
rect 65260 32815 65300 32824
rect 54316 32696 54356 32705
rect 54316 32453 54356 32656
rect 65548 32537 65588 32983
rect 65932 32873 65972 33151
rect 69772 33032 69812 33041
rect 65931 32864 65973 32873
rect 65931 32824 65932 32864
rect 65972 32824 65973 32864
rect 65931 32815 65973 32824
rect 66123 32864 66165 32873
rect 66123 32824 66124 32864
rect 66164 32824 66165 32864
rect 66123 32815 66165 32824
rect 65740 32696 65780 32705
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 65547 32528 65589 32537
rect 65547 32488 65548 32528
rect 65588 32488 65589 32528
rect 65547 32479 65589 32488
rect 53739 32444 53781 32453
rect 53739 32404 53740 32444
rect 53780 32404 53781 32444
rect 53739 32395 53781 32404
rect 54315 32444 54357 32453
rect 54315 32404 54316 32444
rect 54356 32404 54357 32444
rect 54315 32395 54357 32404
rect 53740 30344 53780 32395
rect 65740 31697 65780 32656
rect 66124 32537 66164 32815
rect 69772 32789 69812 32992
rect 70060 32957 70100 32988
rect 70059 32948 70101 32957
rect 70059 32908 70060 32948
rect 70100 32908 70101 32948
rect 70059 32899 70101 32908
rect 70060 32864 70100 32899
rect 69771 32780 69813 32789
rect 69771 32740 69772 32780
rect 69812 32740 69813 32780
rect 69771 32731 69813 32740
rect 70060 32621 70100 32824
rect 70059 32612 70101 32621
rect 70059 32572 70060 32612
rect 70100 32572 70101 32612
rect 70059 32563 70101 32572
rect 66123 32528 66165 32537
rect 66123 32488 66124 32528
rect 66164 32488 66165 32528
rect 66123 32479 66165 32488
rect 65739 31688 65781 31697
rect 65739 31648 65740 31688
rect 65780 31648 65781 31688
rect 65739 31639 65781 31648
rect 52972 30304 53025 30344
rect 53740 30304 53793 30344
rect 49180 29979 49220 30304
rect 52985 29960 53025 30304
rect 53753 29960 53793 30304
rect 18652 5648 18692 6021
rect 20537 5732 20577 6040
rect 22841 5732 22881 6040
rect 23225 5732 23265 6040
rect 23417 5732 23457 6040
rect 23609 5732 23649 6040
rect 23801 5732 23841 6040
rect 23993 5732 24033 6040
rect 25721 5732 25761 6040
rect 20428 5692 20577 5732
rect 22828 5692 22881 5732
rect 23212 5692 23265 5732
rect 23308 5692 23457 5732
rect 23500 5692 23649 5732
rect 23788 5692 23841 5732
rect 23980 5692 24033 5732
rect 25708 5692 25761 5732
rect 18652 5608 18740 5648
rect 14187 4220 14229 4229
rect 14187 4180 14188 4220
rect 14228 4180 14229 4220
rect 14187 4171 14229 4180
rect 13323 4136 13365 4145
rect 13323 4096 13324 4136
rect 13364 4096 13365 4136
rect 13323 4087 13365 4096
rect 12939 4052 12981 4061
rect 12939 4012 12940 4052
rect 12980 4012 12981 4052
rect 12939 4003 12981 4012
rect 8235 3968 8277 3977
rect 8235 3928 8236 3968
rect 8276 3928 8277 3968
rect 8235 3919 8277 3928
rect 7083 3464 7125 3473
rect 7083 3424 7084 3464
rect 7124 3424 7125 3464
rect 7083 3415 7125 3424
rect 12940 3464 12980 4003
rect 13324 3548 13364 4087
rect 14188 3809 14228 4171
rect 16203 4136 16245 4145
rect 16203 4096 16204 4136
rect 16244 4096 16245 4136
rect 16203 4087 16245 4096
rect 14187 3800 14229 3809
rect 14187 3760 14188 3800
rect 14228 3760 14229 3800
rect 14187 3751 14229 3760
rect 13324 3499 13364 3508
rect 12940 3053 12980 3424
rect 13228 3464 13268 3473
rect 12939 3044 12981 3053
rect 12939 3004 12940 3044
rect 12980 3004 12981 3044
rect 12939 2995 12981 3004
rect 13228 2969 13268 3424
rect 13804 3464 13844 3473
rect 13612 3296 13652 3305
rect 13804 3296 13844 3424
rect 14188 3464 14228 3751
rect 16204 3632 16244 4087
rect 18700 3809 18740 5608
rect 17259 3800 17301 3809
rect 17259 3760 17260 3800
rect 17300 3760 17301 3800
rect 17259 3751 17301 3760
rect 17451 3800 17493 3809
rect 17451 3760 17452 3800
rect 17492 3760 17493 3800
rect 17451 3751 17493 3760
rect 18699 3800 18741 3809
rect 18699 3760 18700 3800
rect 18740 3760 18741 3800
rect 18699 3751 18741 3760
rect 19275 3800 19317 3809
rect 19275 3760 19276 3800
rect 19316 3760 19317 3800
rect 19275 3751 19317 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 20331 3800 20373 3809
rect 20331 3760 20332 3800
rect 20372 3760 20373 3800
rect 20331 3751 20373 3760
rect 16204 3583 16244 3592
rect 17260 3477 17300 3751
rect 14188 3415 14228 3424
rect 15052 3464 15092 3473
rect 13652 3256 13844 3296
rect 13612 3247 13652 3256
rect 13227 2960 13269 2969
rect 13227 2920 13228 2960
rect 13268 2920 13269 2960
rect 13227 2911 13269 2920
rect 15052 2885 15092 3424
rect 16876 3464 16916 3473
rect 15051 2876 15093 2885
rect 15051 2836 15052 2876
rect 15092 2836 15093 2876
rect 15051 2827 15093 2836
rect 16876 2876 16916 3424
rect 17260 3137 17300 3437
rect 17259 3128 17301 3137
rect 17259 3088 17260 3128
rect 17300 3088 17301 3128
rect 17259 3079 17301 3088
rect 17355 2960 17397 2969
rect 17452 2960 17492 3751
rect 19276 3632 19316 3751
rect 19276 3583 19316 3592
rect 20332 3548 20372 3751
rect 20332 3499 20372 3508
rect 18124 3464 18164 3473
rect 17355 2920 17356 2960
rect 17396 2920 17492 2960
rect 17547 2960 17589 2969
rect 17547 2920 17548 2960
rect 17588 2920 17589 2960
rect 17355 2911 17397 2920
rect 17547 2911 17589 2920
rect 16876 2827 16916 2836
rect 17356 2792 17396 2911
rect 17164 2752 17396 2792
rect 6891 2708 6933 2717
rect 6891 2668 6892 2708
rect 6932 2668 6933 2708
rect 6891 2659 6933 2668
rect 17164 2624 17204 2752
rect 17164 2575 17204 2584
rect 17259 2624 17301 2633
rect 17259 2584 17260 2624
rect 17300 2584 17301 2624
rect 17259 2575 17301 2584
rect 17548 2624 17588 2911
rect 18124 2885 18164 3424
rect 20428 3464 20468 5692
rect 21291 3968 21333 3977
rect 21291 3928 21292 3968
rect 21332 3928 21333 3968
rect 21291 3919 21333 3928
rect 22155 3968 22197 3977
rect 22155 3928 22156 3968
rect 22196 3928 22197 3968
rect 22155 3919 22197 3928
rect 20044 3212 20084 3221
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 19947 2960 19989 2969
rect 19947 2920 19948 2960
rect 19988 2920 19989 2960
rect 19947 2911 19989 2920
rect 18123 2876 18165 2885
rect 18123 2836 18124 2876
rect 18164 2836 18165 2876
rect 18123 2827 18165 2836
rect 17548 2575 17588 2584
rect 17260 2490 17300 2575
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 18124 1961 18164 2827
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 19948 2120 19988 2911
rect 20044 2624 20084 3172
rect 20140 2624 20180 2633
rect 20044 2584 20140 2624
rect 20140 2575 20180 2584
rect 19660 2080 19988 2120
rect 18123 1952 18165 1961
rect 18123 1912 18124 1952
rect 18164 1912 18165 1952
rect 18123 1903 18165 1912
rect 18604 1700 18644 1709
rect 18644 1660 18740 1700
rect 18604 1651 18644 1660
rect 18700 1541 18740 1660
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 18699 1532 18741 1541
rect 18699 1492 18700 1532
rect 18740 1492 18741 1532
rect 18699 1483 18741 1492
rect 19660 1112 19700 2080
rect 19755 1952 19797 1961
rect 19755 1912 19756 1952
rect 19796 1912 19797 1952
rect 19755 1903 19797 1912
rect 19756 1818 19796 1903
rect 19947 1868 19989 1877
rect 19947 1828 19948 1868
rect 19988 1828 19989 1868
rect 19947 1819 19989 1828
rect 19660 1063 19700 1072
rect 19948 1112 19988 1819
rect 20428 1541 20468 3424
rect 20716 3464 20756 3473
rect 20523 3128 20565 3137
rect 20523 3088 20524 3128
rect 20564 3088 20565 3128
rect 20523 3079 20565 3088
rect 20524 2624 20564 3079
rect 20716 2969 20756 3424
rect 21292 3380 21332 3919
rect 22059 3800 22101 3809
rect 22059 3760 22060 3800
rect 22100 3760 22101 3800
rect 22059 3751 22101 3760
rect 21292 3053 21332 3340
rect 21772 3464 21812 3473
rect 21484 3212 21524 3221
rect 21772 3212 21812 3424
rect 21524 3172 21812 3212
rect 21484 3163 21524 3172
rect 21291 3044 21333 3053
rect 21291 3004 21292 3044
rect 21332 3004 21333 3044
rect 21291 2995 21333 3004
rect 20715 2960 20757 2969
rect 20715 2920 20716 2960
rect 20756 2920 20757 2960
rect 20715 2911 20757 2920
rect 21388 2624 21428 2633
rect 20564 2584 20660 2624
rect 20524 2575 20564 2584
rect 20620 1952 20660 2584
rect 21388 1961 21428 2584
rect 21772 1961 21812 3172
rect 22060 3464 22100 3751
rect 22156 3548 22196 3919
rect 22828 3809 22868 5692
rect 23212 3977 23252 5692
rect 23211 3968 23253 3977
rect 23211 3928 23212 3968
rect 23252 3928 23253 3968
rect 23211 3919 23253 3928
rect 22827 3800 22869 3809
rect 22827 3760 22828 3800
rect 22868 3760 22869 3800
rect 22827 3751 22869 3760
rect 22196 3508 22388 3548
rect 22156 3499 22196 3508
rect 22060 2969 22100 3424
rect 22059 2960 22101 2969
rect 22059 2920 22060 2960
rect 22100 2920 22101 2960
rect 22059 2911 22101 2920
rect 20620 1903 20660 1912
rect 21004 1952 21044 1961
rect 20043 1532 20085 1541
rect 20043 1492 20044 1532
rect 20084 1492 20085 1532
rect 20043 1483 20085 1492
rect 20427 1532 20469 1541
rect 20427 1492 20428 1532
rect 20468 1492 20469 1532
rect 20427 1483 20469 1492
rect 19948 1063 19988 1072
rect 20044 1112 20084 1483
rect 20332 1364 20372 1373
rect 21004 1364 21044 1912
rect 21387 1952 21429 1961
rect 21387 1912 21388 1952
rect 21428 1912 21429 1952
rect 21387 1903 21429 1912
rect 21771 1952 21813 1961
rect 21771 1912 21772 1952
rect 21812 1912 21813 1952
rect 21771 1903 21813 1912
rect 22155 1952 22197 1961
rect 22155 1912 22156 1952
rect 22196 1912 22197 1952
rect 22348 1952 22388 3508
rect 22636 3464 22676 3473
rect 22444 3296 22484 3305
rect 22636 3296 22676 3424
rect 22484 3256 22676 3296
rect 23020 3464 23060 3473
rect 22444 3247 22484 3256
rect 22539 2960 22581 2969
rect 22539 2920 22540 2960
rect 22580 2920 22581 2960
rect 22539 2911 22581 2920
rect 22540 2876 22580 2911
rect 22540 2825 22580 2836
rect 23020 2876 23060 3424
rect 23212 2876 23252 2885
rect 23020 2836 23212 2876
rect 22539 2036 22581 2045
rect 22539 1996 22540 2036
rect 22580 1996 22581 2036
rect 22539 1987 22581 1996
rect 22444 1952 22484 1961
rect 22348 1912 22444 1952
rect 22155 1903 22197 1912
rect 22444 1903 22484 1912
rect 22156 1818 22196 1903
rect 22540 1902 22580 1987
rect 22828 1700 22868 1709
rect 20372 1324 21044 1364
rect 22636 1660 22828 1700
rect 20332 1315 20372 1324
rect 20044 1063 20084 1072
rect 22636 1112 22676 1660
rect 22828 1651 22868 1660
rect 22636 1063 22676 1072
rect 23020 1112 23060 2836
rect 23212 2827 23252 2836
rect 23115 2624 23157 2633
rect 23115 2584 23116 2624
rect 23156 2584 23157 2624
rect 23115 2575 23157 2584
rect 23116 1961 23156 2575
rect 23212 2456 23252 2467
rect 23308 2456 23348 5692
rect 23403 3128 23445 3137
rect 23403 3088 23404 3128
rect 23444 3088 23445 3128
rect 23403 3079 23445 3088
rect 23404 2717 23444 3079
rect 23403 2708 23445 2717
rect 23403 2668 23404 2708
rect 23444 2668 23445 2708
rect 23403 2659 23445 2668
rect 23404 2574 23444 2659
rect 23500 2465 23540 5692
rect 23788 5405 23828 5692
rect 23787 5396 23829 5405
rect 23787 5356 23788 5396
rect 23828 5356 23829 5396
rect 23787 5347 23829 5356
rect 23980 4061 24020 5692
rect 25708 5573 25748 5692
rect 25948 5648 25988 6021
rect 26332 5909 26372 6021
rect 26331 5900 26373 5909
rect 26331 5860 26332 5900
rect 26372 5860 26373 5900
rect 26331 5851 26373 5860
rect 31708 5741 31748 6021
rect 31083 5732 31125 5741
rect 31083 5692 31084 5732
rect 31124 5692 31125 5732
rect 31083 5683 31125 5692
rect 31707 5732 31749 5741
rect 33785 5732 33825 6040
rect 33977 5732 34017 6040
rect 31707 5692 31708 5732
rect 31748 5692 31749 5732
rect 31707 5683 31749 5692
rect 33772 5692 33825 5732
rect 33868 5692 34017 5732
rect 25948 5608 26420 5648
rect 25707 5564 25749 5573
rect 25707 5524 25708 5564
rect 25748 5524 25749 5564
rect 25707 5515 25749 5524
rect 23979 4052 24021 4061
rect 23979 4012 23980 4052
rect 24020 4012 24021 4052
rect 23979 4003 24021 4012
rect 25035 3968 25077 3977
rect 25035 3928 25036 3968
rect 25076 3928 25077 3968
rect 25035 3919 25077 3928
rect 25036 3632 25076 3919
rect 25036 3583 25076 3592
rect 23884 3464 23924 3473
rect 23884 2633 23924 3424
rect 25804 2792 25844 2801
rect 25844 2752 26036 2792
rect 25804 2743 25844 2752
rect 25131 2708 25173 2717
rect 25131 2668 25132 2708
rect 25172 2668 25173 2708
rect 25131 2659 25173 2668
rect 23883 2624 23925 2633
rect 23883 2584 23884 2624
rect 23924 2584 23925 2624
rect 23883 2575 23925 2584
rect 25132 2624 25172 2659
rect 25132 2573 25172 2584
rect 25420 2624 25460 2633
rect 25420 2465 25460 2584
rect 25996 2624 26036 2752
rect 25996 2575 26036 2584
rect 26380 2624 26420 5608
rect 28395 3968 28437 3977
rect 28395 3928 28396 3968
rect 28436 3928 28437 3968
rect 28395 3919 28437 3928
rect 29451 3968 29493 3977
rect 29451 3928 29452 3968
rect 29492 3928 29493 3968
rect 29451 3919 29493 3928
rect 28396 3464 28436 3919
rect 27147 2876 27189 2885
rect 27147 2836 27148 2876
rect 27188 2836 27189 2876
rect 27147 2827 27189 2836
rect 26859 2708 26901 2717
rect 26859 2668 26860 2708
rect 26900 2668 26901 2708
rect 26859 2659 26901 2668
rect 25515 2540 25557 2549
rect 25515 2500 25516 2540
rect 25556 2500 25557 2540
rect 25515 2491 25557 2500
rect 23499 2456 23541 2465
rect 23308 2416 23444 2456
rect 23212 2381 23252 2416
rect 23211 2372 23253 2381
rect 23211 2332 23212 2372
rect 23252 2332 23253 2372
rect 23211 2323 23253 2332
rect 23404 2045 23444 2416
rect 23499 2416 23500 2456
rect 23540 2416 23541 2456
rect 23499 2407 23541 2416
rect 25419 2456 25461 2465
rect 25419 2416 25420 2456
rect 25460 2416 25461 2456
rect 25419 2407 25461 2416
rect 23403 2036 23445 2045
rect 23403 1996 23404 2036
rect 23444 1996 23445 2036
rect 23403 1987 23445 1996
rect 23500 2036 23540 2407
rect 25516 2406 25556 2491
rect 26380 2381 26420 2584
rect 26475 2456 26517 2465
rect 26475 2416 26476 2456
rect 26516 2416 26517 2456
rect 26475 2407 26517 2416
rect 24459 2372 24501 2381
rect 24459 2332 24460 2372
rect 24500 2332 24501 2372
rect 24459 2323 24501 2332
rect 26379 2372 26421 2381
rect 26379 2332 26380 2372
rect 26420 2332 26421 2372
rect 26379 2323 26421 2332
rect 23500 1987 23540 1996
rect 23115 1952 23157 1961
rect 23115 1912 23116 1952
rect 23156 1912 23157 1952
rect 23115 1903 23157 1912
rect 23404 1952 23444 1987
rect 23404 1903 23444 1912
rect 24076 1952 24116 1961
rect 23116 1818 23156 1903
rect 23788 1784 23828 1793
rect 24076 1784 24116 1912
rect 24460 1952 24500 2323
rect 26476 2120 26516 2407
rect 26476 2071 26516 2080
rect 25035 2036 25077 2045
rect 25035 1996 25036 2036
rect 25076 1996 25077 2036
rect 25035 1987 25077 1996
rect 24460 1903 24500 1912
rect 23828 1744 24116 1784
rect 23788 1735 23828 1744
rect 25036 1364 25076 1987
rect 25323 1952 25365 1961
rect 25323 1912 25324 1952
rect 25364 1912 25365 1952
rect 25323 1903 25365 1912
rect 26860 1952 26900 2659
rect 26860 1903 26900 1912
rect 27148 1952 27188 2827
rect 28396 2717 28436 3424
rect 28588 3592 28820 3632
rect 28588 2801 28628 3592
rect 28780 3548 28820 3592
rect 28780 3499 28820 3508
rect 28684 3464 28724 3473
rect 28587 2792 28629 2801
rect 28587 2752 28588 2792
rect 28628 2752 28629 2792
rect 28587 2743 28629 2752
rect 28395 2708 28437 2717
rect 28395 2668 28396 2708
rect 28436 2668 28437 2708
rect 28395 2659 28437 2668
rect 27243 2624 27285 2633
rect 27243 2584 27244 2624
rect 27284 2584 27285 2624
rect 27243 2575 27285 2584
rect 27244 2490 27284 2575
rect 28396 2549 28436 2580
rect 28395 2540 28437 2549
rect 28395 2500 28396 2540
rect 28436 2500 28437 2540
rect 28395 2491 28437 2500
rect 28107 2456 28149 2465
rect 28107 2416 28108 2456
rect 28148 2416 28149 2456
rect 28107 2407 28149 2416
rect 28396 2456 28436 2491
rect 27148 1903 27188 1912
rect 27244 1952 27284 1963
rect 25036 1315 25076 1324
rect 25324 1121 25364 1903
rect 27244 1877 27284 1912
rect 27724 1952 27764 1961
rect 27243 1868 27285 1877
rect 27243 1828 27244 1868
rect 27284 1828 27285 1868
rect 27243 1819 27285 1828
rect 27532 1784 27572 1793
rect 27724 1784 27764 1912
rect 28108 1952 28148 2407
rect 28396 2213 28436 2416
rect 28395 2204 28437 2213
rect 28395 2164 28396 2204
rect 28436 2164 28437 2204
rect 28395 2155 28437 2164
rect 28108 1903 28148 1912
rect 27572 1744 27764 1784
rect 27532 1735 27572 1744
rect 28684 1373 28724 3424
rect 29068 3212 29108 3221
rect 28780 3172 29068 3212
rect 28780 2624 28820 3172
rect 29068 3163 29108 3172
rect 28780 2575 28820 2584
rect 28971 2624 29013 2633
rect 28971 2584 28972 2624
rect 29012 2584 29013 2624
rect 28971 2575 29013 2584
rect 29164 2624 29204 2633
rect 28972 1961 29012 2575
rect 29164 2465 29204 2584
rect 29163 2456 29205 2465
rect 29163 2416 29164 2456
rect 29204 2416 29205 2456
rect 29163 2407 29205 2416
rect 28971 1952 29013 1961
rect 28971 1912 28972 1952
rect 29012 1912 29013 1952
rect 28971 1903 29013 1912
rect 28972 1818 29012 1903
rect 28683 1364 28725 1373
rect 28683 1324 28684 1364
rect 28724 1324 28725 1364
rect 28683 1315 28725 1324
rect 23020 1063 23060 1072
rect 23883 1112 23925 1121
rect 23883 1072 23884 1112
rect 23924 1072 23925 1112
rect 23883 1063 23925 1072
rect 25323 1112 25365 1121
rect 25323 1072 25324 1112
rect 25364 1072 25365 1112
rect 25323 1063 25365 1072
rect 29452 1112 29492 3919
rect 30891 3884 30933 3893
rect 30891 3844 30892 3884
rect 30932 3844 30933 3884
rect 30891 3835 30933 3844
rect 30796 3464 30836 3473
rect 30027 2624 30069 2633
rect 30027 2584 30028 2624
rect 30068 2584 30069 2624
rect 30027 2575 30069 2584
rect 30028 2490 30068 2575
rect 30699 2456 30741 2465
rect 30699 2416 30700 2456
rect 30740 2416 30741 2456
rect 30699 2407 30741 2416
rect 30123 2372 30165 2381
rect 30123 2332 30124 2372
rect 30164 2332 30165 2372
rect 30123 2323 30165 2332
rect 29739 2120 29781 2129
rect 29739 2080 29740 2120
rect 29780 2080 29781 2120
rect 29739 2071 29781 2080
rect 30124 2120 30164 2323
rect 29452 1063 29492 1072
rect 29740 1112 29780 2071
rect 30124 1877 30164 2080
rect 30123 1868 30165 1877
rect 30123 1828 30124 1868
rect 30164 1828 30165 1868
rect 30123 1819 30165 1828
rect 29835 1364 29877 1373
rect 29835 1324 29836 1364
rect 29876 1324 29877 1364
rect 29835 1315 29877 1324
rect 29740 1063 29780 1072
rect 29836 1112 29876 1315
rect 30124 1280 30164 1289
rect 30164 1240 30356 1280
rect 30124 1231 30164 1240
rect 29836 1063 29876 1072
rect 30316 1112 30356 1240
rect 30316 1063 30356 1072
rect 30700 1112 30740 2407
rect 30700 1063 30740 1072
rect 23884 978 23924 1063
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 30796 701 30836 3424
rect 30892 3380 30932 3835
rect 30987 3716 31029 3725
rect 30987 3676 30988 3716
rect 31028 3676 31029 3716
rect 30987 3667 31029 3676
rect 30892 3221 30932 3340
rect 30988 3296 31028 3667
rect 31084 3380 31124 5683
rect 33772 5489 33812 5692
rect 33387 5480 33429 5489
rect 33387 5440 33388 5480
rect 33428 5440 33429 5480
rect 33387 5431 33429 5440
rect 33771 5480 33813 5489
rect 33771 5440 33772 5480
rect 33812 5440 33813 5480
rect 33771 5431 33813 5440
rect 31179 5060 31221 5069
rect 31179 5020 31180 5060
rect 31220 5020 31221 5060
rect 31179 5011 31221 5020
rect 31180 3893 31220 5011
rect 33291 4136 33333 4145
rect 33291 4096 33292 4136
rect 33332 4096 33333 4136
rect 33291 4087 33333 4096
rect 31179 3884 31221 3893
rect 31179 3844 31180 3884
rect 31220 3844 31221 3884
rect 31179 3835 31221 3844
rect 31180 3464 31220 3835
rect 33292 3548 33332 4087
rect 33292 3499 33332 3508
rect 31180 3415 31220 3424
rect 33388 3464 33428 5431
rect 33675 3968 33717 3977
rect 33675 3928 33676 3968
rect 33716 3928 33717 3968
rect 33675 3919 33717 3928
rect 33388 3415 33428 3424
rect 33676 3464 33716 3919
rect 33676 3415 33716 3424
rect 32812 3380 32852 3389
rect 31084 3331 31124 3340
rect 32716 3340 32812 3380
rect 30988 3247 31028 3256
rect 30891 3212 30933 3221
rect 30891 3172 30892 3212
rect 30932 3172 30933 3212
rect 30891 3163 30933 3172
rect 32620 3212 32660 3221
rect 32235 3044 32277 3053
rect 32235 3004 32236 3044
rect 32276 3004 32277 3044
rect 32235 2995 32277 3004
rect 32043 2960 32085 2969
rect 32043 2920 32044 2960
rect 32084 2920 32085 2960
rect 32043 2911 32085 2920
rect 31275 2876 31317 2885
rect 31275 2836 31276 2876
rect 31316 2836 31317 2876
rect 31275 2827 31317 2836
rect 32044 2876 32084 2911
rect 31179 2792 31221 2801
rect 31179 2752 31180 2792
rect 31220 2752 31221 2792
rect 31179 2743 31221 2752
rect 31180 2658 31220 2743
rect 31276 1952 31316 2827
rect 32044 2825 32084 2836
rect 32236 2708 32276 2995
rect 32620 2717 32660 3172
rect 32716 3137 32756 3340
rect 32812 3331 32852 3340
rect 33004 3212 33044 3221
rect 32812 3172 33004 3212
rect 32715 3128 32757 3137
rect 32715 3088 32716 3128
rect 32756 3088 32757 3128
rect 32715 3079 32757 3088
rect 32236 2659 32276 2668
rect 32619 2708 32661 2717
rect 32619 2668 32620 2708
rect 32660 2668 32661 2708
rect 32619 2659 32661 2668
rect 31467 2540 31509 2549
rect 31467 2500 31468 2540
rect 31508 2500 31509 2540
rect 31467 2491 31509 2500
rect 31468 1961 31508 2491
rect 31659 2120 31701 2129
rect 31659 2080 31660 2120
rect 31700 2080 31701 2120
rect 31659 2071 31701 2080
rect 31563 2036 31605 2045
rect 31563 1996 31564 2036
rect 31604 1996 31605 2036
rect 31563 1987 31605 1996
rect 31660 2036 31700 2071
rect 31276 1903 31316 1912
rect 31467 1952 31509 1961
rect 31467 1912 31468 1952
rect 31508 1912 31509 1952
rect 31467 1903 31509 1912
rect 31564 1952 31604 1987
rect 31660 1985 31700 1996
rect 31468 1112 31508 1903
rect 31564 1901 31604 1912
rect 32140 1952 32180 1961
rect 31948 1784 31988 1793
rect 32140 1784 32180 1912
rect 32524 1952 32564 1961
rect 32620 1952 32660 2659
rect 32812 2624 32852 3172
rect 33004 3163 33044 3172
rect 33868 3053 33908 5692
rect 34396 5648 34436 6021
rect 34553 5732 34593 6040
rect 34745 5732 34785 6040
rect 34540 5692 34593 5732
rect 34732 5692 34785 5732
rect 34396 5608 34484 5648
rect 34251 4724 34293 4733
rect 34251 4684 34252 4724
rect 34292 4684 34293 4724
rect 34251 4675 34293 4684
rect 34155 3716 34197 3725
rect 34155 3676 34156 3716
rect 34196 3676 34197 3716
rect 34155 3667 34197 3676
rect 33963 3632 34005 3641
rect 33963 3592 33964 3632
rect 34004 3592 34005 3632
rect 33963 3583 34005 3592
rect 33964 3464 34004 3583
rect 33964 3415 34004 3424
rect 34060 3380 34100 3389
rect 34060 3221 34100 3340
rect 34156 3296 34196 3667
rect 34252 3380 34292 4675
rect 34444 4145 34484 5608
rect 34443 4136 34485 4145
rect 34443 4096 34444 4136
rect 34484 4096 34485 4136
rect 34443 4087 34485 4096
rect 34540 3968 34580 5692
rect 34732 4733 34772 5692
rect 34972 5648 35012 6021
rect 35164 5732 35204 6021
rect 35164 5692 35252 5732
rect 34972 5608 35156 5648
rect 34731 4724 34773 4733
rect 34731 4684 34732 4724
rect 34772 4684 34773 4724
rect 34731 4675 34773 4684
rect 35019 4136 35061 4145
rect 35019 4096 35020 4136
rect 35060 4096 35061 4136
rect 35019 4087 35061 4096
rect 34444 3928 34580 3968
rect 34347 3884 34389 3893
rect 34347 3844 34348 3884
rect 34388 3844 34389 3884
rect 34347 3835 34389 3844
rect 34348 3464 34388 3835
rect 34444 3632 34484 3928
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 34827 3632 34869 3641
rect 35020 3632 35060 4087
rect 34444 3592 34580 3632
rect 34348 3415 34388 3424
rect 34252 3331 34292 3340
rect 34156 3247 34196 3256
rect 34059 3212 34101 3221
rect 34059 3172 34060 3212
rect 34100 3172 34101 3212
rect 34059 3163 34101 3172
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 33867 3044 33909 3053
rect 33867 3004 33868 3044
rect 33908 3004 33909 3044
rect 33867 2995 33909 3004
rect 33195 2708 33237 2717
rect 33195 2668 33196 2708
rect 33236 2668 33237 2708
rect 33195 2659 33237 2668
rect 32812 2575 32852 2584
rect 33196 2624 33236 2659
rect 33196 2573 33236 2584
rect 34060 2624 34100 2633
rect 34060 1961 34100 2584
rect 34540 2456 34580 3592
rect 34827 3592 34828 3632
rect 34868 3592 34869 3632
rect 34827 3583 34869 3592
rect 34924 3592 35060 3632
rect 34636 3464 34676 3473
rect 34636 2969 34676 3424
rect 34635 2960 34677 2969
rect 34635 2920 34636 2960
rect 34676 2920 34677 2960
rect 34635 2911 34677 2920
rect 34828 2801 34868 3583
rect 34924 3464 34964 3592
rect 34924 3137 34964 3424
rect 35020 3464 35060 3473
rect 34923 3128 34965 3137
rect 34923 3088 34924 3128
rect 34964 3088 34965 3128
rect 34923 3079 34965 3088
rect 35020 3053 35060 3424
rect 35019 3044 35061 3053
rect 35019 3004 35020 3044
rect 35060 3004 35061 3044
rect 35019 2995 35061 3004
rect 34827 2792 34869 2801
rect 34827 2752 34828 2792
rect 34868 2752 34869 2792
rect 34827 2743 34869 2752
rect 34444 2416 34580 2456
rect 34444 2129 34484 2416
rect 35116 2381 35156 5608
rect 35212 3641 35252 5692
rect 35356 5648 35396 6021
rect 35513 5732 35553 6040
rect 36665 5732 36705 6040
rect 37433 5732 37473 6040
rect 35500 5692 35553 5732
rect 36556 5692 36705 5732
rect 37420 5692 37473 5732
rect 35356 5608 35444 5648
rect 35211 3632 35253 3641
rect 35211 3592 35212 3632
rect 35252 3592 35253 3632
rect 35211 3583 35253 3592
rect 35308 3212 35348 3221
rect 35211 3128 35253 3137
rect 35211 3088 35212 3128
rect 35252 3088 35253 3128
rect 35211 3079 35253 3088
rect 35212 2876 35252 3079
rect 35212 2827 35252 2836
rect 35308 2801 35348 3172
rect 35307 2792 35349 2801
rect 35307 2752 35308 2792
rect 35348 2752 35349 2792
rect 35307 2743 35349 2752
rect 35115 2372 35157 2381
rect 35115 2332 35116 2372
rect 35156 2332 35157 2372
rect 35115 2323 35157 2332
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 34443 2120 34485 2129
rect 34540 2120 34580 2129
rect 34443 2080 34444 2120
rect 34484 2080 34540 2120
rect 34443 2071 34485 2080
rect 34540 2071 34580 2080
rect 34828 2120 34868 2131
rect 34444 1986 34484 2071
rect 34828 2045 34868 2080
rect 34827 2036 34869 2045
rect 35404 2036 35444 5608
rect 35500 2045 35540 5692
rect 35979 2960 36021 2969
rect 35979 2920 35980 2960
rect 36020 2920 36116 2960
rect 35979 2911 36021 2920
rect 35787 2792 35829 2801
rect 35787 2752 35788 2792
rect 35828 2752 35829 2792
rect 35787 2743 35829 2752
rect 35788 2624 35828 2743
rect 35788 2575 35828 2584
rect 34827 1996 34828 2036
rect 34868 1996 34869 2036
rect 34827 1987 34869 1996
rect 35308 1996 35444 2036
rect 35499 2036 35541 2045
rect 35499 1996 35500 2036
rect 35540 1996 35541 2036
rect 32564 1912 32660 1952
rect 33387 1952 33429 1961
rect 33387 1912 33388 1952
rect 33428 1912 33429 1952
rect 32524 1903 32564 1912
rect 33387 1903 33429 1912
rect 34059 1952 34101 1961
rect 34059 1912 34060 1952
rect 34100 1912 34101 1952
rect 34059 1903 34101 1912
rect 33388 1818 33428 1903
rect 31988 1744 32180 1784
rect 31948 1735 31988 1744
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 35308 1373 35348 1996
rect 35499 1987 35541 1996
rect 35691 2036 35733 2045
rect 35691 1996 35692 2036
rect 35732 1996 35733 2036
rect 35691 1987 35733 1996
rect 35403 1868 35445 1877
rect 35403 1828 35404 1868
rect 35444 1828 35445 1868
rect 35403 1819 35445 1828
rect 32715 1364 32757 1373
rect 32715 1324 32716 1364
rect 32756 1324 32757 1364
rect 32715 1315 32757 1324
rect 35307 1364 35349 1373
rect 35307 1324 35308 1364
rect 35348 1324 35349 1364
rect 35307 1315 35349 1324
rect 35404 1364 35444 1819
rect 35404 1315 35444 1324
rect 32716 1230 32756 1315
rect 31564 1112 31604 1121
rect 31468 1072 31564 1112
rect 31564 1063 31604 1072
rect 35692 1112 35732 1987
rect 35979 1952 36021 1961
rect 35979 1912 35980 1952
rect 36020 1912 36021 1952
rect 35979 1903 36021 1912
rect 35980 1818 36020 1903
rect 36076 1205 36116 2920
rect 36171 2708 36213 2717
rect 36171 2668 36172 2708
rect 36212 2668 36213 2708
rect 36171 2659 36213 2668
rect 36172 2624 36212 2659
rect 36172 2573 36212 2584
rect 36556 1457 36596 5692
rect 36843 5228 36885 5237
rect 36843 5188 36844 5228
rect 36884 5188 36885 5228
rect 36843 5179 36885 5188
rect 36651 5060 36693 5069
rect 36651 5020 36652 5060
rect 36692 5020 36693 5060
rect 36651 5011 36693 5020
rect 36652 3464 36692 5011
rect 36652 3415 36692 3424
rect 36748 3380 36788 3389
rect 36748 3221 36788 3340
rect 36844 3296 36884 5179
rect 37323 5144 37365 5153
rect 37323 5104 37324 5144
rect 37364 5104 37365 5144
rect 37323 5095 37365 5104
rect 36939 4724 36981 4733
rect 36939 4684 36940 4724
rect 36980 4684 36981 4724
rect 36939 4675 36981 4684
rect 36940 3380 36980 4675
rect 37324 4556 37364 5095
rect 37420 4733 37460 5692
rect 37660 5648 37700 6021
rect 39545 5732 39585 6040
rect 39532 5692 39585 5732
rect 37660 5608 37940 5648
rect 37515 4976 37557 4985
rect 37515 4936 37516 4976
rect 37556 4936 37557 4976
rect 37515 4927 37557 4936
rect 37419 4724 37461 4733
rect 37419 4684 37420 4724
rect 37460 4684 37461 4724
rect 37419 4675 37461 4684
rect 37324 4516 37460 4556
rect 37035 3884 37077 3893
rect 37035 3844 37036 3884
rect 37076 3844 37077 3884
rect 37035 3835 37077 3844
rect 37036 3464 37076 3835
rect 37227 3632 37269 3641
rect 37227 3592 37228 3632
rect 37268 3592 37269 3632
rect 37227 3583 37269 3592
rect 37036 3415 37076 3424
rect 37228 3464 37268 3583
rect 37228 3415 37268 3424
rect 36940 3331 36980 3340
rect 37324 3380 37364 3389
rect 36844 3247 36884 3256
rect 37324 3221 37364 3340
rect 37420 3296 37460 4516
rect 37516 3380 37556 4927
rect 37611 3884 37653 3893
rect 37611 3844 37612 3884
rect 37652 3844 37653 3884
rect 37611 3835 37653 3844
rect 37612 3464 37652 3835
rect 37804 3464 37844 3473
rect 37652 3424 37804 3464
rect 37612 3415 37652 3424
rect 37804 3415 37844 3424
rect 37516 3331 37556 3340
rect 37900 3380 37940 5608
rect 39339 3632 39381 3641
rect 39339 3592 39340 3632
rect 39380 3592 39381 3632
rect 39339 3583 39381 3592
rect 38188 3464 38228 3473
rect 39244 3464 39284 3473
rect 38228 3424 38420 3464
rect 38188 3415 38228 3424
rect 37900 3331 37940 3340
rect 38092 3380 38132 3389
rect 37420 3247 37460 3256
rect 37995 3296 38037 3305
rect 37995 3256 37996 3296
rect 38036 3256 38037 3296
rect 37995 3247 38037 3256
rect 36747 3212 36789 3221
rect 36747 3172 36748 3212
rect 36788 3172 36789 3212
rect 36747 3163 36789 3172
rect 37323 3212 37365 3221
rect 37323 3172 37324 3212
rect 37364 3172 37365 3212
rect 37323 3163 37365 3172
rect 37996 3162 38036 3247
rect 38092 3221 38132 3340
rect 38091 3212 38133 3221
rect 38091 3172 38092 3212
rect 38132 3172 38133 3212
rect 38091 3163 38133 3172
rect 38187 3044 38229 3053
rect 38187 3004 38188 3044
rect 38228 3004 38229 3044
rect 38187 2995 38229 3004
rect 37995 2876 38037 2885
rect 37995 2836 37996 2876
rect 38036 2836 38037 2876
rect 37995 2827 38037 2836
rect 38188 2876 38228 2995
rect 38188 2827 38228 2836
rect 36843 2708 36885 2717
rect 36843 2668 36844 2708
rect 36884 2668 36885 2708
rect 36843 2659 36885 2668
rect 36844 2297 36884 2659
rect 37035 2624 37077 2633
rect 37035 2584 37036 2624
rect 37076 2584 37077 2624
rect 37035 2575 37077 2584
rect 37036 2490 37076 2575
rect 36843 2288 36885 2297
rect 36843 2248 36844 2288
rect 36884 2248 36885 2288
rect 36843 2239 36885 2248
rect 36844 1952 36884 2239
rect 36844 1903 36884 1912
rect 37228 1952 37268 1963
rect 37708 1952 37748 1961
rect 37228 1877 37268 1912
rect 37612 1912 37708 1952
rect 37227 1868 37269 1877
rect 37227 1828 37228 1868
rect 37268 1828 37269 1868
rect 37227 1819 37269 1828
rect 36555 1448 36597 1457
rect 36555 1408 36556 1448
rect 36596 1408 36597 1448
rect 36555 1399 36597 1408
rect 37612 1364 37652 1912
rect 37708 1903 37748 1912
rect 37612 1315 37652 1324
rect 37899 1280 37941 1289
rect 37899 1240 37900 1280
rect 37940 1240 37941 1280
rect 37899 1231 37941 1240
rect 36075 1196 36117 1205
rect 36075 1156 36076 1196
rect 36116 1156 36117 1196
rect 36075 1147 36117 1156
rect 35692 1063 35732 1072
rect 35787 1112 35829 1121
rect 35787 1072 35788 1112
rect 35828 1072 35829 1112
rect 35787 1063 35829 1072
rect 36076 1112 36116 1147
rect 37900 1121 37940 1231
rect 35788 978 35828 1063
rect 36076 1061 36116 1072
rect 37899 1112 37941 1121
rect 37899 1072 37900 1112
rect 37940 1072 37941 1112
rect 37899 1063 37941 1072
rect 37996 1112 38036 2827
rect 38091 2540 38133 2549
rect 38091 2500 38092 2540
rect 38132 2500 38133 2540
rect 38091 2491 38133 2500
rect 38092 2297 38132 2491
rect 38091 2288 38133 2297
rect 38091 2248 38092 2288
rect 38132 2248 38133 2288
rect 38091 2239 38133 2248
rect 38092 1952 38132 2239
rect 38092 1903 38132 1912
rect 38283 1196 38325 1205
rect 38283 1156 38284 1196
rect 38324 1156 38325 1196
rect 38283 1147 38325 1156
rect 37996 1063 38036 1072
rect 38284 1112 38324 1147
rect 37900 978 37940 1063
rect 38284 1061 38324 1072
rect 38380 869 38420 3424
rect 38956 3212 38996 3221
rect 38956 2624 38996 3172
rect 39244 2885 39284 3424
rect 39340 3464 39380 3583
rect 39340 3415 39380 3424
rect 39243 2876 39285 2885
rect 39243 2836 39244 2876
rect 39284 2836 39285 2876
rect 39243 2827 39285 2836
rect 38956 2575 38996 2584
rect 39340 2624 39380 2635
rect 39340 2549 39380 2584
rect 39339 2540 39381 2549
rect 39339 2500 39340 2540
rect 39380 2500 39381 2540
rect 39339 2491 39381 2500
rect 38955 2036 38997 2045
rect 38955 1996 38956 2036
rect 38996 1996 38997 2036
rect 38955 1987 38997 1996
rect 38956 1952 38996 1987
rect 38956 1901 38996 1912
rect 39532 1037 39572 5692
rect 39772 5648 39812 6021
rect 39929 5732 39969 6040
rect 39916 5692 39969 5732
rect 39772 5608 39860 5648
rect 39628 3464 39668 3473
rect 39628 2969 39668 3424
rect 39627 2960 39669 2969
rect 39627 2920 39628 2960
rect 39668 2920 39669 2960
rect 39627 2911 39669 2920
rect 39628 1205 39668 2911
rect 39820 2900 39860 5608
rect 39724 2885 39860 2900
rect 39723 2876 39860 2885
rect 39723 2836 39724 2876
rect 39764 2860 39860 2876
rect 39764 2836 39765 2860
rect 39723 2827 39765 2836
rect 39819 2204 39861 2213
rect 39819 2164 39820 2204
rect 39860 2164 39861 2204
rect 39819 2155 39861 2164
rect 39820 1541 39860 2155
rect 39916 2120 39956 5692
rect 40156 5648 40196 6021
rect 40313 5732 40353 6040
rect 40300 5692 40353 5732
rect 40156 5608 40244 5648
rect 40204 2792 40244 5608
rect 40300 3641 40340 5692
rect 40540 5648 40580 6021
rect 40697 5732 40737 6040
rect 40889 5909 40929 6040
rect 40888 5900 40930 5909
rect 40684 5692 40737 5732
rect 40876 5860 40889 5900
rect 40929 5860 40930 5900
rect 40876 5851 40930 5860
rect 40540 5608 40628 5648
rect 40299 3632 40341 3641
rect 40299 3592 40300 3632
rect 40340 3592 40341 3632
rect 40299 3583 40341 3592
rect 40204 2752 40340 2792
rect 40204 2624 40244 2633
rect 40108 2120 40148 2129
rect 39916 2080 40108 2120
rect 39819 1532 39861 1541
rect 39819 1492 39820 1532
rect 39860 1492 39861 1532
rect 39819 1483 39861 1492
rect 39627 1196 39669 1205
rect 39627 1156 39628 1196
rect 39668 1156 39669 1196
rect 39627 1147 39669 1156
rect 39628 1112 39668 1147
rect 39820 1112 39860 1483
rect 39916 1289 39956 2080
rect 40108 2071 40148 2080
rect 40204 2045 40244 2584
rect 40203 2036 40245 2045
rect 40203 1996 40204 2036
rect 40244 1996 40245 2036
rect 40203 1987 40245 1996
rect 40300 1868 40340 2752
rect 40588 2213 40628 5608
rect 40684 4985 40724 5692
rect 40683 4976 40725 4985
rect 40683 4936 40684 4976
rect 40724 4936 40725 4976
rect 40683 4927 40725 4936
rect 40876 2717 40916 5851
rect 43001 5732 43041 6040
rect 42988 5692 43041 5732
rect 42699 3464 42741 3473
rect 42699 3424 42700 3464
rect 42740 3424 42741 3464
rect 42699 3415 42741 3424
rect 42412 3380 42452 3389
rect 42220 3212 42260 3221
rect 41259 2960 41301 2969
rect 41259 2920 41260 2960
rect 41300 2920 41301 2960
rect 41259 2911 41301 2920
rect 40875 2708 40917 2717
rect 40875 2668 40876 2708
rect 40916 2668 40917 2708
rect 40875 2659 40917 2668
rect 40875 2540 40917 2549
rect 40875 2500 40876 2540
rect 40916 2500 40917 2540
rect 40875 2491 40917 2500
rect 40587 2204 40629 2213
rect 40587 2164 40588 2204
rect 40628 2164 40629 2204
rect 40587 2155 40629 2164
rect 40012 1828 40340 1868
rect 40012 1373 40052 1828
rect 40011 1364 40053 1373
rect 40011 1324 40012 1364
rect 40052 1324 40053 1364
rect 40011 1315 40053 1324
rect 39915 1280 39957 1289
rect 39915 1240 39916 1280
rect 39956 1240 39957 1280
rect 39915 1231 39957 1240
rect 39916 1112 39956 1121
rect 39820 1072 39916 1112
rect 39628 1061 39668 1072
rect 39916 1063 39956 1072
rect 40012 1112 40052 1315
rect 40300 1280 40340 1289
rect 40340 1240 40532 1280
rect 40300 1231 40340 1240
rect 40012 1063 40052 1072
rect 40492 1112 40532 1240
rect 40492 1063 40532 1072
rect 40876 1112 40916 2491
rect 41260 1952 41300 2911
rect 42220 2900 42260 3172
rect 42412 2969 42452 3340
rect 42700 3330 42740 3415
rect 42411 2960 42453 2969
rect 42411 2920 42412 2960
rect 42452 2920 42453 2960
rect 42411 2911 42453 2920
rect 41355 2876 41397 2885
rect 41355 2836 41356 2876
rect 41396 2836 41397 2876
rect 42220 2860 42356 2900
rect 41355 2827 41397 2836
rect 41356 2742 41396 2827
rect 42316 2624 42356 2860
rect 42795 2708 42837 2717
rect 42795 2668 42796 2708
rect 42836 2668 42837 2708
rect 42795 2659 42837 2668
rect 42412 2624 42452 2633
rect 42316 2584 42412 2624
rect 41643 2204 41685 2213
rect 41643 2164 41644 2204
rect 41684 2164 41685 2204
rect 41643 2155 41685 2164
rect 42123 2204 42165 2213
rect 42123 2164 42124 2204
rect 42164 2164 42165 2204
rect 42123 2155 42165 2164
rect 41644 2036 41684 2155
rect 42124 2120 42164 2155
rect 42124 2069 42164 2080
rect 41644 1987 41684 1996
rect 41739 2036 41781 2045
rect 41739 1996 41740 2036
rect 41780 1996 41781 2036
rect 41739 1987 41781 1996
rect 41260 1903 41300 1912
rect 41548 1952 41588 1961
rect 41548 1373 41588 1912
rect 41547 1364 41589 1373
rect 41547 1324 41548 1364
rect 41588 1324 41589 1364
rect 41547 1315 41589 1324
rect 40876 1063 40916 1072
rect 41740 1112 41780 1987
rect 41931 1784 41973 1793
rect 41931 1744 41932 1784
rect 41972 1744 41973 1784
rect 41931 1735 41973 1744
rect 41932 1650 41972 1735
rect 42412 1121 42452 2584
rect 42700 2624 42740 2633
rect 42700 2213 42740 2584
rect 42796 2624 42836 2659
rect 42796 2573 42836 2584
rect 42699 2204 42741 2213
rect 42699 2164 42700 2204
rect 42740 2164 42741 2204
rect 42699 2155 42741 2164
rect 42988 1541 43028 5692
rect 46876 5648 46916 6021
rect 47068 5648 47108 6021
rect 47260 5648 47300 6021
rect 47417 5732 47457 6040
rect 47609 5732 47649 6040
rect 47404 5692 47457 5732
rect 47596 5692 47649 5732
rect 46876 5608 46964 5648
rect 47068 5608 47156 5648
rect 47260 5608 47348 5648
rect 44907 3632 44949 3641
rect 44907 3592 44908 3632
rect 44948 3592 44949 3632
rect 44907 3583 44949 3592
rect 44523 3380 44565 3389
rect 44523 3340 44524 3380
rect 44564 3340 44565 3380
rect 44523 3331 44565 3340
rect 44524 3246 44564 3331
rect 43083 2792 43125 2801
rect 43083 2752 43084 2792
rect 43124 2752 43125 2792
rect 43083 2743 43125 2752
rect 43084 2658 43124 2743
rect 43275 2708 43317 2717
rect 43275 2668 43276 2708
rect 43316 2668 43317 2708
rect 43275 2659 43317 2668
rect 43276 2574 43316 2659
rect 44428 2624 44468 2633
rect 44139 2540 44181 2549
rect 44139 2500 44140 2540
rect 44180 2500 44181 2540
rect 44139 2491 44181 2500
rect 43275 2036 43317 2045
rect 43275 1996 43276 2036
rect 43316 1996 43317 2036
rect 43275 1987 43317 1996
rect 43276 1952 43316 1987
rect 43276 1901 43316 1912
rect 44140 1952 44180 2491
rect 44428 2045 44468 2584
rect 44908 2120 44948 3583
rect 46924 3557 46964 5608
rect 47116 3725 47156 5608
rect 47308 3809 47348 5608
rect 47307 3800 47349 3809
rect 47307 3760 47308 3800
rect 47348 3760 47349 3800
rect 47307 3751 47349 3760
rect 47115 3716 47157 3725
rect 47115 3676 47116 3716
rect 47156 3676 47157 3716
rect 47115 3667 47157 3676
rect 46443 3548 46485 3557
rect 46443 3508 46444 3548
rect 46484 3508 46485 3548
rect 46443 3499 46485 3508
rect 46923 3548 46965 3557
rect 46923 3508 46924 3548
rect 46964 3508 46965 3548
rect 46923 3499 46965 3508
rect 46060 3464 46100 3473
rect 45964 3424 46060 3464
rect 45196 3380 45236 3389
rect 45004 3212 45044 3221
rect 45004 2549 45044 3172
rect 45003 2540 45045 2549
rect 45003 2500 45004 2540
rect 45044 2500 45045 2540
rect 45003 2491 45045 2500
rect 45196 2129 45236 3340
rect 45675 2792 45717 2801
rect 45675 2752 45676 2792
rect 45716 2752 45717 2792
rect 45675 2743 45717 2752
rect 45292 2624 45332 2635
rect 45292 2549 45332 2584
rect 45676 2624 45716 2743
rect 45676 2575 45716 2584
rect 45291 2540 45333 2549
rect 45291 2500 45292 2540
rect 45332 2500 45333 2540
rect 45291 2491 45333 2500
rect 44908 2071 44948 2080
rect 45195 2120 45237 2129
rect 45195 2080 45196 2120
rect 45236 2080 45237 2120
rect 45195 2071 45237 2080
rect 44427 2036 44469 2045
rect 44427 1996 44428 2036
rect 44468 1996 44469 2036
rect 44427 1987 44469 1996
rect 44140 1903 44180 1912
rect 44524 1952 44564 1961
rect 44524 1793 44564 1912
rect 44523 1784 44565 1793
rect 44523 1744 44524 1784
rect 44564 1744 44565 1784
rect 44523 1735 44565 1744
rect 44908 1700 44948 1709
rect 42987 1532 43029 1541
rect 42987 1492 42988 1532
rect 43028 1492 43029 1532
rect 42987 1483 43029 1492
rect 42891 1364 42933 1373
rect 42891 1324 42892 1364
rect 42932 1324 42933 1364
rect 42891 1315 42933 1324
rect 42892 1230 42932 1315
rect 41740 1063 41780 1072
rect 42411 1112 42453 1121
rect 42411 1072 42412 1112
rect 42452 1072 42453 1112
rect 42411 1063 42453 1072
rect 44427 1112 44469 1121
rect 44427 1072 44428 1112
rect 44468 1072 44469 1112
rect 44427 1063 44469 1072
rect 44716 1112 44756 1123
rect 39531 1028 39573 1037
rect 39531 988 39532 1028
rect 39572 988 39573 1028
rect 39531 979 39573 988
rect 44428 978 44468 1063
rect 44716 1037 44756 1072
rect 44812 1112 44852 1121
rect 44908 1112 44948 1660
rect 45099 1364 45141 1373
rect 45099 1324 45100 1364
rect 45140 1324 45141 1364
rect 45099 1315 45141 1324
rect 45100 1230 45140 1315
rect 45964 1121 46004 3424
rect 46060 3415 46100 3424
rect 46348 3464 46388 3473
rect 46348 3053 46388 3424
rect 46444 3414 46484 3499
rect 46732 3212 46772 3221
rect 46347 3044 46389 3053
rect 46347 3004 46348 3044
rect 46388 3004 46389 3044
rect 46347 2995 46389 3004
rect 46059 2708 46101 2717
rect 46059 2668 46060 2708
rect 46100 2668 46101 2708
rect 46059 2659 46101 2668
rect 46060 1952 46100 2659
rect 46732 2624 46772 3172
rect 46732 2575 46772 2584
rect 47116 2624 47156 2635
rect 47116 2549 47156 2584
rect 46923 2540 46965 2549
rect 46923 2500 46924 2540
rect 46964 2500 46965 2540
rect 46923 2491 46965 2500
rect 47115 2540 47157 2549
rect 47115 2500 47116 2540
rect 47156 2500 47157 2540
rect 47115 2491 47157 2500
rect 46060 1903 46100 1912
rect 46924 1952 46964 2491
rect 46924 1903 46964 1912
rect 47308 1952 47348 1961
rect 47211 1448 47253 1457
rect 47211 1408 47212 1448
rect 47252 1408 47253 1448
rect 47211 1399 47253 1408
rect 44852 1072 44948 1112
rect 45963 1112 46005 1121
rect 45963 1072 45964 1112
rect 46004 1072 46005 1112
rect 44812 1063 44852 1072
rect 45963 1063 46005 1072
rect 46923 1112 46965 1121
rect 46923 1072 46924 1112
rect 46964 1072 46965 1112
rect 46923 1063 46965 1072
rect 47212 1112 47252 1399
rect 47308 1373 47348 1912
rect 47307 1364 47349 1373
rect 47307 1324 47308 1364
rect 47348 1324 47349 1364
rect 47307 1315 47349 1324
rect 47404 1205 47444 5692
rect 47596 3641 47636 5692
rect 48939 3968 48981 3977
rect 48939 3928 48940 3968
rect 48980 3928 48981 3968
rect 48939 3919 48981 3928
rect 48651 3716 48693 3725
rect 48651 3676 48652 3716
rect 48692 3676 48693 3716
rect 48940 3716 48980 3919
rect 52395 3884 52437 3893
rect 52395 3844 52396 3884
rect 52436 3844 52437 3884
rect 52395 3835 52437 3844
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 52299 3800 52341 3809
rect 52299 3760 52300 3800
rect 52340 3760 52341 3800
rect 52299 3751 52341 3760
rect 49611 3716 49653 3725
rect 48940 3676 49076 3716
rect 48651 3667 48693 3676
rect 47595 3632 47637 3641
rect 47595 3592 47596 3632
rect 47636 3592 47637 3632
rect 47595 3583 47637 3592
rect 48652 3464 48692 3667
rect 48747 3632 48789 3641
rect 48747 3592 48748 3632
rect 48788 3592 48980 3632
rect 48747 3583 48789 3592
rect 48652 3415 48692 3424
rect 48940 3464 48980 3592
rect 49036 3557 49076 3676
rect 49611 3676 49612 3716
rect 49652 3676 49653 3716
rect 49611 3667 49653 3676
rect 51819 3716 51861 3725
rect 51819 3676 51820 3716
rect 51860 3676 51861 3716
rect 51819 3667 51861 3676
rect 49035 3548 49077 3557
rect 49035 3508 49036 3548
rect 49076 3508 49077 3548
rect 49035 3499 49077 3508
rect 48940 3296 48980 3424
rect 49036 3414 49076 3499
rect 49612 3296 49652 3667
rect 51820 3464 51860 3667
rect 52203 3632 52245 3641
rect 52203 3592 52204 3632
rect 52244 3592 52245 3632
rect 52203 3583 52245 3592
rect 52107 3548 52149 3557
rect 52107 3508 52108 3548
rect 52148 3508 52149 3548
rect 52107 3499 52149 3508
rect 52204 3548 52244 3583
rect 51820 3415 51860 3424
rect 52108 3464 52148 3499
rect 52204 3497 52244 3508
rect 48940 3256 49172 3296
rect 49612 3256 49748 3296
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 49132 2876 49172 3256
rect 49324 3212 49364 3221
rect 49364 3172 49652 3212
rect 49324 3163 49364 3172
rect 49132 2827 49172 2836
rect 47979 2792 48021 2801
rect 47979 2752 47980 2792
rect 48020 2752 48021 2792
rect 47979 2743 48021 2752
rect 48651 2792 48693 2801
rect 48651 2752 48652 2792
rect 48692 2752 48693 2792
rect 48651 2743 48693 2752
rect 47980 2624 48020 2743
rect 47980 2575 48020 2584
rect 48652 1952 48692 2743
rect 49612 2624 49652 3172
rect 49612 2575 49652 2584
rect 49515 2540 49557 2549
rect 49515 2500 49516 2540
rect 49556 2500 49557 2540
rect 49515 2491 49557 2500
rect 48652 1903 48692 1912
rect 49516 1952 49556 2491
rect 49708 2456 49748 3256
rect 52012 2876 52052 2885
rect 52108 2876 52148 3424
rect 52300 2969 52340 3751
rect 52396 3557 52436 3835
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 54603 3716 54645 3725
rect 54603 3676 54604 3716
rect 54644 3676 54645 3716
rect 54603 3667 54645 3676
rect 57771 3716 57813 3725
rect 57771 3676 57772 3716
rect 57812 3676 57813 3716
rect 57771 3667 57813 3676
rect 52395 3548 52437 3557
rect 52395 3508 52396 3548
rect 52436 3508 52437 3548
rect 52395 3499 52437 3508
rect 52299 2960 52341 2969
rect 52299 2920 52300 2960
rect 52340 2920 52341 2960
rect 52299 2911 52341 2920
rect 52052 2836 52148 2876
rect 52012 2827 52052 2836
rect 50859 2792 50901 2801
rect 50859 2752 50860 2792
rect 50900 2752 50901 2792
rect 50859 2743 50901 2752
rect 51243 2792 51285 2801
rect 51243 2752 51244 2792
rect 51284 2752 51285 2792
rect 51243 2743 51285 2752
rect 49996 2624 50036 2635
rect 49996 2549 50036 2584
rect 50860 2624 50900 2743
rect 50860 2575 50900 2584
rect 49995 2540 50037 2549
rect 49995 2500 49996 2540
rect 50036 2500 50037 2540
rect 49995 2491 50037 2500
rect 49516 1903 49556 1912
rect 49612 2416 49748 2456
rect 47500 1700 47540 1709
rect 47403 1196 47445 1205
rect 47403 1156 47404 1196
rect 47444 1156 47445 1196
rect 47403 1147 47445 1156
rect 47212 1063 47252 1072
rect 44715 1028 44757 1037
rect 44715 988 44716 1028
rect 44756 988 44757 1028
rect 44715 979 44757 988
rect 46924 978 46964 1063
rect 47500 1037 47540 1660
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 47595 1364 47637 1373
rect 47595 1324 47596 1364
rect 47636 1324 47637 1364
rect 47595 1315 47637 1324
rect 47596 1230 47636 1315
rect 49612 1289 49652 2416
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 49900 1952 49940 1961
rect 49900 1373 49940 1912
rect 51244 1952 51284 2743
rect 52107 2540 52149 2549
rect 52107 2500 52108 2540
rect 52148 2500 52149 2540
rect 52107 2491 52149 2500
rect 51244 1903 51284 1912
rect 52108 1952 52148 2491
rect 52108 1903 52148 1912
rect 50283 1868 50325 1877
rect 50283 1828 50284 1868
rect 50324 1828 50325 1868
rect 50283 1819 50325 1828
rect 50092 1700 50132 1709
rect 49996 1660 50092 1700
rect 49996 1457 50036 1660
rect 50092 1651 50132 1660
rect 49995 1448 50037 1457
rect 49995 1408 49996 1448
rect 50036 1408 50037 1448
rect 49995 1399 50037 1408
rect 49899 1364 49941 1373
rect 49899 1324 49900 1364
rect 49940 1324 49941 1364
rect 49899 1315 49941 1324
rect 49611 1280 49653 1289
rect 49611 1240 49612 1280
rect 49652 1240 49653 1280
rect 49611 1231 49653 1240
rect 49612 1112 49652 1231
rect 49899 1196 49941 1205
rect 49899 1156 49900 1196
rect 49940 1156 49941 1196
rect 49899 1147 49941 1156
rect 49612 1063 49652 1072
rect 49900 1112 49940 1147
rect 49900 1061 49940 1072
rect 49996 1112 50036 1399
rect 50284 1364 50324 1819
rect 50284 1315 50324 1324
rect 49996 1063 50036 1072
rect 52108 1112 52148 1121
rect 52300 1112 52340 2911
rect 52148 1072 52340 1112
rect 52396 1112 52436 3499
rect 54604 3464 54644 3667
rect 54891 3632 54933 3641
rect 54891 3592 54892 3632
rect 54932 3592 54933 3632
rect 54891 3583 54933 3592
rect 55179 3632 55221 3641
rect 55179 3592 55180 3632
rect 55220 3592 55221 3632
rect 55179 3583 55221 3592
rect 54604 3415 54644 3424
rect 54892 3464 54932 3583
rect 54987 3548 55029 3557
rect 54987 3508 54988 3548
rect 55028 3508 55029 3548
rect 54987 3499 55029 3508
rect 54892 3415 54932 3424
rect 54988 3414 55028 3499
rect 52492 3212 52532 3221
rect 52532 3172 52820 3212
rect 52492 3163 52532 3172
rect 52780 2624 52820 3172
rect 55180 2876 55220 3583
rect 55180 2827 55220 2836
rect 55276 3212 55316 3221
rect 53835 2708 53877 2717
rect 53835 2668 53836 2708
rect 53876 2668 53877 2708
rect 53835 2659 53877 2668
rect 54027 2708 54069 2717
rect 54027 2668 54028 2708
rect 54068 2668 54093 2708
rect 54027 2659 54093 2668
rect 52780 2575 52820 2584
rect 53164 2624 53204 2635
rect 53164 2549 53204 2584
rect 53163 2540 53205 2549
rect 53163 2500 53164 2540
rect 53204 2500 53205 2540
rect 53163 2491 53205 2500
rect 52492 1952 52532 1963
rect 52492 1877 52532 1912
rect 53836 1952 53876 2659
rect 54053 2624 54093 2659
rect 55276 2624 55316 3172
rect 55755 2876 55797 2885
rect 55755 2836 55756 2876
rect 55796 2836 55797 2876
rect 55755 2827 55797 2836
rect 57772 2876 57812 3667
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 57772 2827 57812 2836
rect 55372 2624 55412 2633
rect 55276 2584 55372 2624
rect 54053 2575 54093 2584
rect 55372 2575 55412 2584
rect 55756 2624 55796 2827
rect 56619 2708 56661 2717
rect 56619 2668 56620 2708
rect 56660 2668 56661 2708
rect 56619 2659 56661 2668
rect 55756 2129 55796 2584
rect 56620 2624 56660 2659
rect 71980 2633 72020 33655
rect 80812 33545 80852 34252
rect 80811 33536 80853 33545
rect 80811 33496 80812 33536
rect 80852 33496 80853 33536
rect 80811 33487 80853 33496
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 80715 32780 80757 32789
rect 80715 32740 80716 32780
rect 80756 32740 80757 32780
rect 80715 32731 80757 32740
rect 78507 32612 78549 32621
rect 78507 32572 78508 32612
rect 78548 32572 78549 32612
rect 78507 32563 78549 32572
rect 74187 30932 74229 30941
rect 74187 30892 74188 30932
rect 74228 30892 74229 30932
rect 74187 30883 74229 30892
rect 74188 17072 74228 30883
rect 78508 30689 78548 32563
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 78316 30680 78356 30689
rect 78316 30437 78356 30640
rect 78507 30680 78549 30689
rect 78507 30640 78508 30680
rect 78548 30640 78549 30680
rect 78507 30631 78549 30640
rect 78699 30680 78741 30689
rect 78699 30640 78700 30680
rect 78740 30640 78741 30680
rect 78699 30631 78741 30640
rect 78700 30546 78740 30631
rect 78892 30437 78932 30522
rect 78315 30428 78357 30437
rect 78315 30388 78316 30428
rect 78356 30388 78357 30428
rect 78315 30379 78357 30388
rect 78891 30428 78933 30437
rect 78891 30388 78892 30428
rect 78932 30388 78933 30428
rect 78891 30379 78933 30388
rect 78316 27380 78356 30379
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 78028 27340 78356 27380
rect 80716 27380 80756 32731
rect 80811 32192 80853 32201
rect 80811 32152 80812 32192
rect 80852 32152 80853 32192
rect 80811 32143 80853 32152
rect 81196 32192 81236 34336
rect 82060 34376 82100 34385
rect 81867 33788 81909 33797
rect 81867 33748 81868 33788
rect 81908 33748 81909 33788
rect 81867 33739 81909 33748
rect 81868 33654 81908 33739
rect 81964 33704 82004 33713
rect 81579 33536 81621 33545
rect 81579 33496 81580 33536
rect 81620 33496 81621 33536
rect 81579 33487 81621 33496
rect 81580 33402 81620 33487
rect 80812 32058 80852 32143
rect 80907 31268 80949 31277
rect 80907 31228 80908 31268
rect 80948 31228 80949 31268
rect 80907 31219 80949 31228
rect 80811 27656 80853 27665
rect 80811 27616 80812 27656
rect 80852 27616 80853 27656
rect 80811 27607 80853 27616
rect 80812 27522 80852 27607
rect 80716 27340 80852 27380
rect 75627 23120 75669 23129
rect 75627 23080 75628 23120
rect 75668 23080 75669 23120
rect 75627 23071 75669 23080
rect 74188 17023 74228 17032
rect 75628 16988 75668 23071
rect 75628 13805 75668 16948
rect 77451 15560 77493 15569
rect 77451 15520 77452 15560
rect 77492 15520 77493 15560
rect 77451 15511 77493 15520
rect 76395 14720 76437 14729
rect 76395 14680 76396 14720
rect 76436 14680 76437 14720
rect 76395 14671 76437 14680
rect 76396 13964 76436 14671
rect 76396 13915 76436 13924
rect 74091 13796 74133 13805
rect 74091 13756 74092 13796
rect 74132 13756 74133 13796
rect 74091 13747 74133 13756
rect 75627 13796 75669 13805
rect 76204 13796 76244 13805
rect 75627 13756 75628 13796
rect 75668 13756 75669 13796
rect 75627 13747 75669 13756
rect 76012 13756 76204 13796
rect 73419 7916 73461 7925
rect 73419 7876 73420 7916
rect 73460 7876 73461 7916
rect 73419 7867 73461 7876
rect 73420 5825 73460 7867
rect 72747 5816 72789 5825
rect 72747 5776 72748 5816
rect 72788 5776 72789 5816
rect 72747 5767 72789 5776
rect 73419 5816 73461 5825
rect 73419 5776 73420 5816
rect 73460 5776 73461 5816
rect 73419 5767 73461 5776
rect 56620 2573 56660 2584
rect 71979 2624 72021 2633
rect 71979 2584 71980 2624
rect 72020 2584 72021 2624
rect 71979 2575 72021 2584
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 54699 2120 54741 2129
rect 54699 2080 54700 2120
rect 54740 2080 54741 2120
rect 54699 2071 54741 2080
rect 55755 2120 55797 2129
rect 55755 2080 55756 2120
rect 55796 2080 55797 2120
rect 55755 2071 55797 2080
rect 53836 1903 53876 1912
rect 54700 1952 54740 2071
rect 54700 1903 54740 1912
rect 55084 1952 55124 1963
rect 55084 1877 55124 1912
rect 72748 1952 72788 5767
rect 72748 1903 72788 1912
rect 74092 1952 74132 13747
rect 75916 13208 75956 13217
rect 76012 13208 76052 13756
rect 76204 13747 76244 13756
rect 76588 13376 76628 13385
rect 76628 13336 76820 13376
rect 76588 13327 76628 13336
rect 76204 13208 76244 13217
rect 75956 13168 76052 13208
rect 76108 13168 76204 13208
rect 75628 13040 75668 13049
rect 75628 12368 75668 13000
rect 75916 12545 75956 13168
rect 75915 12536 75957 12545
rect 75915 12496 75916 12536
rect 75956 12496 75957 12536
rect 75915 12487 75957 12496
rect 76108 12368 76148 13168
rect 76204 13159 76244 13168
rect 76780 13208 76820 13336
rect 76780 13159 76820 13168
rect 77164 13208 77204 13217
rect 76300 13124 76340 13133
rect 76300 12965 76340 13084
rect 76299 12956 76341 12965
rect 76299 12916 76300 12956
rect 76340 12916 76341 12956
rect 76299 12907 76341 12916
rect 77164 12881 77204 13168
rect 77163 12872 77205 12881
rect 77163 12832 77164 12872
rect 77204 12832 77205 12872
rect 77163 12823 77205 12832
rect 77164 12704 77204 12823
rect 77260 12704 77300 12713
rect 77164 12664 77260 12704
rect 77260 12655 77300 12664
rect 77452 12452 77492 15511
rect 78028 13217 78068 27340
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 79756 24632 79796 24641
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 79756 23129 79796 24592
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 79755 23120 79797 23129
rect 79755 23080 79756 23120
rect 79796 23080 79797 23120
rect 79755 23071 79797 23080
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 80715 20096 80757 20105
rect 80715 20056 80716 20096
rect 80756 20056 80757 20096
rect 80715 20047 80757 20056
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 79468 15560 79508 15569
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 79468 14972 79508 15520
rect 79851 15560 79893 15569
rect 79851 15520 79852 15560
rect 79892 15520 79893 15560
rect 79851 15511 79893 15520
rect 80716 15560 80756 20047
rect 80812 17300 80852 27340
rect 80908 19340 80948 31219
rect 81196 27656 81236 32152
rect 81387 32192 81429 32201
rect 81387 32152 81388 32192
rect 81428 32152 81429 32192
rect 81387 32143 81429 32152
rect 81388 31604 81428 32143
rect 81964 32033 82004 33664
rect 82060 32192 82100 34336
rect 82252 33881 82292 35092
rect 82443 34964 82485 34973
rect 82443 34924 82444 34964
rect 82484 34924 82485 34964
rect 82443 34915 82485 34924
rect 82444 34830 82484 34915
rect 83212 34544 83252 36175
rect 91600 36142 91601 36182
rect 91641 36142 91642 36182
rect 91600 36133 91642 36142
rect 82251 33872 82293 33881
rect 82251 33832 82252 33872
rect 82292 33832 82293 33872
rect 82251 33823 82293 33832
rect 83212 33797 83252 34504
rect 83211 33788 83253 33797
rect 83211 33748 83212 33788
rect 83252 33748 83253 33788
rect 83211 33739 83253 33748
rect 81675 32024 81717 32033
rect 81675 31984 81676 32024
rect 81716 31984 81717 32024
rect 81675 31975 81717 31984
rect 81963 32024 82005 32033
rect 81963 31984 81964 32024
rect 82004 31984 82005 32024
rect 81963 31975 82005 31984
rect 81388 31555 81428 31564
rect 81676 31352 81716 31975
rect 81771 31688 81813 31697
rect 81771 31648 81772 31688
rect 81812 31648 81813 31688
rect 81771 31639 81813 31648
rect 81676 31303 81716 31312
rect 81772 31352 81812 31639
rect 82060 31520 82100 32152
rect 81003 21692 81045 21701
rect 81003 21652 81004 21692
rect 81044 21652 81045 21692
rect 81003 21643 81045 21652
rect 81004 20096 81044 21643
rect 81196 20189 81236 27616
rect 81387 27656 81429 27665
rect 81387 27616 81388 27656
rect 81428 27616 81429 27656
rect 81387 27607 81429 27616
rect 81388 27068 81428 27607
rect 81772 27380 81812 31312
rect 81868 31480 82100 31520
rect 82252 33704 82292 33713
rect 81868 30680 81908 31480
rect 82060 31352 82100 31361
rect 82252 31352 82292 33664
rect 83211 32024 83253 32033
rect 83211 31984 83212 32024
rect 83252 31984 83253 32024
rect 83211 31975 83253 31984
rect 83212 31890 83252 31975
rect 83211 31688 83253 31697
rect 83211 31648 83212 31688
rect 83252 31648 83253 31688
rect 83211 31639 83253 31648
rect 82100 31312 82484 31352
rect 82060 31303 82100 31312
rect 81868 30521 81908 30640
rect 82251 30680 82293 30689
rect 82251 30640 82252 30680
rect 82292 30640 82293 30680
rect 82251 30631 82293 30640
rect 82252 30546 82292 30631
rect 81867 30512 81909 30521
rect 81867 30472 81868 30512
rect 81908 30472 81909 30512
rect 81867 30463 81909 30472
rect 82059 30512 82101 30521
rect 82059 30472 82060 30512
rect 82100 30472 82101 30512
rect 82059 30463 82101 30472
rect 82060 27665 82100 30463
rect 82059 27656 82101 27665
rect 82059 27616 82060 27656
rect 82100 27616 82101 27656
rect 82059 27607 82101 27616
rect 82060 27522 82100 27607
rect 82444 27380 82484 31312
rect 82539 30512 82581 30521
rect 82539 30472 82540 30512
rect 82580 30472 82581 30512
rect 82539 30463 82581 30472
rect 82540 30378 82580 30463
rect 83212 27824 83252 31639
rect 83212 27775 83252 27784
rect 83115 27656 83157 27665
rect 83115 27616 83116 27656
rect 83156 27616 83157 27656
rect 83115 27607 83157 27616
rect 97515 27656 97557 27665
rect 97515 27616 97516 27656
rect 97556 27616 97557 27656
rect 97515 27607 97557 27616
rect 81388 27019 81428 27028
rect 81676 27340 81812 27380
rect 82060 27340 82484 27380
rect 81676 26816 81716 27340
rect 81676 26767 81716 26776
rect 81772 26816 81812 26825
rect 81772 24716 81812 26776
rect 81388 24676 81812 24716
rect 82060 26816 82100 27340
rect 81195 20180 81237 20189
rect 81195 20140 81196 20180
rect 81236 20140 81237 20180
rect 81195 20131 81237 20140
rect 81388 20180 81428 24676
rect 81771 24548 81813 24557
rect 81771 24508 81772 24548
rect 81812 24508 81813 24548
rect 81771 24499 81813 24508
rect 81772 24414 81812 24499
rect 82060 21701 82100 26776
rect 81483 21692 81525 21701
rect 81483 21652 81484 21692
rect 81524 21652 81525 21692
rect 81483 21643 81525 21652
rect 82059 21692 82101 21701
rect 82059 21652 82060 21692
rect 82100 21652 82101 21692
rect 82059 21643 82101 21652
rect 81004 20047 81044 20056
rect 81292 20096 81332 20105
rect 81292 19508 81332 20056
rect 81388 20021 81428 20140
rect 81387 20012 81429 20021
rect 81387 19972 81388 20012
rect 81428 19972 81429 20012
rect 81387 19963 81429 19972
rect 81484 19508 81524 21643
rect 81579 20180 81621 20189
rect 81579 20140 81580 20180
rect 81620 20140 81621 20180
rect 81579 20131 81621 20140
rect 82251 20180 82293 20189
rect 82251 20140 82252 20180
rect 82292 20140 82293 20180
rect 82251 20131 82293 20140
rect 81292 19468 81428 19508
rect 81292 19340 81332 19349
rect 80908 19300 81292 19340
rect 81292 19291 81332 19300
rect 80812 17260 80948 17300
rect 80811 15896 80853 15905
rect 80811 15856 80812 15896
rect 80852 15856 80853 15896
rect 80811 15847 80853 15856
rect 80716 15511 80756 15520
rect 79852 15426 79892 15511
rect 80812 15392 80852 15847
rect 80716 15352 80852 15392
rect 80428 14972 80468 14981
rect 79468 14932 80428 14972
rect 80428 14923 80468 14932
rect 80716 14720 80756 15352
rect 80716 14671 80756 14680
rect 80812 14720 80852 14729
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 78027 13208 78069 13217
rect 78027 13168 78028 13208
rect 78068 13168 78069 13208
rect 78027 13159 78069 13168
rect 79852 13208 79892 13217
rect 78028 13074 78068 13159
rect 79468 13124 79508 13133
rect 79180 13040 79220 13049
rect 79180 12965 79220 13000
rect 79179 12956 79221 12965
rect 79179 12916 79180 12956
rect 79220 12916 79221 12956
rect 79179 12907 79221 12916
rect 79084 12536 79124 12547
rect 79180 12536 79220 12907
rect 79468 12713 79508 13084
rect 79852 12881 79892 13168
rect 80715 13208 80757 13217
rect 80715 13168 80716 13208
rect 80756 13168 80757 13208
rect 80715 13159 80757 13168
rect 79851 12872 79893 12881
rect 79851 12832 79852 12872
rect 79892 12832 79893 12872
rect 79851 12823 79893 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 79467 12704 79509 12713
rect 79467 12664 79468 12704
rect 79508 12664 79509 12704
rect 79467 12655 79509 12664
rect 79372 12536 79412 12545
rect 79180 12496 79372 12536
rect 79084 12461 79124 12496
rect 77452 12403 77492 12412
rect 79083 12452 79125 12461
rect 79083 12412 79084 12452
rect 79124 12412 79125 12452
rect 79083 12403 79125 12412
rect 79372 12377 79412 12496
rect 79467 12536 79509 12545
rect 79467 12496 79468 12536
rect 79508 12496 79509 12536
rect 79467 12487 79509 12496
rect 79468 12402 79508 12487
rect 75628 12328 76148 12368
rect 74283 10184 74325 10193
rect 74283 10144 74284 10184
rect 74324 10144 74325 10184
rect 74283 10135 74325 10144
rect 74284 5741 74324 10135
rect 74283 5732 74325 5741
rect 74283 5692 74284 5732
rect 74324 5692 74325 5732
rect 74283 5683 74325 5692
rect 76108 5657 76148 12328
rect 79371 12368 79413 12377
rect 79371 12328 79372 12368
rect 79412 12328 79413 12368
rect 79371 12319 79413 12328
rect 79756 12284 79796 12293
rect 79468 12244 79756 12284
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 79468 11696 79508 12244
rect 79756 12235 79796 12244
rect 79468 11647 79508 11656
rect 79852 11696 79892 12823
rect 79947 12704 79989 12713
rect 79947 12664 79948 12704
rect 79988 12664 79989 12704
rect 79947 12655 79989 12664
rect 80235 12704 80277 12713
rect 80235 12664 80236 12704
rect 80276 12664 80277 12704
rect 80235 12655 80277 12664
rect 80427 12704 80469 12713
rect 80427 12664 80428 12704
rect 80468 12664 80469 12704
rect 80427 12655 80469 12664
rect 79948 12368 79988 12655
rect 80236 12620 80276 12655
rect 80236 12569 80276 12580
rect 80331 12536 80373 12545
rect 80331 12496 80332 12536
rect 80372 12496 80373 12536
rect 80331 12487 80373 12496
rect 80332 12402 80372 12487
rect 79948 12319 79988 12328
rect 79852 11024 79892 11656
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 80140 11024 80180 11033
rect 79852 10984 79988 11024
rect 79852 10772 79892 10781
rect 79468 10732 79852 10772
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 79468 10184 79508 10732
rect 79852 10723 79892 10732
rect 79468 10135 79508 10144
rect 79852 10184 79892 10193
rect 79948 10184 79988 10984
rect 79892 10144 79988 10184
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 79467 6488 79509 6497
rect 79467 6448 79468 6488
rect 79508 6448 79509 6488
rect 79467 6439 79509 6448
rect 79852 6488 79892 10144
rect 80140 9974 80180 10984
rect 80236 11024 80276 11033
rect 80428 11024 80468 12655
rect 80620 12536 80660 12545
rect 80620 12461 80660 12496
rect 80619 12452 80661 12461
rect 80619 12412 80620 12452
rect 80660 12412 80661 12452
rect 80619 12403 80661 12412
rect 80276 10984 80468 11024
rect 80524 11024 80564 11033
rect 80620 11024 80660 12403
rect 80564 10984 80660 11024
rect 80716 11696 80756 13159
rect 80236 10975 80276 10984
rect 80428 10025 80468 10098
rect 80427 10016 80469 10025
rect 80427 9976 80428 10016
rect 80468 9976 80469 10016
rect 80427 9974 80469 9976
rect 80140 9967 80469 9974
rect 80140 9934 80468 9967
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 79468 6354 79508 6439
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 76107 5648 76149 5657
rect 76107 5608 76108 5648
rect 76148 5608 76149 5648
rect 76107 5599 76149 5608
rect 79852 4892 79892 6448
rect 80139 6488 80181 6497
rect 80139 6448 80140 6488
rect 80180 6448 80181 6488
rect 80139 6439 80181 6448
rect 80140 5900 80180 6439
rect 80428 6068 80468 9934
rect 80140 5851 80180 5860
rect 80332 6028 80468 6068
rect 80332 5480 80372 6028
rect 80427 5900 80469 5909
rect 80427 5860 80428 5900
rect 80468 5860 80469 5900
rect 80427 5851 80469 5860
rect 80428 5648 80468 5851
rect 80524 5825 80564 10984
rect 80716 10184 80756 11656
rect 80716 6488 80756 10144
rect 80812 9857 80852 14680
rect 80811 9848 80853 9857
rect 80811 9808 80812 9848
rect 80852 9808 80853 9848
rect 80811 9799 80853 9808
rect 80908 7220 80948 17260
rect 81388 17081 81428 19468
rect 81484 19459 81524 19468
rect 81484 19088 81524 19097
rect 81387 17072 81429 17081
rect 81387 17032 81388 17072
rect 81428 17032 81429 17072
rect 81387 17023 81429 17032
rect 81484 14729 81524 19048
rect 81580 15569 81620 20131
rect 81868 20096 81908 20105
rect 81676 19928 81716 19937
rect 81868 19928 81908 20056
rect 82252 20096 82292 20131
rect 83116 20105 83156 27607
rect 97516 24557 97556 27607
rect 97515 24548 97557 24557
rect 97515 24508 97516 24548
rect 97556 24508 97557 24548
rect 97515 24499 97557 24508
rect 82252 20045 82292 20056
rect 83115 20096 83157 20105
rect 83115 20056 83116 20096
rect 83156 20056 83157 20096
rect 83115 20047 83157 20056
rect 83116 19962 83156 20047
rect 91468 20021 91508 24240
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 84267 20012 84309 20021
rect 84267 19972 84268 20012
rect 84308 19972 84309 20012
rect 84267 19963 84309 19972
rect 91467 20012 91509 20021
rect 91467 19972 91468 20012
rect 91508 19972 91509 20012
rect 91467 19963 91509 19972
rect 81716 19888 81908 19928
rect 81676 19879 81716 19888
rect 84268 19878 84308 19963
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 90776 17240 90818 17249
rect 90776 17200 90777 17240
rect 90817 17200 90818 17240
rect 90776 17191 90818 17200
rect 95384 17240 95426 17249
rect 95384 17200 95385 17240
rect 95425 17200 95426 17240
rect 95384 17191 95426 17200
rect 81867 17072 81909 17081
rect 81867 17032 81868 17072
rect 81908 17032 81909 17072
rect 81867 17023 81909 17032
rect 81868 15905 81908 17023
rect 82731 16988 82773 16997
rect 82731 16948 82732 16988
rect 82772 16948 82773 16988
rect 90777 16979 90817 17191
rect 93848 17156 93890 17165
rect 93848 17116 93849 17156
rect 93889 17116 93890 17156
rect 93848 17107 93890 17116
rect 94232 17156 94274 17165
rect 94232 17116 94233 17156
rect 94273 17116 94274 17156
rect 94232 17107 94274 17116
rect 93849 16979 93889 17107
rect 94233 16979 94273 17107
rect 95000 16988 95042 16997
rect 82731 16939 82773 16948
rect 95000 16948 95001 16988
rect 95041 16948 95042 16988
rect 95385 16979 95425 17191
rect 95000 16939 95042 16948
rect 81963 16820 82005 16829
rect 81963 16780 81964 16820
rect 82004 16780 82005 16820
rect 81963 16771 82005 16780
rect 81867 15896 81909 15905
rect 81867 15856 81868 15896
rect 81908 15856 81909 15896
rect 81867 15847 81909 15856
rect 81868 15728 81908 15847
rect 81868 15679 81908 15688
rect 81579 15560 81621 15569
rect 81579 15520 81580 15560
rect 81620 15520 81621 15560
rect 81579 15511 81621 15520
rect 81099 14720 81141 14729
rect 81099 14680 81100 14720
rect 81140 14680 81141 14720
rect 81099 14671 81141 14680
rect 81483 14720 81525 14729
rect 81483 14680 81484 14720
rect 81524 14680 81525 14720
rect 81483 14671 81525 14680
rect 81100 14586 81140 14671
rect 81868 13460 81908 13469
rect 81964 13460 82004 16771
rect 81908 13420 82004 13460
rect 81868 13411 81908 13420
rect 81868 13040 81908 13049
rect 81868 12713 81908 13000
rect 81867 12704 81909 12713
rect 81867 12664 81868 12704
rect 81908 12664 81909 12704
rect 81867 12655 81909 12664
rect 81867 12536 81909 12545
rect 81867 12496 81868 12536
rect 81908 12496 81909 12536
rect 81867 12487 81909 12496
rect 81868 11780 81908 12487
rect 81868 11537 81908 11740
rect 81867 11528 81909 11537
rect 81867 11488 81868 11528
rect 81908 11488 81909 11528
rect 81867 11479 81909 11488
rect 81868 10268 81908 10277
rect 81868 10025 81908 10228
rect 81867 10016 81909 10025
rect 81867 9976 81868 10016
rect 81908 9976 81909 10016
rect 81867 9967 81909 9976
rect 81867 9848 81909 9857
rect 81867 9808 81868 9848
rect 81908 9808 81909 9848
rect 81867 9799 81909 9808
rect 81868 8849 81908 9799
rect 81867 8840 81909 8849
rect 81867 8800 81868 8840
rect 81908 8800 81909 8840
rect 81867 8791 81909 8800
rect 80716 6439 80756 6448
rect 80812 7180 80948 7220
rect 80523 5816 80565 5825
rect 80812 5816 80852 7180
rect 81868 6656 81908 8791
rect 82732 7925 82772 16939
rect 82731 7916 82773 7925
rect 82731 7876 82732 7916
rect 82772 7876 82773 7916
rect 82731 7867 82773 7876
rect 81868 6607 81908 6616
rect 81868 6236 81908 6245
rect 81868 5909 81908 6196
rect 81867 5900 81909 5909
rect 81867 5860 81868 5900
rect 81908 5860 81909 5900
rect 81867 5851 81909 5860
rect 80523 5776 80524 5816
rect 80564 5776 80565 5816
rect 80523 5767 80565 5776
rect 80716 5776 80852 5816
rect 80428 5599 80468 5608
rect 80524 5648 80564 5657
rect 80564 5608 80660 5648
rect 80524 5599 80564 5608
rect 80523 5480 80565 5489
rect 80332 5440 80468 5480
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 80139 4976 80181 4985
rect 80139 4936 80140 4976
rect 80180 4936 80181 4976
rect 80139 4927 80181 4936
rect 80236 4976 80276 4985
rect 80428 4976 80468 5440
rect 80523 5440 80524 5480
rect 80564 5440 80565 5480
rect 80523 5431 80565 5440
rect 80276 4936 80468 4976
rect 80524 4976 80564 5431
rect 80236 4927 80276 4936
rect 79852 4852 79988 4892
rect 79852 4724 79892 4733
rect 79468 4684 79852 4724
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 79468 4136 79508 4684
rect 79852 4675 79892 4684
rect 79468 4087 79508 4096
rect 79852 4136 79892 4145
rect 79948 4136 79988 4852
rect 80140 4842 80180 4927
rect 79892 4096 79988 4136
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 79852 2624 79892 4096
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 79468 2540 79508 2549
rect 79508 2500 79604 2540
rect 79468 2491 79508 2500
rect 74092 1903 74132 1912
rect 78604 1952 78644 1961
rect 52491 1868 52533 1877
rect 52491 1828 52492 1868
rect 52532 1828 52533 1868
rect 52491 1819 52533 1828
rect 52779 1868 52821 1877
rect 52779 1828 52780 1868
rect 52820 1828 52821 1868
rect 52779 1819 52821 1828
rect 55083 1868 55125 1877
rect 55083 1828 55084 1868
rect 55124 1828 55125 1868
rect 55083 1819 55125 1828
rect 52684 1700 52724 1709
rect 52684 1205 52724 1660
rect 52780 1364 52820 1819
rect 78604 1625 78644 1912
rect 78892 1952 78932 1961
rect 78892 1700 78932 1912
rect 78987 1952 79029 1961
rect 78987 1912 78988 1952
rect 79028 1912 79029 1952
rect 78987 1903 79029 1912
rect 79468 1952 79508 1961
rect 78988 1818 79028 1903
rect 79276 1784 79316 1793
rect 79468 1784 79508 1912
rect 79316 1744 79508 1784
rect 79276 1735 79316 1744
rect 78892 1660 79220 1700
rect 78603 1616 78645 1625
rect 78603 1576 78604 1616
rect 78644 1576 78645 1616
rect 78603 1567 78645 1576
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 79180 1457 79220 1660
rect 79179 1448 79221 1457
rect 79179 1408 79180 1448
rect 79220 1408 79221 1448
rect 79179 1399 79221 1408
rect 52780 1315 52820 1324
rect 79564 1364 79604 2500
rect 79852 1952 79892 2584
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 79852 1903 79892 1912
rect 79947 1952 79989 1961
rect 79947 1912 79948 1952
rect 79988 1912 79989 1952
rect 79947 1903 79989 1912
rect 79948 1541 79988 1903
rect 80524 1625 80564 4936
rect 80235 1616 80277 1625
rect 80235 1576 80236 1616
rect 80276 1576 80277 1616
rect 80235 1567 80277 1576
rect 80523 1616 80565 1625
rect 80523 1576 80524 1616
rect 80564 1576 80565 1616
rect 80523 1567 80565 1576
rect 79947 1532 79989 1541
rect 79947 1492 79948 1532
rect 79988 1492 79989 1532
rect 79947 1483 79989 1492
rect 79564 1315 79604 1324
rect 52491 1196 52533 1205
rect 52491 1156 52492 1196
rect 52532 1156 52533 1196
rect 52491 1147 52533 1156
rect 52683 1196 52725 1205
rect 52683 1156 52684 1196
rect 52724 1156 52725 1196
rect 52683 1147 52725 1156
rect 52108 1063 52148 1072
rect 52396 1063 52436 1072
rect 52492 1112 52532 1147
rect 52492 1061 52532 1072
rect 79948 1112 79988 1483
rect 79948 1063 79988 1072
rect 80236 1112 80276 1567
rect 80236 1063 80276 1072
rect 80620 1037 80660 5608
rect 80716 4136 80756 5776
rect 80812 5648 80852 5657
rect 80812 5489 80852 5608
rect 80811 5480 80853 5489
rect 80811 5440 80812 5480
rect 80852 5440 80853 5480
rect 80811 5431 80853 5440
rect 81867 4976 81909 4985
rect 81867 4936 81868 4976
rect 81908 4936 81909 4976
rect 81867 4927 81909 4936
rect 81868 4388 81908 4927
rect 81868 4339 81908 4348
rect 80716 2717 80756 4096
rect 81868 3968 81908 3977
rect 81908 3928 82100 3968
rect 81868 3919 81908 3928
rect 80715 2708 80757 2717
rect 80715 2668 80716 2708
rect 80756 2668 80757 2708
rect 80715 2659 80757 2668
rect 80716 2624 80756 2659
rect 80716 1952 80756 2584
rect 81868 2456 81908 2465
rect 81908 2416 82004 2456
rect 81868 2407 81908 2416
rect 80716 1903 80756 1912
rect 81868 1700 81908 1709
rect 81868 1541 81908 1660
rect 81867 1532 81909 1541
rect 81867 1492 81868 1532
rect 81908 1492 81909 1532
rect 81867 1483 81909 1492
rect 47307 1028 47349 1037
rect 47307 988 47308 1028
rect 47348 988 47349 1028
rect 47307 979 47349 988
rect 47499 1028 47541 1037
rect 47499 988 47500 1028
rect 47540 988 47541 1028
rect 47499 979 47541 988
rect 79851 1028 79893 1037
rect 79851 988 79852 1028
rect 79892 988 79893 1028
rect 79851 979 79893 988
rect 80619 1028 80661 1037
rect 80619 988 80620 1028
rect 80660 988 80661 1028
rect 80619 979 80661 988
rect 47308 894 47348 979
rect 79852 894 79892 979
rect 38379 860 38421 869
rect 38379 820 38380 860
rect 38420 820 38421 860
rect 38379 811 38421 820
rect 81868 785 81908 1483
rect 81964 1037 82004 2416
rect 82060 1457 82100 3928
rect 82059 1448 82101 1457
rect 82059 1408 82060 1448
rect 82100 1408 82101 1448
rect 82059 1399 82101 1408
rect 81963 1028 82005 1037
rect 81963 988 81964 1028
rect 82004 988 82005 1028
rect 81963 979 82005 988
rect 82060 953 82100 1399
rect 89048 1041 89106 1042
rect 89048 1001 89057 1041
rect 89097 1001 89106 1041
rect 89048 1000 89106 1001
rect 82059 944 82101 953
rect 82059 904 82060 944
rect 82100 904 82101 944
rect 82059 895 82101 904
rect 89260 869 89300 1021
rect 89259 860 89301 869
rect 89259 820 89260 860
rect 89300 820 89301 860
rect 89259 811 89301 820
rect 90777 785 90817 1021
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 81867 776 81909 785
rect 81867 736 81868 776
rect 81908 736 81909 776
rect 81867 727 81909 736
rect 90776 776 90818 785
rect 90776 736 90777 776
rect 90817 736 90818 776
rect 90776 727 90818 736
rect 90988 701 91028 1021
rect 94233 953 94273 1021
rect 94232 944 94274 953
rect 94232 904 94233 944
rect 94273 904 94274 944
rect 94232 895 94274 904
rect 30795 692 30837 701
rect 30795 652 30796 692
rect 30836 652 30837 692
rect 30795 643 30837 652
rect 90987 692 91029 701
rect 90987 652 90988 692
rect 91028 652 91029 692
rect 90987 643 91029 652
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 652 37528 692 37568
rect 268 35848 308 35888
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 5740 36688 5780 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 5548 33832 5588 33872
rect 3532 33664 3572 33704
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 1708 33160 1748 33200
rect 844 32068 884 32108
rect 1420 31900 1460 31940
rect 1900 32068 1940 32108
rect 2092 31900 2132 31940
rect 2956 31900 2996 31940
rect 1612 31396 1652 31436
rect 1900 31396 1940 31436
rect 2764 31396 2804 31436
rect 1516 30724 1556 30764
rect 1132 30220 1172 30260
rect 940 29716 980 29756
rect 748 28876 788 28916
rect 652 26188 692 26228
rect 652 24928 692 24968
rect 1228 29968 1268 30008
rect 1612 30220 1652 30260
rect 2476 30892 2516 30932
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 2092 29884 2132 29924
rect 1804 29800 1844 29840
rect 1612 29716 1652 29756
rect 1228 29128 1268 29168
rect 1420 29128 1460 29168
rect 2092 29296 2132 29336
rect 1612 28960 1652 29000
rect 1516 28876 1556 28916
rect 2572 29800 2612 29840
rect 2668 29716 2708 29756
rect 2956 29716 2996 29756
rect 2476 29212 2516 29252
rect 1900 28960 1940 29000
rect 1996 28708 2036 28748
rect 2188 29128 2228 29168
rect 2380 28708 2420 28748
rect 1420 27448 1460 27488
rect 1036 26104 1076 26144
rect 2092 27616 2132 27656
rect 1996 27448 2036 27488
rect 1996 27280 2036 27320
rect 1228 26104 1268 26144
rect 844 23668 884 23708
rect 652 23248 692 23288
rect 652 23080 692 23120
rect 1516 26776 1556 26816
rect 1612 26188 1652 26228
rect 1900 26776 1940 26816
rect 2380 27616 2420 27656
rect 2764 29296 2804 29336
rect 2956 29296 2996 29336
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 5260 32404 5300 32444
rect 3820 31396 3860 31436
rect 3628 31312 3668 31352
rect 3628 30892 3668 30932
rect 3532 29464 3572 29504
rect 4876 31312 4916 31352
rect 4780 31144 4820 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3820 30220 3860 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3724 29296 3764 29336
rect 2668 29212 2708 29252
rect 3052 29128 3092 29168
rect 3340 29128 3380 29168
rect 3436 28876 3476 28916
rect 2860 28708 2900 28748
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 3148 28540 3188 28580
rect 3532 28540 3572 28580
rect 3916 29128 3956 29168
rect 4492 29128 4532 29168
rect 3628 28456 3668 28496
rect 2860 27616 2900 27656
rect 4396 28876 4436 28916
rect 3916 28456 3956 28496
rect 3436 27532 3476 27572
rect 3052 27448 3092 27488
rect 3628 27448 3668 27488
rect 3532 27364 3572 27404
rect 2668 26776 2708 26816
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3052 26776 3092 26816
rect 1996 25936 2036 25976
rect 2572 26104 2612 26144
rect 2188 25264 2228 25304
rect 1132 24508 1172 24548
rect 1420 24508 1460 24548
rect 1900 24508 1940 24548
rect 1036 24088 1076 24128
rect 1228 23668 1268 23708
rect 1132 23584 1172 23624
rect 1324 23080 1364 23120
rect 1036 22324 1076 22364
rect 652 21568 692 21608
rect 1612 23752 1652 23792
rect 1708 23668 1748 23708
rect 1612 23584 1652 23624
rect 1996 23752 2036 23792
rect 2092 23668 2132 23708
rect 1996 23248 2036 23288
rect 2284 23164 2324 23204
rect 1900 23080 1940 23120
rect 1516 21484 1556 21524
rect 652 20728 692 20768
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 1228 18628 1268 18668
rect 844 18544 884 18584
rect 652 18208 692 18248
rect 1228 17704 1268 17744
rect 652 17368 692 17408
rect 1036 16528 1076 16568
rect 1228 15856 1268 15896
rect 652 15688 692 15728
rect 460 15520 500 15560
rect 1420 17620 1460 17660
rect 1612 18544 1652 18584
rect 2092 20896 2132 20936
rect 2476 20644 2516 20684
rect 1900 18292 1940 18332
rect 3340 26692 3380 26732
rect 3628 26776 3668 26816
rect 4108 28120 4148 28160
rect 4300 28120 4340 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 4588 27616 4628 27656
rect 4204 27364 4244 27404
rect 4588 27364 4628 27404
rect 4108 27280 4148 27320
rect 4300 27280 4340 27320
rect 3820 26608 3860 26648
rect 3724 26524 3764 26564
rect 3532 26104 3572 26144
rect 4012 26776 4052 26816
rect 4684 27028 4724 27068
rect 4300 26692 4340 26732
rect 4204 26608 4244 26648
rect 4492 26608 4532 26648
rect 4108 26524 4148 26564
rect 3724 26188 3764 26228
rect 3436 26020 3476 26060
rect 3340 25936 3380 25976
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3916 26188 3956 26228
rect 4684 26272 4724 26312
rect 2956 25096 2996 25136
rect 3340 24592 3380 24632
rect 3436 24424 3476 24464
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 3724 25096 3764 25136
rect 4108 25852 4148 25892
rect 4012 25264 4052 25304
rect 3916 24592 3956 24632
rect 3724 24508 3764 24548
rect 4492 26104 4532 26144
rect 4300 25852 4340 25892
rect 4684 25264 4724 25304
rect 4492 25096 4532 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 4396 24760 4436 24800
rect 4108 24424 4148 24464
rect 4204 24340 4244 24380
rect 3052 23248 3092 23288
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 4396 23248 4436 23288
rect 4588 23164 4628 23204
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 3532 21568 3572 21608
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4684 23080 4724 23120
rect 3820 21568 3860 21608
rect 2764 20644 2804 20684
rect 2860 20560 2900 20600
rect 3148 20056 3188 20096
rect 4588 22996 4628 23036
rect 4204 22828 4244 22868
rect 4972 27616 5012 27656
rect 4876 26104 4916 26144
rect 4876 25852 4916 25892
rect 4972 25264 5012 25304
rect 4972 24424 5012 24464
rect 4780 22828 4820 22868
rect 4108 20896 4148 20936
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 4684 21736 4724 21776
rect 4300 21652 4340 21692
rect 4396 21568 4436 21608
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3436 19972 3476 20012
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4780 20056 4820 20096
rect 4300 19972 4340 20012
rect 4588 19552 4628 19592
rect 4684 19048 4724 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 5260 24508 5300 24548
rect 5068 23080 5108 23120
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 83212 36184 83252 36224
rect 12172 35848 12212 35888
rect 12460 35848 12500 35888
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 13324 34336 13364 34376
rect 5932 34168 5972 34208
rect 14380 34168 14420 34208
rect 13324 33832 13364 33872
rect 11116 33664 11156 33704
rect 5932 33160 5972 33200
rect 5740 32992 5780 33032
rect 9292 33076 9332 33116
rect 7084 32992 7124 33032
rect 7276 32992 7316 33032
rect 7084 32824 7124 32864
rect 6604 32656 6644 32696
rect 5740 32488 5780 32528
rect 6028 31816 6068 31856
rect 5452 30220 5492 30260
rect 5836 29128 5876 29168
rect 5836 27028 5876 27068
rect 5932 26188 5972 26228
rect 5836 25096 5876 25136
rect 5740 24508 5780 24548
rect 4972 21568 5012 21608
rect 5260 20560 5300 20600
rect 4972 20056 5012 20096
rect 4972 19048 5012 19088
rect 4588 18712 4628 18752
rect 3820 18628 3860 18668
rect 2860 18292 2900 18332
rect 3244 18292 3284 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4012 18292 4052 18332
rect 1804 17620 1844 17660
rect 2284 17704 2324 17744
rect 2668 17620 2708 17660
rect 1420 16024 1460 16064
rect 844 15436 884 15476
rect 652 14848 692 14888
rect 652 14008 692 14048
rect 1228 14512 1268 14552
rect 1516 15520 1556 15560
rect 1900 16192 1940 16232
rect 1900 15940 1940 15980
rect 1708 15604 1748 15644
rect 1132 13672 1172 13712
rect 1420 13672 1460 13712
rect 844 13588 884 13628
rect 652 13168 692 13208
rect 844 13000 884 13040
rect 1420 13504 1460 13544
rect 652 12328 692 12368
rect 556 11488 596 11528
rect 652 9808 692 9848
rect 1804 15520 1844 15560
rect 2092 16192 2132 16232
rect 2284 16024 2324 16064
rect 2284 15856 2324 15896
rect 2092 15604 2132 15644
rect 1996 15520 2036 15560
rect 2092 15436 2132 15476
rect 2092 14680 2132 14720
rect 1708 13672 1748 13712
rect 1900 13588 1940 13628
rect 1804 13504 1844 13544
rect 1516 13000 1556 13040
rect 1996 13000 2036 13040
rect 1708 12496 1748 12536
rect 1612 11824 1652 11864
rect 940 11236 980 11276
rect 1612 11236 1652 11276
rect 844 10900 884 10940
rect 844 10060 884 10100
rect 1708 11152 1748 11192
rect 1036 10732 1076 10772
rect 1420 10900 1460 10940
rect 1228 10312 1268 10352
rect 1324 10144 1364 10184
rect 652 8968 692 9008
rect 844 8800 884 8840
rect 652 7288 692 7328
rect 1996 10984 2036 11024
rect 1612 10144 1652 10184
rect 1804 10144 1844 10184
rect 1516 10060 1556 10100
rect 1420 8800 1460 8840
rect 2188 14428 2228 14468
rect 2572 15772 2612 15812
rect 2572 14512 2612 14552
rect 2284 13924 2324 13964
rect 2188 12496 2228 12536
rect 2188 10312 2228 10352
rect 2572 13168 2612 13208
rect 4300 17704 4340 17744
rect 4012 17620 4052 17660
rect 4300 17536 4340 17576
rect 2764 16780 2804 16820
rect 2764 15856 2804 15896
rect 2476 11824 2516 11864
rect 1900 8884 1940 8924
rect 1036 8128 1076 8168
rect 940 7120 980 7160
rect 556 7036 596 7076
rect 652 6448 692 6488
rect 2380 8884 2420 8924
rect 652 5608 692 5648
rect 1228 5608 1268 5648
rect 268 5524 308 5564
rect 652 4768 692 4808
rect 652 3928 692 3968
rect 1708 8464 1748 8504
rect 1612 7120 1652 7160
rect 1516 5104 1556 5144
rect 1900 7036 1940 7076
rect 1708 3676 1748 3716
rect 1420 3592 1460 3632
rect 2284 7120 2324 7160
rect 2092 7036 2132 7076
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4876 17704 4916 17744
rect 5068 18712 5108 18752
rect 4972 17536 5012 17576
rect 5932 21652 5972 21692
rect 5836 19972 5876 20012
rect 5836 17536 5876 17576
rect 4972 17284 5012 17324
rect 5740 17284 5780 17324
rect 6412 31060 6452 31100
rect 6892 31228 6932 31268
rect 6604 27616 6644 27656
rect 6412 22996 6452 23036
rect 6028 19972 6068 20012
rect 6028 19552 6068 19592
rect 3244 17032 3284 17072
rect 4780 17032 4820 17072
rect 3052 16780 3092 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4396 16528 4436 16568
rect 3628 15856 3668 15896
rect 3532 15436 3572 15476
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4396 16192 4436 16232
rect 3820 15940 3860 15980
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4492 15604 4532 15644
rect 4588 15520 4628 15560
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4972 15604 5012 15644
rect 4684 14680 4724 14720
rect 3820 14512 3860 14552
rect 3436 12328 3476 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3436 10816 3476 10856
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3916 14092 3956 14132
rect 4012 14008 4052 14048
rect 4204 14008 4244 14048
rect 4012 13420 4052 13460
rect 3628 12916 3668 12956
rect 3820 12916 3860 12956
rect 3916 12328 3956 12368
rect 4300 13924 4340 13964
rect 4684 13168 4724 13208
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3724 10816 3764 10856
rect 4588 11488 4628 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 4012 11236 4052 11276
rect 4204 11236 4244 11276
rect 4396 10984 4436 11024
rect 4588 10984 4628 11024
rect 4108 10900 4148 10940
rect 4108 10564 4148 10604
rect 3820 10312 3860 10352
rect 3244 10144 3284 10184
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 5932 15100 5972 15140
rect 5836 14512 5876 14552
rect 5836 14092 5876 14132
rect 5932 14008 5972 14048
rect 4876 11488 4916 11528
rect 4972 11404 5012 11444
rect 4876 10984 4916 11024
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 4396 9472 4436 9512
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4108 8632 4148 8672
rect 4780 8632 4820 8672
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 4684 7960 4724 8000
rect 3820 7120 3860 7160
rect 4204 7036 4244 7076
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 5836 11320 5876 11360
rect 5260 11068 5300 11108
rect 4972 9472 5012 9512
rect 4876 7960 4916 8000
rect 4876 7036 4916 7076
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 4492 5020 4532 5060
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 2956 4180 2996 4220
rect 4588 4096 4628 4136
rect 2572 4012 2612 4052
rect 2476 3844 2516 3884
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 1996 3256 2036 3296
rect 652 3088 692 3128
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 5836 10900 5876 10940
rect 6604 15520 6644 15560
rect 6028 10564 6068 10604
rect 5260 8884 5300 8924
rect 5932 7120 5972 7160
rect 4972 5692 5012 5732
rect 5836 5692 5876 5732
rect 6604 5860 6644 5900
rect 5932 5356 5972 5396
rect 4972 5020 5012 5060
rect 4780 2836 4820 2876
rect 7276 32656 7316 32696
rect 8908 32488 8948 32528
rect 7756 32404 7796 32444
rect 7948 32320 7988 32360
rect 7852 31732 7892 31772
rect 7660 15285 7700 15325
rect 7660 14512 7700 14552
rect 7564 10732 7604 10772
rect 7564 10144 7604 10184
rect 7852 8632 7892 8672
rect 7660 5608 7700 5648
rect 9196 31816 9236 31856
rect 8236 30976 8276 31016
rect 7948 5440 7988 5480
rect 12268 33076 12308 33116
rect 13996 33076 14036 33116
rect 14476 33076 14516 33116
rect 12268 32656 12308 32696
rect 14092 32656 14132 32696
rect 14188 32572 14228 32612
rect 13804 32488 13844 32528
rect 32620 35008 32660 35048
rect 15052 34336 15092 34376
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 20812 34504 20852 34544
rect 21580 34504 21620 34544
rect 22732 34504 22772 34544
rect 25324 34504 25364 34544
rect 15244 33832 15284 33872
rect 15244 33664 15284 33704
rect 14860 33580 14900 33620
rect 14860 33328 14900 33368
rect 15820 34168 15860 34208
rect 16684 34168 16724 34208
rect 16012 33832 16052 33872
rect 16972 33832 17012 33872
rect 15724 33748 15764 33788
rect 17356 33748 17396 33788
rect 16972 33580 17012 33620
rect 16396 33076 16436 33116
rect 15148 32656 15188 32696
rect 14668 31732 14708 31772
rect 11116 31312 11156 31352
rect 17260 33076 17300 33116
rect 16396 32572 16436 32612
rect 16300 32488 16340 32528
rect 15628 32236 15668 32276
rect 18412 34084 18452 34124
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 17644 33076 17684 33116
rect 19276 34168 19316 34208
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 20428 33748 20468 33788
rect 20620 33580 20660 33620
rect 20428 33496 20468 33536
rect 19372 33412 19412 33452
rect 19276 33076 19316 33116
rect 18796 32656 18836 32696
rect 17548 32488 17588 32528
rect 17452 32236 17492 32276
rect 18028 32236 18068 32276
rect 20524 33076 20564 33116
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 22348 34336 22388 34376
rect 21100 33748 21140 33788
rect 22060 34168 22100 34208
rect 21772 34000 21812 34040
rect 21388 33832 21428 33872
rect 21580 33832 21620 33872
rect 21196 33580 21236 33620
rect 21004 33076 21044 33116
rect 20812 31900 20852 31940
rect 22348 33748 22388 33788
rect 22636 33748 22676 33788
rect 21964 33412 22004 33452
rect 22444 33412 22484 33452
rect 23116 34420 23156 34460
rect 23692 34336 23732 34376
rect 23020 33580 23060 33620
rect 22924 33412 22964 33452
rect 22828 33328 22868 33368
rect 23020 32404 23060 32444
rect 21196 31228 21236 31268
rect 24940 33832 24980 33872
rect 24076 33748 24116 33788
rect 25804 34420 25844 34460
rect 27820 34168 27860 34208
rect 25804 34084 25844 34124
rect 25612 34000 25652 34040
rect 27532 33832 27572 33872
rect 23980 33496 24020 33536
rect 23116 30976 23156 31016
rect 25516 33412 25556 33452
rect 26572 33412 26612 33452
rect 27532 33160 27572 33200
rect 25708 32656 25748 32696
rect 27436 32488 27476 32528
rect 28396 33664 28436 33704
rect 31468 34336 31508 34376
rect 32716 34336 32756 34376
rect 29644 34168 29684 34208
rect 29644 33916 29684 33956
rect 30220 33916 30260 33956
rect 30604 33664 30644 33704
rect 29260 33496 29300 33536
rect 30508 33496 30548 33536
rect 33004 35008 33044 35048
rect 32812 34168 32852 34208
rect 30604 33412 30644 33452
rect 30220 33328 30260 33368
rect 29740 33160 29780 33200
rect 29644 32488 29684 32528
rect 27532 31144 27572 31184
rect 29548 31144 29588 31184
rect 31564 33664 31604 33704
rect 31468 33160 31508 33200
rect 31756 33496 31796 33536
rect 32332 33412 32372 33452
rect 10252 30220 10292 30260
rect 18233 30052 18273 30092
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 33100 33916 33140 33956
rect 33484 33664 33524 33704
rect 34060 35008 34100 35048
rect 33772 34084 33812 34124
rect 33772 33916 33812 33956
rect 34156 33748 34196 33788
rect 34060 33664 34100 33704
rect 33580 33412 33620 33452
rect 34156 33328 34196 33368
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 34732 35008 34772 35048
rect 34252 33076 34292 33116
rect 33100 32992 33140 33032
rect 33964 32656 34004 32696
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 35692 34336 35732 34376
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 34444 33664 34484 33704
rect 35308 33664 35348 33704
rect 35692 33664 35732 33704
rect 37900 34168 37940 34208
rect 37708 33748 37748 33788
rect 36940 33580 36980 33620
rect 35596 33412 35636 33452
rect 36556 33412 36596 33452
rect 36748 33076 36788 33116
rect 37708 33412 37748 33452
rect 37324 32824 37364 32864
rect 49996 34504 50036 34544
rect 81196 34924 81236 34964
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 42124 34420 42164 34460
rect 38188 34168 38228 34208
rect 38476 34084 38516 34124
rect 38476 33832 38516 33872
rect 38284 33664 38324 33704
rect 38860 34336 38900 34376
rect 40588 34336 40628 34376
rect 38860 33916 38900 33956
rect 40300 33832 40340 33872
rect 39148 33664 39188 33704
rect 38572 33160 38612 33200
rect 38092 32656 38132 32696
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 34444 32404 34484 32444
rect 34252 32320 34292 32360
rect 42124 33832 42164 33872
rect 40876 33412 40916 33452
rect 42028 33580 42068 33620
rect 42892 33664 42932 33704
rect 42316 33580 42356 33620
rect 43084 32992 43124 33032
rect 45292 33580 45332 33620
rect 40972 32824 41012 32864
rect 44044 32824 44084 32864
rect 44716 32824 44756 32864
rect 42700 32656 42740 32696
rect 45388 32656 45428 32696
rect 44044 32488 44084 32528
rect 49324 34336 49364 34376
rect 45580 33160 45620 33200
rect 47308 33244 47348 33284
rect 48748 33664 48788 33704
rect 47884 33580 47924 33620
rect 49708 34252 49748 34292
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 50092 33748 50132 33788
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 47980 33160 48020 33200
rect 45964 32656 46004 32696
rect 46156 32656 46196 32696
rect 45676 32572 45716 32612
rect 47500 32572 47540 32612
rect 47596 32404 47636 32444
rect 45964 32236 46004 32276
rect 47884 32236 47924 32276
rect 45484 31228 45524 31268
rect 38764 30892 38804 30932
rect 49132 32992 49172 33032
rect 51532 34336 51572 34376
rect 51820 34336 51860 34376
rect 50764 33664 50804 33704
rect 51340 33664 51380 33704
rect 50476 33580 50516 33620
rect 50284 32992 50324 33032
rect 49900 32656 49940 32696
rect 50764 32992 50804 33032
rect 49324 32572 49364 32612
rect 50572 32572 50612 32612
rect 48940 32488 48980 32528
rect 48652 31060 48692 31100
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 51820 33664 51860 33704
rect 52492 34252 52532 34292
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 52684 33664 52724 33704
rect 71980 33664 72020 33704
rect 53164 33580 53204 33620
rect 52492 33412 52532 33452
rect 52972 33412 53012 33452
rect 52300 32572 52340 32612
rect 51628 32404 51668 32444
rect 51532 32236 51572 32276
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 65932 33160 65972 33200
rect 65548 32992 65588 33032
rect 65932 32824 65972 32864
rect 66124 32824 66164 32864
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 65548 32488 65588 32528
rect 53740 32404 53780 32444
rect 54316 32404 54356 32444
rect 70060 32908 70100 32948
rect 69772 32740 69812 32780
rect 70060 32572 70100 32612
rect 66124 32488 66164 32528
rect 65740 31648 65780 31688
rect 14188 4180 14228 4220
rect 13324 4096 13364 4136
rect 12940 4012 12980 4052
rect 8236 3928 8276 3968
rect 7084 3424 7124 3464
rect 16204 4096 16244 4136
rect 14188 3760 14228 3800
rect 12940 3004 12980 3044
rect 17260 3760 17300 3800
rect 17452 3760 17492 3800
rect 18700 3760 18740 3800
rect 19276 3760 19316 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 20332 3760 20372 3800
rect 13228 2920 13268 2960
rect 15052 2836 15092 2876
rect 17260 3088 17300 3128
rect 17356 2920 17396 2960
rect 17548 2920 17588 2960
rect 6892 2668 6932 2708
rect 17260 2584 17300 2624
rect 21292 3928 21332 3968
rect 22156 3928 22196 3968
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 19948 2920 19988 2960
rect 18124 2836 18164 2876
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 18124 1912 18164 1952
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 18700 1492 18740 1532
rect 19756 1912 19796 1952
rect 19948 1828 19988 1868
rect 20524 3088 20564 3128
rect 22060 3760 22100 3800
rect 21292 3004 21332 3044
rect 20716 2920 20756 2960
rect 23212 3928 23252 3968
rect 22828 3760 22868 3800
rect 22060 2920 22100 2960
rect 20044 1492 20084 1532
rect 20428 1492 20468 1532
rect 21388 1912 21428 1952
rect 21772 1912 21812 1952
rect 22156 1912 22196 1952
rect 22540 2920 22580 2960
rect 22540 1996 22580 2036
rect 23116 2584 23156 2624
rect 23404 3088 23444 3128
rect 23404 2668 23444 2708
rect 23788 5356 23828 5396
rect 26332 5860 26372 5900
rect 31084 5692 31124 5732
rect 31708 5692 31748 5732
rect 25708 5524 25748 5564
rect 23980 4012 24020 4052
rect 25036 3928 25076 3968
rect 25132 2668 25172 2708
rect 23884 2584 23924 2624
rect 28396 3928 28436 3968
rect 29452 3928 29492 3968
rect 27148 2836 27188 2876
rect 26860 2668 26900 2708
rect 25516 2500 25556 2540
rect 23212 2332 23252 2372
rect 23500 2416 23540 2456
rect 25420 2416 25460 2456
rect 23404 1996 23444 2036
rect 26476 2416 26516 2456
rect 24460 2332 24500 2372
rect 26380 2332 26420 2372
rect 23116 1912 23156 1952
rect 25036 1996 25076 2036
rect 25324 1912 25364 1952
rect 28588 2752 28628 2792
rect 28396 2668 28436 2708
rect 27244 2584 27284 2624
rect 28396 2500 28436 2540
rect 28108 2416 28148 2456
rect 27244 1828 27284 1868
rect 28396 2164 28436 2204
rect 28972 2584 29012 2624
rect 29164 2416 29204 2456
rect 28972 1912 29012 1952
rect 28684 1324 28724 1364
rect 23884 1072 23924 1112
rect 25324 1072 25364 1112
rect 30892 3844 30932 3884
rect 30028 2584 30068 2624
rect 30700 2416 30740 2456
rect 30124 2332 30164 2372
rect 29740 2080 29780 2120
rect 30124 1828 30164 1868
rect 29836 1324 29876 1364
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 30988 3676 31028 3716
rect 33388 5440 33428 5480
rect 33772 5440 33812 5480
rect 31180 5020 31220 5060
rect 33292 4096 33332 4136
rect 31180 3844 31220 3884
rect 33676 3928 33716 3968
rect 30892 3172 30932 3212
rect 32236 3004 32276 3044
rect 32044 2920 32084 2960
rect 31276 2836 31316 2876
rect 31180 2752 31220 2792
rect 32716 3088 32756 3128
rect 32620 2668 32660 2708
rect 31468 2500 31508 2540
rect 31660 2080 31700 2120
rect 31564 1996 31604 2036
rect 31468 1912 31508 1952
rect 34252 4684 34292 4724
rect 34156 3676 34196 3716
rect 33964 3592 34004 3632
rect 34444 4096 34484 4136
rect 34732 4684 34772 4724
rect 35020 4096 35060 4136
rect 34348 3844 34388 3884
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 34060 3172 34100 3212
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 33868 3004 33908 3044
rect 33196 2668 33236 2708
rect 34828 3592 34868 3632
rect 34636 2920 34676 2960
rect 34924 3088 34964 3128
rect 35020 3004 35060 3044
rect 34828 2752 34868 2792
rect 35212 3592 35252 3632
rect 35212 3088 35252 3128
rect 35308 2752 35348 2792
rect 35116 2332 35156 2372
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 34444 2080 34484 2120
rect 35980 2920 36020 2960
rect 35788 2752 35828 2792
rect 34828 1996 34868 2036
rect 35500 1996 35540 2036
rect 33388 1912 33428 1952
rect 34060 1912 34100 1952
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 35692 1996 35732 2036
rect 35404 1828 35444 1868
rect 32716 1324 32756 1364
rect 35308 1324 35348 1364
rect 35980 1912 36020 1952
rect 36172 2668 36212 2708
rect 36844 5188 36884 5228
rect 36652 5020 36692 5060
rect 37324 5104 37364 5144
rect 36940 4684 36980 4724
rect 37516 4936 37556 4976
rect 37420 4684 37460 4724
rect 37036 3844 37076 3884
rect 37228 3592 37268 3632
rect 37612 3844 37652 3884
rect 39340 3592 39380 3632
rect 37996 3256 38036 3296
rect 36748 3172 36788 3212
rect 37324 3172 37364 3212
rect 38092 3172 38132 3212
rect 38188 3004 38228 3044
rect 37996 2836 38036 2876
rect 36844 2668 36884 2708
rect 37036 2584 37076 2624
rect 36844 2248 36884 2288
rect 37228 1828 37268 1868
rect 36556 1408 36596 1448
rect 37900 1240 37940 1280
rect 36076 1156 36116 1196
rect 35788 1072 35828 1112
rect 37900 1072 37940 1112
rect 38092 2500 38132 2540
rect 38092 2248 38132 2288
rect 38284 1156 38324 1196
rect 39244 2836 39284 2876
rect 39340 2500 39380 2540
rect 38956 1996 38996 2036
rect 39628 2920 39668 2960
rect 39724 2836 39764 2876
rect 39820 2164 39860 2204
rect 40889 5860 40929 5900
rect 40300 3592 40340 3632
rect 39820 1492 39860 1532
rect 39628 1156 39668 1196
rect 40204 1996 40244 2036
rect 40684 4936 40724 4976
rect 42700 3424 42740 3464
rect 41260 2920 41300 2960
rect 40876 2668 40916 2708
rect 40876 2500 40916 2540
rect 40588 2164 40628 2204
rect 40012 1324 40052 1364
rect 39916 1240 39956 1280
rect 42412 2920 42452 2960
rect 41356 2836 41396 2876
rect 42796 2668 42836 2708
rect 41644 2164 41684 2204
rect 42124 2164 42164 2204
rect 41740 1996 41780 2036
rect 41548 1324 41588 1364
rect 41932 1744 41972 1784
rect 42700 2164 42740 2204
rect 44908 3592 44948 3632
rect 44524 3340 44564 3380
rect 43084 2752 43124 2792
rect 43276 2668 43316 2708
rect 44140 2500 44180 2540
rect 43276 1996 43316 2036
rect 47308 3760 47348 3800
rect 47116 3676 47156 3716
rect 46444 3508 46484 3548
rect 46924 3508 46964 3548
rect 45004 2500 45044 2540
rect 45676 2752 45716 2792
rect 45292 2500 45332 2540
rect 45196 2080 45236 2120
rect 44428 1996 44468 2036
rect 44524 1744 44564 1784
rect 42988 1492 43028 1532
rect 42892 1324 42932 1364
rect 42412 1072 42452 1112
rect 44428 1072 44468 1112
rect 39532 988 39572 1028
rect 45100 1324 45140 1364
rect 46348 3004 46388 3044
rect 46060 2668 46100 2708
rect 46924 2500 46964 2540
rect 47116 2500 47156 2540
rect 47212 1408 47252 1448
rect 45964 1072 46004 1112
rect 46924 1072 46964 1112
rect 47308 1324 47348 1364
rect 48940 3928 48980 3968
rect 48652 3676 48692 3716
rect 52396 3844 52436 3884
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 52300 3760 52340 3800
rect 47596 3592 47636 3632
rect 48748 3592 48788 3632
rect 49612 3676 49652 3716
rect 51820 3676 51860 3716
rect 49036 3508 49076 3548
rect 52204 3592 52244 3632
rect 52108 3508 52148 3548
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 47980 2752 48020 2792
rect 48652 2752 48692 2792
rect 49516 2500 49556 2540
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 54604 3676 54644 3716
rect 57772 3676 57812 3716
rect 52396 3508 52436 3548
rect 52300 2920 52340 2960
rect 50860 2752 50900 2792
rect 51244 2752 51284 2792
rect 49996 2500 50036 2540
rect 47404 1156 47444 1196
rect 44716 988 44756 1028
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 47596 1324 47636 1364
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 52108 2500 52148 2540
rect 50284 1828 50324 1868
rect 49996 1408 50036 1448
rect 49900 1324 49940 1364
rect 49612 1240 49652 1280
rect 49900 1156 49940 1196
rect 54892 3592 54932 3632
rect 55180 3592 55220 3632
rect 54988 3508 55028 3548
rect 53836 2668 53876 2708
rect 54028 2668 54068 2708
rect 53164 2500 53204 2540
rect 55756 2836 55796 2876
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 56620 2668 56660 2708
rect 80812 33496 80852 33536
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 80716 32740 80756 32780
rect 78508 32572 78548 32612
rect 74188 30892 74228 30932
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 78508 30640 78548 30680
rect 78700 30640 78740 30680
rect 78316 30388 78356 30428
rect 78892 30388 78932 30428
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 80812 32152 80852 32192
rect 81868 33748 81908 33788
rect 81580 33496 81620 33536
rect 80908 31228 80948 31268
rect 80812 27616 80852 27656
rect 75628 23080 75668 23120
rect 77452 15520 77492 15560
rect 76396 14680 76436 14720
rect 74092 13756 74132 13796
rect 75628 13756 75668 13796
rect 73420 7876 73460 7916
rect 72748 5776 72788 5816
rect 73420 5776 73460 5816
rect 71980 2584 72020 2624
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 54700 2080 54740 2120
rect 55756 2080 55796 2120
rect 75916 12496 75956 12536
rect 76300 12916 76340 12956
rect 77164 12832 77204 12872
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 79756 23080 79796 23120
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 80716 20056 80756 20096
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 79852 15520 79892 15560
rect 81388 32152 81428 32192
rect 82444 34924 82484 34964
rect 91601 36142 91641 36182
rect 82252 33832 82292 33872
rect 83212 33748 83252 33788
rect 81676 31984 81716 32024
rect 81964 31984 82004 32024
rect 81772 31648 81812 31688
rect 81004 21652 81044 21692
rect 81388 27616 81428 27656
rect 83212 31984 83252 32024
rect 83212 31648 83252 31688
rect 82252 30640 82292 30680
rect 81868 30472 81908 30512
rect 82060 30472 82100 30512
rect 82060 27616 82100 27656
rect 82540 30472 82580 30512
rect 83116 27616 83156 27656
rect 97516 27616 97556 27656
rect 81196 20140 81236 20180
rect 81772 24508 81812 24548
rect 81484 21652 81524 21692
rect 82060 21652 82100 21692
rect 81388 19972 81428 20012
rect 81580 20140 81620 20180
rect 82252 20140 82292 20180
rect 80812 15856 80852 15896
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 78028 13168 78068 13208
rect 79180 12916 79220 12956
rect 80716 13168 80756 13208
rect 79852 12832 79892 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 79468 12664 79508 12704
rect 79084 12412 79124 12452
rect 79468 12496 79508 12536
rect 74284 10144 74324 10184
rect 74284 5692 74324 5732
rect 79372 12328 79412 12368
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 79948 12664 79988 12704
rect 80236 12664 80276 12704
rect 80428 12664 80468 12704
rect 80332 12496 80372 12536
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 79468 6448 79508 6488
rect 80620 12412 80660 12452
rect 80428 9976 80468 10016
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 76108 5608 76148 5648
rect 80140 6448 80180 6488
rect 80428 5860 80468 5900
rect 80812 9808 80852 9848
rect 81388 17032 81428 17072
rect 97516 24508 97556 24548
rect 83116 20056 83156 20096
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 84268 19972 84308 20012
rect 91468 19972 91508 20012
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 90777 17200 90817 17240
rect 95385 17200 95425 17240
rect 81868 17032 81908 17072
rect 82732 16948 82772 16988
rect 93849 17116 93889 17156
rect 94233 17116 94273 17156
rect 95001 16948 95041 16988
rect 81964 16780 82004 16820
rect 81868 15856 81908 15896
rect 81580 15520 81620 15560
rect 81100 14680 81140 14720
rect 81484 14680 81524 14720
rect 81868 12664 81908 12704
rect 81868 12496 81908 12536
rect 81868 11488 81908 11528
rect 81868 9976 81908 10016
rect 81868 9808 81908 9848
rect 81868 8800 81908 8840
rect 82732 7876 82772 7916
rect 81868 5860 81908 5900
rect 80524 5776 80564 5816
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 80140 4936 80180 4976
rect 80524 5440 80564 5480
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 52492 1828 52532 1868
rect 52780 1828 52820 1868
rect 55084 1828 55124 1868
rect 78988 1912 79028 1952
rect 78604 1576 78644 1616
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 79180 1408 79220 1448
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 79948 1912 79988 1952
rect 80236 1576 80276 1616
rect 80524 1576 80564 1616
rect 79948 1492 79988 1532
rect 52492 1156 52532 1196
rect 52684 1156 52724 1196
rect 80812 5440 80852 5480
rect 81868 4936 81908 4976
rect 80716 2668 80756 2708
rect 81868 1492 81908 1532
rect 47308 988 47348 1028
rect 47500 988 47540 1028
rect 79852 988 79892 1028
rect 80620 988 80660 1028
rect 38380 820 38420 860
rect 82060 1408 82100 1448
rect 81964 988 82004 1028
rect 89057 1001 89097 1041
rect 82060 904 82100 944
rect 89260 820 89300 860
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 81868 736 81908 776
rect 90777 736 90817 776
rect 94233 904 94273 944
rect 30796 652 30836 692
rect 90988 652 91028 692
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 0 37568 80 37588
rect 0 37528 652 37568
rect 692 37528 701 37568
rect 0 37508 80 37528
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 0 36728 80 36748
rect 0 36688 5740 36728
rect 5780 36688 5789 36728
rect 0 36668 80 36688
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 83203 36184 83212 36224
rect 83252 36184 91220 36224
rect 91180 36182 91220 36184
rect 91180 36142 91601 36182
rect 91641 36142 91650 36182
rect 0 35888 80 35908
rect 4771 35888 4829 35889
rect 0 35848 268 35888
rect 308 35848 317 35888
rect 4771 35848 4780 35888
rect 4820 35848 12172 35888
rect 12212 35848 12460 35888
rect 12500 35848 12509 35888
rect 0 35828 80 35848
rect 4771 35847 4829 35848
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 0 34988 80 35068
rect 32611 35008 32620 35048
rect 32660 35008 33004 35048
rect 33044 35008 34060 35048
rect 34100 35008 34732 35048
rect 34772 35008 34781 35048
rect 81187 34924 81196 34964
rect 81236 34924 82444 34964
rect 82484 34924 82493 34964
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 20803 34544 20861 34545
rect 50179 34544 50237 34545
rect 20718 34504 20812 34544
rect 20852 34504 20861 34544
rect 21571 34504 21580 34544
rect 21620 34504 22004 34544
rect 22723 34504 22732 34544
rect 22772 34504 25324 34544
rect 25364 34504 25373 34544
rect 49987 34504 49996 34544
rect 50036 34504 50188 34544
rect 50228 34504 50237 34544
rect 20803 34503 20861 34504
rect 21964 34460 22004 34504
rect 50179 34503 50237 34504
rect 42115 34460 42173 34461
rect 21964 34420 23116 34460
rect 23156 34420 25804 34460
rect 25844 34420 25853 34460
rect 42030 34420 42124 34460
rect 42164 34420 42173 34460
rect 42115 34419 42173 34420
rect 13315 34336 13324 34376
rect 13364 34336 15052 34376
rect 15092 34336 21812 34376
rect 22339 34336 22348 34376
rect 22388 34336 23692 34376
rect 23732 34336 23741 34376
rect 31459 34336 31468 34376
rect 31508 34336 32716 34376
rect 32756 34336 35692 34376
rect 35732 34336 35741 34376
rect 38851 34336 38860 34376
rect 38900 34336 40588 34376
rect 40628 34336 40637 34376
rect 49315 34336 49324 34376
rect 49364 34336 51532 34376
rect 51572 34336 51581 34376
rect 51811 34336 51820 34376
rect 51860 34336 51869 34376
rect 0 34148 80 34228
rect 5923 34168 5932 34208
rect 5972 34168 14380 34208
rect 14420 34168 15820 34208
rect 15860 34168 15869 34208
rect 16675 34168 16684 34208
rect 16724 34168 19276 34208
rect 19316 34168 19325 34208
rect 15820 34124 15860 34168
rect 15820 34084 18412 34124
rect 18452 34084 18461 34124
rect 21772 34040 21812 34336
rect 51820 34292 51860 34336
rect 49699 34252 49708 34292
rect 49748 34252 52492 34292
rect 52532 34252 52541 34292
rect 22051 34168 22060 34208
rect 22100 34168 27820 34208
rect 27860 34168 29644 34208
rect 29684 34168 29693 34208
rect 32803 34168 32812 34208
rect 32852 34168 37460 34208
rect 37891 34168 37900 34208
rect 37940 34168 38188 34208
rect 38228 34168 38237 34208
rect 37420 34124 37460 34168
rect 25795 34084 25804 34124
rect 25844 34084 33772 34124
rect 33812 34084 33821 34124
rect 37420 34084 38476 34124
rect 38516 34084 38525 34124
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 21763 34000 21772 34040
rect 21812 34000 25612 34040
rect 25652 34000 25661 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 29635 33916 29644 33956
rect 29684 33916 30220 33956
rect 30260 33916 33100 33956
rect 33140 33916 33772 33956
rect 33812 33916 38860 33956
rect 38900 33916 38909 33956
rect 5539 33832 5548 33872
rect 5588 33832 13324 33872
rect 13364 33832 13373 33872
rect 15235 33832 15244 33872
rect 15284 33832 16012 33872
rect 16052 33832 16972 33872
rect 17012 33832 17021 33872
rect 21379 33832 21388 33872
rect 21428 33832 21580 33872
rect 21620 33832 24940 33872
rect 24980 33832 27532 33872
rect 27572 33832 27581 33872
rect 38467 33832 38476 33872
rect 38516 33832 40300 33872
rect 40340 33832 40349 33872
rect 42115 33832 42124 33872
rect 42164 33832 82252 33872
rect 82292 33832 82301 33872
rect 50179 33788 50237 33789
rect 15715 33748 15724 33788
rect 15764 33748 17356 33788
rect 17396 33748 20428 33788
rect 20468 33748 20477 33788
rect 21091 33748 21100 33788
rect 21140 33748 22348 33788
rect 22388 33748 22397 33788
rect 22627 33748 22636 33788
rect 22676 33748 24076 33788
rect 24116 33748 28436 33788
rect 34147 33748 34156 33788
rect 34196 33748 37708 33788
rect 37748 33748 37757 33788
rect 50083 33748 50092 33788
rect 50132 33748 50188 33788
rect 50228 33748 50237 33788
rect 81859 33748 81868 33788
rect 81908 33748 83212 33788
rect 83252 33748 83261 33788
rect 28396 33704 28436 33748
rect 50179 33747 50237 33748
rect 3523 33664 3532 33704
rect 3572 33664 7220 33704
rect 11107 33664 11116 33704
rect 11156 33664 15244 33704
rect 15284 33664 27380 33704
rect 28387 33664 28396 33704
rect 28436 33664 28445 33704
rect 30595 33664 30604 33704
rect 30644 33664 31564 33704
rect 31604 33664 33484 33704
rect 33524 33664 34060 33704
rect 34100 33664 34109 33704
rect 34435 33664 34444 33704
rect 34484 33664 35308 33704
rect 35348 33664 35357 33704
rect 35683 33664 35692 33704
rect 35732 33664 38284 33704
rect 38324 33664 38333 33704
rect 39139 33664 39148 33704
rect 39188 33664 42892 33704
rect 42932 33664 48748 33704
rect 48788 33664 50764 33704
rect 50804 33664 51340 33704
rect 51380 33664 51389 33704
rect 51811 33664 51820 33704
rect 51860 33664 52684 33704
rect 52724 33664 71980 33704
rect 72020 33664 72029 33704
rect 7180 33620 7220 33664
rect 27340 33620 27380 33664
rect 51340 33620 51380 33664
rect 7180 33580 14860 33620
rect 14900 33580 14909 33620
rect 16963 33580 16972 33620
rect 17012 33580 20620 33620
rect 20660 33580 20669 33620
rect 21187 33580 21196 33620
rect 21236 33580 23020 33620
rect 23060 33580 23069 33620
rect 27340 33580 36940 33620
rect 36980 33580 36989 33620
rect 42019 33580 42028 33620
rect 42068 33580 42316 33620
rect 42356 33580 45292 33620
rect 45332 33580 47884 33620
rect 47924 33580 50476 33620
rect 50516 33580 50525 33620
rect 51340 33580 53164 33620
rect 53204 33580 53213 33620
rect 20419 33496 20428 33536
rect 20468 33496 23980 33536
rect 24020 33496 24029 33536
rect 29251 33496 29260 33536
rect 29300 33496 30508 33536
rect 30548 33496 31756 33536
rect 31796 33496 31805 33536
rect 80803 33496 80812 33536
rect 80852 33496 81580 33536
rect 81620 33496 81629 33536
rect 22915 33452 22973 33453
rect 19363 33412 19372 33452
rect 19412 33412 21964 33452
rect 22004 33412 22013 33452
rect 22435 33412 22444 33452
rect 22484 33412 22924 33452
rect 22964 33412 22973 33452
rect 25507 33412 25516 33452
rect 25556 33412 26572 33452
rect 26612 33412 30604 33452
rect 30644 33412 32332 33452
rect 32372 33412 33580 33452
rect 33620 33412 35596 33452
rect 35636 33412 36556 33452
rect 36596 33412 36605 33452
rect 37699 33412 37708 33452
rect 37748 33412 40876 33452
rect 40916 33412 40925 33452
rect 52483 33412 52492 33452
rect 52532 33412 52972 33452
rect 53012 33412 53021 33452
rect 22915 33411 22973 33412
rect 0 33308 80 33388
rect 14851 33328 14860 33368
rect 14900 33328 22828 33368
rect 22868 33328 22877 33368
rect 30211 33328 30220 33368
rect 30260 33328 34156 33368
rect 34196 33328 34205 33368
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 47299 33244 47308 33284
rect 47348 33244 47357 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 47308 33200 47348 33244
rect 1699 33160 1708 33200
rect 1748 33160 5932 33200
rect 5972 33160 5981 33200
rect 27523 33160 27532 33200
rect 27572 33160 29740 33200
rect 29780 33160 31468 33200
rect 31508 33160 31517 33200
rect 38563 33160 38572 33200
rect 38612 33160 45580 33200
rect 45620 33160 47980 33200
rect 48020 33160 48029 33200
rect 65923 33160 65932 33200
rect 65972 33160 66356 33200
rect 17443 33116 17501 33117
rect 66316 33116 66356 33160
rect 68803 33116 68861 33117
rect 9283 33076 9292 33116
rect 9332 33076 12268 33116
rect 12308 33076 12317 33116
rect 13987 33076 13996 33116
rect 14036 33076 14476 33116
rect 14516 33076 14525 33116
rect 16387 33076 16396 33116
rect 16436 33076 17260 33116
rect 17300 33076 17452 33116
rect 17492 33076 17501 33116
rect 17635 33076 17644 33116
rect 17684 33076 19276 33116
rect 19316 33076 20524 33116
rect 20564 33076 21004 33116
rect 21044 33076 21053 33116
rect 34243 33076 34252 33116
rect 34292 33076 36748 33116
rect 36788 33076 36797 33116
rect 66316 33076 68812 33116
rect 68852 33076 68861 33116
rect 17443 33075 17501 33076
rect 68803 33075 68861 33076
rect 5731 32992 5740 33032
rect 5780 32992 7084 33032
rect 7124 32992 7133 33032
rect 7267 32992 7276 33032
rect 7316 32992 33100 33032
rect 33140 32992 33149 33032
rect 43075 32992 43084 33032
rect 43124 32992 49132 33032
rect 49172 32992 50284 33032
rect 50324 32992 50764 33032
rect 50804 32992 65548 33032
rect 65588 32992 65597 33032
rect 67660 32908 70060 32948
rect 70100 32908 70109 32948
rect 67660 32864 67700 32908
rect 7075 32824 7084 32864
rect 7124 32824 37324 32864
rect 37364 32824 37373 32864
rect 40963 32824 40972 32864
rect 41012 32824 44044 32864
rect 44084 32824 44093 32864
rect 44707 32824 44716 32864
rect 44756 32824 65932 32864
rect 65972 32824 65981 32864
rect 66115 32824 66124 32864
rect 66164 32824 67700 32864
rect 69763 32740 69772 32780
rect 69812 32740 80716 32780
rect 80756 32740 80765 32780
rect 17443 32696 17501 32697
rect 69091 32696 69149 32697
rect 6595 32656 6604 32696
rect 6644 32656 7276 32696
rect 7316 32656 7325 32696
rect 12259 32656 12268 32696
rect 12308 32656 12980 32696
rect 14083 32656 14092 32696
rect 14132 32656 15148 32696
rect 15188 32656 15197 32696
rect 17443 32656 17452 32696
rect 17492 32656 18796 32696
rect 18836 32656 18845 32696
rect 25699 32656 25708 32696
rect 25748 32656 33964 32696
rect 34004 32656 38092 32696
rect 38132 32656 42700 32696
rect 42740 32656 42749 32696
rect 45379 32656 45388 32696
rect 45428 32656 45964 32696
rect 46004 32656 46013 32696
rect 46147 32656 46156 32696
rect 46196 32656 49900 32696
rect 49940 32656 69100 32696
rect 69140 32656 69149 32696
rect 12940 32612 12980 32656
rect 14092 32612 14132 32656
rect 17443 32655 17501 32656
rect 69091 32655 69149 32656
rect 61987 32612 62045 32613
rect 12940 32572 14132 32612
rect 14179 32572 14188 32612
rect 14228 32572 16396 32612
rect 16436 32572 16445 32612
rect 45667 32572 45676 32612
rect 45716 32572 47500 32612
rect 47540 32572 49324 32612
rect 49364 32572 49373 32612
rect 50563 32572 50572 32612
rect 50612 32572 52300 32612
rect 52340 32572 61996 32612
rect 62036 32572 62045 32612
rect 70051 32572 70060 32612
rect 70100 32572 78508 32612
rect 78548 32572 78557 32612
rect 61987 32571 62045 32572
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 5731 32488 5740 32528
rect 5780 32488 8908 32528
rect 8948 32488 13804 32528
rect 13844 32488 13853 32528
rect 16291 32488 16300 32528
rect 16340 32488 17548 32528
rect 17588 32488 17597 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 27427 32488 27436 32528
rect 27476 32488 29644 32528
rect 29684 32488 29693 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 44035 32488 44044 32528
rect 44084 32488 48940 32528
rect 48980 32488 48989 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 65539 32488 65548 32528
rect 65588 32488 66124 32528
rect 66164 32488 66173 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 16300 32444 16340 32488
rect 5251 32404 5260 32444
rect 5300 32404 7756 32444
rect 7796 32404 16340 32444
rect 23011 32404 23020 32444
rect 23060 32404 34444 32444
rect 34484 32404 34493 32444
rect 47587 32404 47596 32444
rect 47636 32404 51628 32444
rect 51668 32404 53740 32444
rect 53780 32404 54316 32444
rect 54356 32404 54365 32444
rect 7939 32320 7948 32360
rect 7988 32320 34252 32360
rect 34292 32320 34301 32360
rect 4963 32276 5021 32277
rect 66211 32276 66269 32277
rect 4963 32236 4972 32276
rect 5012 32236 15628 32276
rect 15668 32236 17452 32276
rect 17492 32236 18028 32276
rect 18068 32236 18077 32276
rect 45955 32236 45964 32276
rect 46004 32236 47884 32276
rect 47924 32236 51532 32276
rect 51572 32236 66220 32276
rect 66260 32236 66269 32276
rect 4963 32235 5021 32236
rect 66211 32235 66269 32236
rect 80803 32152 80812 32192
rect 80852 32152 81388 32192
rect 81428 32152 81437 32192
rect 835 32068 844 32108
rect 884 32068 1900 32108
rect 1940 32068 1949 32108
rect 81667 31984 81676 32024
rect 81716 31984 81964 32024
rect 82004 31984 83212 32024
rect 83252 31984 85421 32024
rect 1411 31900 1420 31940
rect 1460 31900 2092 31940
rect 2132 31900 2956 31940
rect 2996 31900 20812 31940
rect 20852 31900 20861 31940
rect 6019 31816 6028 31856
rect 6068 31816 9196 31856
rect 9236 31816 9245 31856
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 7843 31732 7852 31772
rect 7892 31732 14668 31772
rect 14708 31732 14717 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 0 31628 80 31708
rect 69283 31688 69341 31689
rect 65731 31648 65740 31688
rect 65780 31648 69292 31688
rect 69332 31648 69341 31688
rect 81763 31648 81772 31688
rect 81812 31648 83212 31688
rect 83252 31648 85421 31688
rect 69283 31647 69341 31648
rect 1603 31396 1612 31436
rect 1652 31396 1900 31436
rect 1940 31396 2764 31436
rect 2804 31396 3820 31436
rect 3860 31396 3869 31436
rect 3619 31312 3628 31352
rect 3668 31312 4876 31352
rect 4916 31312 11116 31352
rect 11156 31312 11165 31352
rect 6883 31228 6892 31268
rect 6932 31228 21196 31268
rect 21236 31228 21245 31268
rect 43180 31228 45484 31268
rect 45524 31228 80908 31268
rect 80948 31228 80957 31268
rect 4771 31144 4780 31184
rect 4820 31144 27532 31184
rect 27572 31144 29548 31184
rect 29588 31144 29597 31184
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 2467 30892 2476 30932
rect 2516 30892 3628 30932
rect 3668 30892 3677 30932
rect 0 30788 80 30868
rect 4780 30764 4820 31144
rect 43180 31100 43220 31228
rect 69187 31100 69245 31101
rect 6403 31060 6412 31100
rect 6452 31060 43220 31100
rect 48643 31060 48652 31100
rect 48692 31060 69196 31100
rect 69236 31060 69245 31100
rect 69187 31059 69245 31060
rect 8227 30976 8236 31016
rect 8276 30976 23116 31016
rect 23156 30976 23165 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 38755 30892 38764 30932
rect 38804 30892 74188 30932
rect 74228 30892 74237 30932
rect 1507 30724 1516 30764
rect 1556 30724 4820 30764
rect 78499 30640 78508 30680
rect 78548 30640 78700 30680
rect 78740 30640 82252 30680
rect 82292 30640 82301 30680
rect 97320 30512 97362 30521
rect 81859 30472 81868 30512
rect 81908 30472 82060 30512
rect 82100 30472 82540 30512
rect 82580 30472 82589 30512
rect 97320 30472 97321 30512
rect 97361 30472 97362 30512
rect 97320 30463 97362 30472
rect 78307 30388 78316 30428
rect 78356 30388 78892 30428
rect 78932 30388 78941 30428
rect 1123 30220 1132 30260
rect 1172 30220 1612 30260
rect 1652 30220 1661 30260
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 3811 30220 3820 30260
rect 3860 30220 5452 30260
rect 5492 30220 10252 30260
rect 10292 30220 10301 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 7843 30092 7901 30093
rect 22915 30092 22973 30093
rect 7843 30052 7852 30092
rect 7892 30052 18233 30092
rect 18273 30052 22924 30092
rect 22964 30052 22973 30092
rect 7843 30051 7901 30052
rect 22915 30051 22973 30052
rect 0 29948 80 30028
rect 1219 29968 1228 30008
rect 1268 29968 2132 30008
rect 2092 29924 2132 29968
rect 2083 29884 2092 29924
rect 2132 29884 2141 29924
rect 1795 29800 1804 29840
rect 1844 29800 2572 29840
rect 2612 29800 2621 29840
rect 931 29716 940 29756
rect 980 29716 1612 29756
rect 1652 29716 1661 29756
rect 2659 29716 2668 29756
rect 2708 29716 2956 29756
rect 2996 29716 3005 29756
rect 3523 29504 3581 29505
rect 3438 29464 3532 29504
rect 3572 29464 3581 29504
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 3523 29463 3581 29464
rect 2083 29296 2092 29336
rect 2132 29296 2764 29336
rect 2804 29296 2813 29336
rect 2947 29296 2956 29336
rect 2996 29296 3724 29336
rect 3764 29296 3773 29336
rect 2467 29212 2476 29252
rect 2516 29212 2668 29252
rect 2708 29212 3380 29252
rect 0 29108 80 29188
rect 3340 29168 3380 29212
rect 1219 29128 1228 29168
rect 1268 29128 1420 29168
rect 1460 29128 2188 29168
rect 2228 29128 2237 29168
rect 2860 29128 3052 29168
rect 3092 29128 3101 29168
rect 3331 29128 3340 29168
rect 3380 29128 3389 29168
rect 3907 29128 3916 29168
rect 3956 29128 4492 29168
rect 4532 29128 5836 29168
rect 5876 29128 5885 29168
rect 2188 29084 2228 29128
rect 2860 29084 2900 29128
rect 2188 29044 2900 29084
rect 1603 28960 1612 29000
rect 1652 28960 1900 29000
rect 1940 28960 1949 29000
rect 739 28876 748 28916
rect 788 28876 1516 28916
rect 1556 28876 1565 28916
rect 3427 28876 3436 28916
rect 3476 28876 4396 28916
rect 4436 28876 4445 28916
rect 1987 28708 1996 28748
rect 2036 28708 2380 28748
rect 2420 28708 2860 28748
rect 2900 28708 2909 28748
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 3139 28540 3148 28580
rect 3188 28540 3532 28580
rect 3572 28540 3581 28580
rect 3619 28456 3628 28496
rect 3668 28456 3916 28496
rect 3956 28456 3965 28496
rect 0 28268 80 28348
rect 4099 28120 4108 28160
rect 4148 28120 4300 28160
rect 4340 28120 4349 28160
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 2083 27616 2092 27656
rect 2132 27616 2380 27656
rect 2420 27616 2860 27656
rect 2900 27616 2909 27656
rect 4579 27616 4588 27656
rect 4628 27616 4972 27656
rect 5012 27616 6604 27656
rect 6644 27616 6653 27656
rect 80803 27616 80812 27656
rect 80852 27616 81388 27656
rect 81428 27616 81437 27656
rect 82051 27616 82060 27656
rect 82100 27616 83116 27656
rect 83156 27616 83165 27656
rect 97379 27616 97516 27656
rect 97556 27616 97565 27656
rect 3427 27532 3436 27572
rect 3476 27532 3764 27572
rect 0 27428 80 27508
rect 1411 27448 1420 27488
rect 1460 27448 1996 27488
rect 2036 27448 2045 27488
rect 3043 27448 3052 27488
rect 3092 27448 3628 27488
rect 3668 27448 3677 27488
rect 3523 27364 3532 27404
rect 3572 27364 3581 27404
rect 3532 27320 3572 27364
rect 1987 27280 1996 27320
rect 2036 27280 3572 27320
rect 3724 27320 3764 27532
rect 4195 27364 4204 27404
rect 4244 27364 4588 27404
rect 4628 27364 4637 27404
rect 3724 27280 4108 27320
rect 4148 27280 4300 27320
rect 4340 27280 4349 27320
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 4675 27028 4684 27068
rect 4724 27028 5836 27068
rect 5876 27028 5885 27068
rect 1507 26776 1516 26816
rect 1556 26776 1900 26816
rect 1940 26776 2668 26816
rect 2708 26776 3052 26816
rect 3092 26776 3101 26816
rect 3619 26776 3628 26816
rect 3668 26776 4012 26816
rect 4052 26776 4061 26816
rect 3331 26692 3340 26732
rect 3380 26692 4300 26732
rect 4340 26692 4820 26732
rect 0 26588 80 26668
rect 3811 26608 3820 26648
rect 3860 26608 4204 26648
rect 4244 26608 4492 26648
rect 4532 26608 4541 26648
rect 3715 26524 3724 26564
rect 3764 26524 4108 26564
rect 4148 26524 4157 26564
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 4780 26396 4820 26692
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 4684 26356 4820 26396
rect 4684 26312 4724 26356
rect 4675 26272 4684 26312
rect 4724 26272 4733 26312
rect 4195 26228 4253 26229
rect 643 26188 652 26228
rect 692 26188 1612 26228
rect 1652 26188 1661 26228
rect 2476 26188 3724 26228
rect 3764 26188 3773 26228
rect 3907 26188 3916 26228
rect 3956 26188 4204 26228
rect 4244 26188 5932 26228
rect 5972 26188 5981 26228
rect 2476 26144 2516 26188
rect 4195 26187 4253 26188
rect 1027 26104 1036 26144
rect 1076 26104 1228 26144
rect 1268 26104 2516 26144
rect 2563 26104 2572 26144
rect 2612 26104 3532 26144
rect 3572 26104 3581 26144
rect 4483 26104 4492 26144
rect 4532 26104 4876 26144
rect 4916 26104 4925 26144
rect 3427 26020 3436 26060
rect 3476 26020 3485 26060
rect 3436 25976 3476 26020
rect 1987 25936 1996 25976
rect 2036 25936 3340 25976
rect 3380 25936 3389 25976
rect 3436 25936 4916 25976
rect 4876 25892 4916 25936
rect 4099 25852 4108 25892
rect 4148 25852 4300 25892
rect 4340 25852 4349 25892
rect 4867 25852 4876 25892
rect 4916 25852 4925 25892
rect 0 25748 80 25828
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 2179 25264 2188 25304
rect 2228 25264 4012 25304
rect 4052 25264 4684 25304
rect 4724 25264 4972 25304
rect 5012 25264 5021 25304
rect 2947 25096 2956 25136
rect 2996 25096 3724 25136
rect 3764 25096 3773 25136
rect 4483 25096 4492 25136
rect 4532 25096 5836 25136
rect 5876 25096 5885 25136
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 0 24908 80 24928
rect 4780 24884 4820 25096
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 4396 24844 4820 24884
rect 4396 24800 4436 24844
rect 4387 24760 4396 24800
rect 4436 24760 4445 24800
rect 3331 24592 3340 24632
rect 3380 24592 3916 24632
rect 3956 24592 3965 24632
rect 1123 24508 1132 24548
rect 1172 24508 1420 24548
rect 1460 24508 1900 24548
rect 1940 24508 1949 24548
rect 3715 24508 3724 24548
rect 3764 24508 5260 24548
rect 5300 24508 5309 24548
rect 5731 24508 5740 24548
rect 5780 24508 8040 24548
rect 81763 24508 81772 24548
rect 81812 24508 97516 24548
rect 97556 24508 97565 24548
rect 4963 24464 5021 24465
rect 3427 24424 3436 24464
rect 3476 24424 4108 24464
rect 4148 24424 4157 24464
rect 4878 24424 4972 24464
rect 5012 24424 5021 24464
rect 4963 24423 5021 24424
rect 3523 24380 3581 24381
rect 3523 24340 3532 24380
rect 3572 24340 4204 24380
rect 4244 24340 4253 24380
rect 3523 24339 3581 24340
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 0 24128 80 24148
rect 0 24088 1036 24128
rect 1076 24088 1085 24128
rect 0 24068 80 24088
rect 1603 23752 1612 23792
rect 1652 23752 1996 23792
rect 2036 23752 2045 23792
rect 835 23668 844 23708
rect 884 23668 1228 23708
rect 1268 23668 1708 23708
rect 1748 23668 2092 23708
rect 2132 23668 2141 23708
rect 1123 23584 1132 23624
rect 1172 23584 1612 23624
rect 1652 23584 1661 23624
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 0 23288 80 23308
rect 4195 23288 4253 23289
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 1987 23248 1996 23288
rect 2036 23248 3052 23288
rect 3092 23248 3101 23288
rect 4195 23248 4204 23288
rect 4244 23248 4396 23288
rect 4436 23248 4445 23288
rect 0 23228 80 23248
rect 4195 23247 4253 23248
rect 2275 23164 2284 23204
rect 2324 23164 4588 23204
rect 4628 23164 4637 23204
rect 643 23080 652 23120
rect 692 23080 1324 23120
rect 1364 23080 1373 23120
rect 1891 23080 1900 23120
rect 1940 23080 4684 23120
rect 4724 23080 5068 23120
rect 5108 23080 5117 23120
rect 75619 23080 75628 23120
rect 75668 23080 79756 23120
rect 79796 23080 79805 23120
rect 4579 22996 4588 23036
rect 4628 22996 6412 23036
rect 6452 22996 6461 23036
rect 4195 22828 4204 22868
rect 4244 22828 4780 22868
rect 4820 22828 4829 22868
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 0 22448 80 22468
rect 0 22408 1076 22448
rect 0 22388 80 22408
rect 1036 22364 1076 22408
rect 1027 22324 1036 22364
rect 1076 22324 1085 22364
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 4195 21776 4253 21777
rect 4195 21736 4204 21776
rect 4244 21736 4684 21776
rect 4724 21736 4733 21776
rect 4195 21735 4253 21736
rect 4291 21652 4300 21692
rect 4340 21652 5932 21692
rect 5972 21652 5981 21692
rect 80995 21652 81004 21692
rect 81044 21652 81484 21692
rect 81524 21652 82060 21692
rect 82100 21652 82109 21692
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 3523 21568 3532 21608
rect 3572 21568 3820 21608
rect 3860 21568 3869 21608
rect 4387 21568 4396 21608
rect 4436 21568 4972 21608
rect 5012 21568 5021 21608
rect 0 21548 80 21568
rect 6403 21524 6461 21525
rect 1507 21484 1516 21524
rect 1556 21484 6412 21524
rect 6452 21484 6461 21524
rect 6403 21483 6461 21484
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 2083 20896 2092 20936
rect 2132 20896 4108 20936
rect 4148 20896 4157 20936
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 0 20708 80 20728
rect 2467 20644 2476 20684
rect 2516 20644 2764 20684
rect 2804 20644 2813 20684
rect 2851 20560 2860 20600
rect 2900 20560 5260 20600
rect 5300 20571 7604 20600
rect 5300 20560 8021 20571
rect 7564 20531 8021 20560
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 81187 20140 81196 20180
rect 81236 20140 81580 20180
rect 81620 20140 82252 20180
rect 82292 20140 82301 20180
rect 3139 20056 3148 20096
rect 3188 20056 4780 20096
rect 4820 20056 4972 20096
rect 5012 20056 5021 20096
rect 80707 20056 80716 20096
rect 80756 20056 83116 20096
rect 83156 20056 83165 20096
rect 3427 19972 3436 20012
rect 3476 19972 4300 20012
rect 4340 19972 4349 20012
rect 5827 19972 5836 20012
rect 5876 19972 6028 20012
rect 6068 19972 6077 20012
rect 81379 19972 81388 20012
rect 81428 19972 84268 20012
rect 84308 19972 91468 20012
rect 91508 19972 91517 20012
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 0 19868 80 19888
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 4579 19552 4588 19592
rect 4628 19552 6028 19592
rect 6068 19563 7604 19592
rect 6068 19552 8021 19563
rect 7564 19523 8021 19552
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 4675 19048 4684 19088
rect 4724 19048 4972 19088
rect 5012 19048 5021 19088
rect 0 19028 80 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 4579 18712 4588 18752
rect 4628 18712 5068 18752
rect 5108 18712 5117 18752
rect 1219 18628 1228 18668
rect 1268 18628 3820 18668
rect 3860 18628 3869 18668
rect 835 18544 844 18584
rect 884 18544 1612 18584
rect 1652 18544 1661 18584
rect 1891 18292 1900 18332
rect 1940 18292 2860 18332
rect 2900 18292 3244 18332
rect 3284 18292 4012 18332
rect 4052 18292 4061 18332
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 1219 17704 1228 17744
rect 1268 17704 2284 17744
rect 2324 17704 2333 17744
rect 4291 17704 4300 17744
rect 4340 17704 4876 17744
rect 4916 17704 4925 17744
rect 1411 17620 1420 17660
rect 1460 17620 1804 17660
rect 1844 17620 2668 17660
rect 2708 17620 2717 17660
rect 4003 17620 4012 17660
rect 4052 17620 8040 17660
rect 4291 17536 4300 17576
rect 4340 17536 4972 17576
rect 5012 17536 5836 17576
rect 5876 17547 7604 17576
rect 5876 17536 8021 17547
rect 7564 17507 8021 17536
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 0 17348 80 17368
rect 4963 17284 4972 17324
rect 5012 17284 5740 17324
rect 5780 17284 5789 17324
rect 76963 17240 77021 17241
rect 76963 17200 76972 17240
rect 77012 17200 90777 17240
rect 90817 17200 90826 17240
rect 90892 17200 95385 17240
rect 95425 17200 95434 17240
rect 76963 17199 77021 17200
rect 82915 17156 82973 17157
rect 90892 17156 90932 17200
rect 82915 17116 82924 17156
rect 82964 17116 90932 17156
rect 91075 17156 91133 17157
rect 91075 17116 91084 17156
rect 91124 17116 93849 17156
rect 93889 17116 93898 17156
rect 93964 17116 94233 17156
rect 94273 17116 94282 17156
rect 82915 17115 82973 17116
rect 91075 17115 91133 17116
rect 93964 17072 94004 17116
rect 3235 17032 3244 17072
rect 3284 17032 4780 17072
rect 4820 17032 4829 17072
rect 81379 17032 81388 17072
rect 81428 17032 81868 17072
rect 81908 17032 94004 17072
rect 82723 16948 82732 16988
rect 82772 16948 95001 16988
rect 95041 16948 95050 16988
rect 91075 16820 91133 16821
rect 2755 16780 2764 16820
rect 2804 16780 3052 16820
rect 3092 16780 3101 16820
rect 81955 16780 81964 16820
rect 82004 16780 91084 16820
rect 91124 16780 91133 16820
rect 91075 16779 91133 16780
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 0 16568 80 16588
rect 0 16528 1036 16568
rect 1076 16528 1085 16568
rect 4387 16528 4396 16568
rect 4436 16539 7604 16568
rect 4436 16528 8021 16539
rect 0 16508 80 16528
rect 7564 16499 8021 16528
rect 1891 16192 1900 16232
rect 1940 16192 2092 16232
rect 2132 16192 4396 16232
rect 4436 16192 4445 16232
rect 1411 16024 1420 16064
rect 1460 16024 2284 16064
rect 2324 16024 2333 16064
rect 1900 15980 1940 16024
rect 1891 15940 1900 15980
rect 1940 15940 1980 15980
rect 3811 15940 3820 15980
rect 3860 15940 3869 15980
rect 1219 15856 1228 15896
rect 1268 15856 2284 15896
rect 2324 15856 2333 15896
rect 2755 15856 2764 15896
rect 2804 15856 3628 15896
rect 3668 15856 3677 15896
rect 3820 15812 3860 15940
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 80803 15856 80812 15896
rect 80852 15856 81868 15896
rect 81908 15856 81917 15896
rect 2563 15772 2572 15812
rect 2612 15772 3860 15812
rect 0 15728 80 15748
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 0 15668 80 15688
rect 1699 15604 1708 15644
rect 1748 15604 2092 15644
rect 2132 15604 3572 15644
rect 4483 15604 4492 15644
rect 4532 15604 4972 15644
rect 5012 15604 5021 15644
rect 451 15520 460 15560
rect 500 15520 1516 15560
rect 1556 15520 1565 15560
rect 1795 15520 1804 15560
rect 1844 15520 1996 15560
rect 2036 15520 2045 15560
rect 3532 15476 3572 15604
rect 4579 15520 4588 15560
rect 4628 15520 6604 15560
rect 6644 15520 6653 15560
rect 77443 15520 77452 15560
rect 77492 15520 79852 15560
rect 79892 15520 81580 15560
rect 81620 15520 81629 15560
rect 835 15436 844 15476
rect 884 15436 2092 15476
rect 2132 15436 2141 15476
rect 3523 15436 3532 15476
rect 3572 15436 8040 15476
rect 7651 15285 7660 15325
rect 7700 15285 8021 15325
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 5923 15100 5932 15140
rect 5972 15100 8040 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 0 14828 80 14848
rect 2083 14680 2092 14720
rect 2132 14680 4684 14720
rect 4724 14680 4733 14720
rect 76387 14680 76396 14720
rect 76436 14680 81100 14720
rect 81140 14680 81484 14720
rect 81524 14680 81533 14720
rect 1219 14512 1228 14552
rect 1268 14512 2572 14552
rect 2612 14512 3820 14552
rect 3860 14512 3869 14552
rect 5827 14512 5836 14552
rect 5876 14512 7660 14552
rect 7700 14512 7709 14552
rect 6403 14468 6461 14469
rect 2179 14428 2188 14468
rect 2228 14428 6412 14468
rect 6452 14428 6461 14468
rect 6403 14427 6461 14428
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 3907 14092 3916 14132
rect 3956 14092 5836 14132
rect 5876 14092 5885 14132
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 4003 14008 4012 14048
rect 4052 14008 4204 14048
rect 4244 14008 5932 14048
rect 5972 14008 5981 14048
rect 0 13988 80 14008
rect 2275 13924 2284 13964
rect 2324 13924 4300 13964
rect 4340 13924 4349 13964
rect 74083 13756 74092 13796
rect 74132 13756 75628 13796
rect 75668 13756 75677 13796
rect 1123 13672 1132 13712
rect 1172 13672 1420 13712
rect 1460 13672 1708 13712
rect 1748 13672 1757 13712
rect 835 13588 844 13628
rect 884 13588 1900 13628
rect 1940 13588 1949 13628
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 1411 13504 1420 13544
rect 1460 13504 1804 13544
rect 1844 13504 4052 13544
rect 4012 13460 4052 13504
rect 4003 13420 4012 13460
rect 4052 13420 8040 13460
rect 0 13208 80 13228
rect 4771 13208 4829 13209
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 2563 13168 2572 13208
rect 2612 13168 4684 13208
rect 4724 13168 4780 13208
rect 4820 13168 4829 13208
rect 78019 13168 78028 13208
rect 78068 13168 80716 13208
rect 80756 13168 80765 13208
rect 0 13148 80 13168
rect 4771 13167 4829 13168
rect 6595 13040 6653 13041
rect 835 13000 844 13040
rect 884 13000 1516 13040
rect 1556 13000 1565 13040
rect 1987 13000 1996 13040
rect 2036 13000 6604 13040
rect 6644 13000 6653 13040
rect 6595 12999 6653 13000
rect 3619 12916 3628 12956
rect 3668 12916 3820 12956
rect 3860 12916 3869 12956
rect 76291 12916 76300 12956
rect 76340 12916 79180 12956
rect 79220 12916 79229 12956
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 77155 12832 77164 12872
rect 77204 12832 79852 12872
rect 79892 12832 79901 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 79459 12664 79468 12704
rect 79508 12664 79948 12704
rect 79988 12664 79997 12704
rect 80227 12664 80236 12704
rect 80276 12664 80428 12704
rect 80468 12664 81868 12704
rect 81908 12664 81917 12704
rect 1699 12496 1708 12536
rect 1748 12496 2188 12536
rect 2228 12496 2237 12536
rect 75907 12496 75916 12536
rect 75956 12496 75965 12536
rect 79459 12496 79468 12536
rect 79508 12496 80332 12536
rect 80372 12496 81868 12536
rect 81908 12496 81917 12536
rect 75916 12452 75956 12496
rect 75916 12412 79084 12452
rect 79124 12412 80620 12452
rect 80660 12412 80669 12452
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 3427 12328 3436 12368
rect 3476 12328 3916 12368
rect 3956 12328 3965 12368
rect 79363 12328 79372 12368
rect 79412 12328 84021 12368
rect 0 12308 80 12328
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 1603 11824 1612 11864
rect 1652 11824 2476 11864
rect 2516 11824 2525 11864
rect 0 11528 80 11548
rect 0 11488 556 11528
rect 596 11488 605 11528
rect 4579 11488 4588 11528
rect 4628 11488 4876 11528
rect 4916 11488 4925 11528
rect 81859 11488 81868 11528
rect 81908 11488 84021 11528
rect 99931 11501 99989 11502
rect 0 11468 80 11488
rect 99931 11461 99940 11501
rect 99980 11461 99989 11501
rect 99931 11460 99989 11461
rect 4963 11404 4972 11444
rect 5012 11404 8040 11444
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 5827 11320 5836 11360
rect 5876 11331 7604 11360
rect 5876 11320 8021 11331
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 5836 11276 5876 11320
rect 7564 11291 8021 11320
rect 931 11236 940 11276
rect 980 11236 1612 11276
rect 1652 11236 1661 11276
rect 4003 11236 4012 11276
rect 4052 11236 4204 11276
rect 4244 11236 5876 11276
rect 1795 11192 1853 11193
rect 1699 11152 1708 11192
rect 1748 11152 1804 11192
rect 1844 11152 1853 11192
rect 1795 11151 1853 11152
rect 5251 11068 5260 11108
rect 5300 11068 8040 11108
rect 1987 10984 1996 11024
rect 2036 10984 4396 11024
rect 4436 10984 4588 11024
rect 4628 10984 4876 11024
rect 4916 10984 4925 11024
rect 835 10900 844 10940
rect 884 10900 1420 10940
rect 1460 10900 1469 10940
rect 4099 10900 4108 10940
rect 4148 10900 5836 10940
rect 5876 10900 8040 10940
rect 3427 10816 3436 10856
rect 3476 10816 3724 10856
rect 3764 10816 3773 10856
rect 1027 10732 1036 10772
rect 1076 10732 1085 10772
rect 7555 10732 7564 10772
rect 7604 10732 8040 10772
rect 0 10688 80 10708
rect 1036 10688 1076 10732
rect 0 10648 1076 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 4099 10564 4108 10604
rect 4148 10564 6028 10604
rect 6068 10564 8040 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 1219 10312 1228 10352
rect 1268 10312 2188 10352
rect 2228 10312 3820 10352
rect 3860 10312 3869 10352
rect 1315 10144 1324 10184
rect 1364 10144 1612 10184
rect 1652 10144 1661 10184
rect 1795 10144 1804 10184
rect 1844 10144 3244 10184
rect 3284 10144 7564 10184
rect 7604 10144 7613 10184
rect 74275 10144 74284 10184
rect 74324 10144 84021 10184
rect 835 10060 844 10100
rect 884 10060 1516 10100
rect 1556 10060 1565 10100
rect 80419 9976 80428 10016
rect 80468 9976 81868 10016
rect 81908 9976 84021 10016
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 80803 9808 80812 9848
rect 80852 9808 81868 9848
rect 81908 9808 81917 9848
rect 0 9788 80 9808
rect 4387 9472 4396 9512
rect 4436 9472 4972 9512
rect 5012 9472 5021 9512
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 0 9008 80 9028
rect 99920 9008 99962 9017
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 99920 8968 99921 9008
rect 99961 8968 99962 9008
rect 0 8948 80 8968
rect 99920 8959 99962 8968
rect 1891 8884 1900 8924
rect 1940 8884 2380 8924
rect 2420 8884 5260 8924
rect 5300 8884 5309 8924
rect 83491 8840 83549 8841
rect 835 8800 844 8840
rect 884 8800 1420 8840
rect 1460 8800 1469 8840
rect 81859 8800 81868 8840
rect 81908 8800 83500 8840
rect 83540 8800 83549 8840
rect 83491 8799 83549 8800
rect 99931 8813 99989 8814
rect 99931 8773 99940 8813
rect 99980 8773 99989 8813
rect 99931 8772 99989 8773
rect 4099 8632 4108 8672
rect 4148 8632 4780 8672
rect 4820 8632 7852 8672
rect 7892 8632 7901 8672
rect 1699 8504 1757 8505
rect 1614 8464 1708 8504
rect 1748 8464 1757 8504
rect 1699 8463 1757 8464
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 0 8168 80 8188
rect 0 8128 1036 8168
rect 1076 8128 1085 8168
rect 0 8108 80 8128
rect 4675 7960 4684 8000
rect 4724 7960 4876 8000
rect 4916 7960 4925 8000
rect 73411 7876 73420 7916
rect 73460 7876 82732 7916
rect 82772 7876 82781 7916
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 0 7268 80 7288
rect 931 7120 940 7160
rect 980 7120 1612 7160
rect 1652 7120 1661 7160
rect 2275 7120 2284 7160
rect 2324 7120 3820 7160
rect 3860 7120 5932 7160
rect 5972 7120 5981 7160
rect 547 7036 556 7076
rect 596 7036 1900 7076
rect 1940 7036 1949 7076
rect 2083 7036 2092 7076
rect 2132 7036 4204 7076
rect 4244 7036 4876 7076
rect 4916 7036 4925 7076
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 79459 6448 79468 6488
rect 79508 6448 80140 6488
rect 80180 6448 80189 6488
rect 0 6428 80 6448
rect 99931 6293 99989 6294
rect 99931 6253 99940 6293
rect 99980 6253 99989 6293
rect 99931 6252 99989 6253
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 7180 5944 27380 5984
rect 7180 5900 7220 5944
rect 26851 5900 26909 5901
rect 6595 5860 6604 5900
rect 6644 5860 7220 5900
rect 26323 5860 26332 5900
rect 26372 5860 26860 5900
rect 26900 5860 26909 5900
rect 27340 5900 27380 5944
rect 27340 5860 40889 5900
rect 40929 5860 40938 5900
rect 80419 5860 80428 5900
rect 80468 5860 81868 5900
rect 81908 5860 81917 5900
rect 26851 5859 26909 5860
rect 72739 5816 72797 5817
rect 72654 5776 72748 5816
rect 72788 5776 73420 5816
rect 73460 5776 73469 5816
rect 80515 5776 80524 5816
rect 80564 5776 80573 5816
rect 72739 5775 72797 5776
rect 4963 5692 4972 5732
rect 5012 5692 5836 5732
rect 5876 5692 5885 5732
rect 7180 5692 31028 5732
rect 31075 5692 31084 5732
rect 31124 5692 31708 5732
rect 31748 5692 31757 5732
rect 31852 5692 74284 5732
rect 74324 5692 74333 5732
rect 0 5648 80 5668
rect 7180 5648 7220 5692
rect 30988 5648 31028 5692
rect 31852 5648 31892 5692
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 1219 5608 1228 5648
rect 1268 5608 7220 5648
rect 7651 5608 7660 5648
rect 7700 5608 27380 5648
rect 30988 5608 31892 5648
rect 37420 5608 76108 5648
rect 76148 5608 76157 5648
rect 0 5588 80 5608
rect 27340 5564 27380 5608
rect 37420 5564 37460 5608
rect 259 5524 268 5564
rect 308 5524 25708 5564
rect 25748 5524 25757 5564
rect 27340 5524 37460 5564
rect 80524 5480 80564 5776
rect 7939 5440 7948 5480
rect 7988 5440 33388 5480
rect 33428 5440 33772 5480
rect 33812 5440 33821 5480
rect 80515 5440 80524 5480
rect 80564 5440 80812 5480
rect 80852 5440 80861 5480
rect 5923 5356 5932 5396
rect 5972 5356 23788 5396
rect 23828 5356 23837 5396
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 6595 5228 6653 5229
rect 6595 5188 6604 5228
rect 6644 5188 36844 5228
rect 36884 5188 36893 5228
rect 6595 5187 6653 5188
rect 6403 5144 6461 5145
rect 1507 5104 1516 5144
rect 1556 5104 5108 5144
rect 5068 5060 5108 5104
rect 6403 5104 6412 5144
rect 6452 5104 37324 5144
rect 37364 5104 37373 5144
rect 6403 5103 6461 5104
rect 73027 5060 73085 5061
rect 4483 5020 4492 5060
rect 4532 5020 4972 5060
rect 5012 5020 5021 5060
rect 5068 5020 31180 5060
rect 31220 5020 31229 5060
rect 36643 5020 36652 5060
rect 36692 5020 73036 5060
rect 73076 5020 73085 5060
rect 73027 5019 73085 5020
rect 37507 4936 37516 4976
rect 37556 4936 40684 4976
rect 40724 4936 40733 4976
rect 80131 4936 80140 4976
rect 80180 4936 81868 4976
rect 81908 4936 81917 4976
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 34243 4684 34252 4724
rect 34292 4684 34732 4724
rect 34772 4684 34781 4724
rect 36931 4684 36940 4724
rect 36980 4684 37420 4724
rect 37460 4684 37469 4724
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 2947 4180 2956 4220
rect 2996 4180 14188 4220
rect 14228 4180 14237 4220
rect 4579 4096 4588 4136
rect 4628 4096 13324 4136
rect 13364 4096 16204 4136
rect 16244 4096 17300 4136
rect 33283 4096 33292 4136
rect 33332 4096 34444 4136
rect 34484 4096 35020 4136
rect 35060 4096 35069 4136
rect 17260 4052 17300 4096
rect 2563 4012 2572 4052
rect 2612 4012 12940 4052
rect 12980 4012 12989 4052
rect 17260 4012 23980 4052
rect 24020 4012 24029 4052
rect 0 3968 80 3988
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 8227 3928 8236 3968
rect 8276 3928 21292 3968
rect 21332 3928 21341 3968
rect 22147 3928 22156 3968
rect 22196 3928 23212 3968
rect 23252 3928 25036 3968
rect 25076 3928 25085 3968
rect 28387 3928 28396 3968
rect 28436 3928 29452 3968
rect 29492 3928 33676 3968
rect 33716 3928 33725 3968
rect 47500 3928 48940 3968
rect 48980 3928 48989 3968
rect 0 3908 80 3928
rect 2467 3844 2476 3884
rect 2516 3844 30892 3884
rect 30932 3844 30941 3884
rect 31171 3844 31180 3884
rect 31220 3844 34348 3884
rect 34388 3844 37036 3884
rect 37076 3844 37612 3884
rect 37652 3844 37661 3884
rect 47500 3800 47540 3928
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 14179 3760 14188 3800
rect 14228 3760 17260 3800
rect 17300 3760 17309 3800
rect 17443 3760 17452 3800
rect 17492 3760 18700 3800
rect 18740 3760 19276 3800
rect 19316 3760 19325 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 20323 3760 20332 3800
rect 20372 3760 22060 3800
rect 22100 3760 22828 3800
rect 22868 3760 22877 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 47299 3760 47308 3800
rect 47348 3760 47540 3800
rect 48460 3844 52396 3884
rect 52436 3844 52445 3884
rect 48460 3716 48500 3844
rect 63331 3800 63389 3801
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 52291 3760 52300 3800
rect 52340 3760 63340 3800
rect 63380 3760 63389 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 63331 3759 63389 3760
rect 1699 3676 1708 3716
rect 1748 3676 30988 3716
rect 31028 3676 31037 3716
rect 31084 3676 34156 3716
rect 34196 3676 34205 3716
rect 47107 3676 47116 3716
rect 47156 3676 48500 3716
rect 48643 3676 48652 3716
rect 48692 3676 49612 3716
rect 49652 3676 51820 3716
rect 51860 3676 54604 3716
rect 54644 3676 54653 3716
rect 57580 3676 57772 3716
rect 57812 3676 57821 3716
rect 31084 3632 31124 3676
rect 33955 3632 34013 3633
rect 37219 3632 37277 3633
rect 1411 3592 1420 3632
rect 1460 3592 31124 3632
rect 33870 3592 33964 3632
rect 34004 3592 34013 3632
rect 34819 3592 34828 3632
rect 34868 3592 35212 3632
rect 35252 3592 35261 3632
rect 37134 3592 37228 3632
rect 37268 3592 37277 3632
rect 39331 3592 39340 3632
rect 39380 3592 40300 3632
rect 40340 3592 44908 3632
rect 44948 3592 44957 3632
rect 46444 3592 47596 3632
rect 47636 3592 48748 3632
rect 48788 3592 48797 3632
rect 48940 3592 52204 3632
rect 52244 3592 54892 3632
rect 54932 3592 55180 3632
rect 55220 3592 55229 3632
rect 33955 3591 34013 3592
rect 37219 3591 37277 3592
rect 46444 3548 46484 3592
rect 48940 3548 48980 3592
rect 57580 3548 57620 3676
rect 46435 3508 46444 3548
rect 46484 3508 46493 3548
rect 46915 3508 46924 3548
rect 46964 3508 48980 3548
rect 49027 3508 49036 3548
rect 49076 3508 52108 3548
rect 52148 3508 52157 3548
rect 52387 3508 52396 3548
rect 52436 3508 54988 3548
rect 55028 3508 57620 3548
rect 7075 3424 7084 3464
rect 7124 3424 42700 3464
rect 42740 3424 42749 3464
rect 68803 3380 68861 3381
rect 44515 3340 44524 3380
rect 44564 3340 68812 3380
rect 68852 3340 68861 3380
rect 68803 3339 68861 3340
rect 1987 3256 1996 3296
rect 2036 3256 37996 3296
rect 38036 3256 38045 3296
rect 30883 3172 30892 3212
rect 30932 3172 34060 3212
rect 34100 3172 36748 3212
rect 36788 3172 37324 3212
rect 37364 3172 38092 3212
rect 38132 3172 38141 3212
rect 0 3128 80 3148
rect 0 3088 652 3128
rect 692 3088 701 3128
rect 17251 3088 17260 3128
rect 17300 3088 20524 3128
rect 20564 3088 20573 3128
rect 23395 3088 23404 3128
rect 23444 3088 32716 3128
rect 32756 3088 32765 3128
rect 34915 3088 34924 3128
rect 34964 3088 35212 3128
rect 35252 3088 35261 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 12931 3004 12940 3044
rect 12980 3004 17588 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 21283 3004 21292 3044
rect 21332 3004 32236 3044
rect 32276 3004 32285 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 33859 3004 33868 3044
rect 33908 3004 35020 3044
rect 35060 3004 38188 3044
rect 38228 3004 46348 3044
rect 46388 3004 46397 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 17548 2960 17588 3004
rect 13219 2920 13228 2960
rect 13268 2920 17356 2960
rect 17396 2920 17405 2960
rect 17539 2920 17548 2960
rect 17588 2920 19948 2960
rect 19988 2920 20716 2960
rect 20756 2920 20765 2960
rect 22051 2920 22060 2960
rect 22100 2920 22540 2960
rect 22580 2920 22589 2960
rect 32035 2920 32044 2960
rect 32084 2920 34636 2960
rect 34676 2920 35980 2960
rect 36020 2920 36029 2960
rect 39619 2920 39628 2960
rect 39668 2920 41260 2960
rect 41300 2920 41309 2960
rect 42403 2920 42412 2960
rect 42452 2920 52300 2960
rect 52340 2920 52349 2960
rect 32044 2876 32084 2920
rect 55747 2876 55805 2877
rect 4771 2836 4780 2876
rect 4820 2836 15052 2876
rect 15092 2836 18124 2876
rect 18164 2836 18173 2876
rect 27139 2836 27148 2876
rect 27188 2836 28628 2876
rect 31267 2836 31276 2876
rect 31316 2836 32084 2876
rect 37987 2836 37996 2876
rect 38036 2836 39244 2876
rect 39284 2836 39724 2876
rect 39764 2836 41356 2876
rect 41396 2836 41405 2876
rect 55662 2836 55756 2876
rect 55796 2836 55805 2876
rect 28588 2792 28628 2836
rect 55747 2835 55805 2836
rect 69283 2792 69341 2793
rect 28579 2752 28588 2792
rect 28628 2752 31180 2792
rect 31220 2752 34828 2792
rect 34868 2752 34877 2792
rect 35299 2752 35308 2792
rect 35348 2752 35788 2792
rect 35828 2752 35837 2792
rect 43075 2752 43084 2792
rect 43124 2752 45676 2792
rect 45716 2752 45725 2792
rect 47500 2752 47980 2792
rect 48020 2752 48652 2792
rect 48692 2752 50860 2792
rect 50900 2752 51244 2792
rect 51284 2752 69292 2792
rect 69332 2752 69341 2792
rect 47500 2708 47540 2752
rect 69283 2751 69341 2752
rect 6883 2668 6892 2708
rect 6932 2668 23404 2708
rect 23444 2668 23453 2708
rect 23500 2668 25132 2708
rect 25172 2668 26860 2708
rect 26900 2668 28396 2708
rect 28436 2668 28445 2708
rect 32611 2668 32620 2708
rect 32660 2668 33196 2708
rect 33236 2668 36172 2708
rect 36212 2668 36844 2708
rect 36884 2668 36893 2708
rect 40867 2668 40876 2708
rect 40916 2668 42796 2708
rect 42836 2668 43276 2708
rect 43316 2668 43325 2708
rect 46051 2668 46060 2708
rect 46100 2668 47540 2708
rect 53827 2668 53836 2708
rect 53876 2668 54028 2708
rect 54068 2668 56620 2708
rect 56660 2668 80716 2708
rect 80756 2668 80765 2708
rect 7843 2624 7901 2625
rect 23500 2624 23540 2668
rect 7843 2584 7852 2624
rect 7892 2584 17260 2624
rect 17300 2584 17309 2624
rect 23107 2584 23116 2624
rect 23156 2584 23540 2624
rect 23875 2584 23884 2624
rect 23924 2584 27244 2624
rect 27284 2584 28916 2624
rect 28963 2584 28972 2624
rect 29012 2584 30028 2624
rect 30068 2584 37036 2624
rect 37076 2584 71980 2624
rect 72020 2584 72029 2624
rect 7843 2583 7901 2584
rect 28876 2540 28916 2584
rect 25507 2500 25516 2540
rect 25556 2500 28396 2540
rect 28436 2500 28445 2540
rect 28876 2500 31468 2540
rect 31508 2500 31517 2540
rect 38083 2500 38092 2540
rect 38132 2500 39340 2540
rect 39380 2500 40876 2540
rect 40916 2500 40925 2540
rect 44131 2500 44140 2540
rect 44180 2500 45004 2540
rect 45044 2500 45292 2540
rect 45332 2500 46924 2540
rect 46964 2500 47116 2540
rect 47156 2500 49516 2540
rect 49556 2500 49996 2540
rect 50036 2500 52108 2540
rect 52148 2500 53164 2540
rect 53204 2500 53213 2540
rect 23491 2416 23500 2456
rect 23540 2416 25420 2456
rect 25460 2416 26476 2456
rect 26516 2416 26525 2456
rect 28099 2416 28108 2456
rect 28148 2416 29164 2456
rect 29204 2416 30700 2456
rect 30740 2416 30749 2456
rect 28108 2372 28148 2416
rect 23203 2332 23212 2372
rect 23252 2332 24460 2372
rect 24500 2332 26380 2372
rect 26420 2332 28148 2372
rect 30115 2332 30124 2372
rect 30164 2332 35116 2372
rect 35156 2332 35165 2372
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 36835 2248 36844 2288
rect 36884 2248 38092 2288
rect 38132 2248 38141 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 0 2228 80 2248
rect 28387 2164 28396 2204
rect 28436 2164 39820 2204
rect 39860 2164 39869 2204
rect 40579 2164 40588 2204
rect 40628 2164 41644 2204
rect 41684 2164 42124 2204
rect 42164 2164 42700 2204
rect 42740 2164 42749 2204
rect 29731 2080 29740 2120
rect 29780 2080 31660 2120
rect 31700 2080 34444 2120
rect 34484 2080 34493 2120
rect 45187 2080 45196 2120
rect 45236 2080 54700 2120
rect 54740 2080 55756 2120
rect 55796 2080 55805 2120
rect 69091 2036 69149 2037
rect 22531 1996 22540 2036
rect 22580 1996 23404 2036
rect 23444 1996 25036 2036
rect 25076 1996 25085 2036
rect 31555 1996 31564 2036
rect 31604 1996 34828 2036
rect 34868 1996 35500 2036
rect 35540 1996 35692 2036
rect 35732 1996 35741 2036
rect 38947 1996 38956 2036
rect 38996 1996 40204 2036
rect 40244 1996 41740 2036
rect 41780 1996 43276 2036
rect 43316 1996 44428 2036
rect 44468 1996 69100 2036
rect 69140 1996 69149 2036
rect 69091 1995 69149 1996
rect 69187 1952 69245 1953
rect 18115 1912 18124 1952
rect 18164 1912 19756 1952
rect 19796 1912 21388 1952
rect 21428 1912 21437 1952
rect 21763 1912 21772 1952
rect 21812 1912 22156 1952
rect 22196 1912 23116 1952
rect 23156 1912 23165 1952
rect 25315 1912 25324 1952
rect 25364 1912 28972 1952
rect 29012 1912 29021 1952
rect 31459 1912 31468 1952
rect 31508 1912 33388 1952
rect 33428 1912 34060 1952
rect 34100 1912 35980 1952
rect 36020 1912 69196 1952
rect 69236 1912 69245 1952
rect 78979 1912 78988 1952
rect 79028 1912 79948 1952
rect 79988 1912 79997 1952
rect 69187 1911 69245 1912
rect 19939 1828 19948 1868
rect 19988 1828 27244 1868
rect 27284 1828 30124 1868
rect 30164 1828 30173 1868
rect 35395 1828 35404 1868
rect 35444 1828 37228 1868
rect 37268 1828 37277 1868
rect 50275 1828 50284 1868
rect 50324 1828 52492 1868
rect 52532 1828 52541 1868
rect 52771 1828 52780 1868
rect 52820 1828 55084 1868
rect 55124 1828 55133 1868
rect 41923 1744 41932 1784
rect 41972 1744 44524 1784
rect 44564 1744 44573 1784
rect 78595 1576 78604 1616
rect 78644 1576 80236 1616
rect 80276 1576 80524 1616
rect 80564 1576 80573 1616
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 18691 1492 18700 1532
rect 18740 1492 20044 1532
rect 20084 1492 20428 1532
rect 20468 1492 20477 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 39811 1492 39820 1532
rect 39860 1492 42988 1532
rect 43028 1492 43037 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 79939 1492 79948 1532
rect 79988 1492 81868 1532
rect 81908 1492 81917 1532
rect 36547 1408 36556 1448
rect 36596 1408 47212 1448
rect 47252 1408 49996 1448
rect 50036 1408 50045 1448
rect 79171 1408 79180 1448
rect 79220 1408 82060 1448
rect 82100 1408 82109 1448
rect 28675 1324 28684 1364
rect 28724 1324 29836 1364
rect 29876 1324 32716 1364
rect 32756 1324 35308 1364
rect 35348 1324 35357 1364
rect 40003 1324 40012 1364
rect 40052 1324 41548 1364
rect 41588 1324 42892 1364
rect 42932 1324 42941 1364
rect 45091 1324 45100 1364
rect 45140 1324 47308 1364
rect 47348 1324 47357 1364
rect 47587 1324 47596 1364
rect 47636 1324 49900 1364
rect 49940 1324 49949 1364
rect 37891 1240 37900 1280
rect 37940 1240 39916 1280
rect 39956 1240 39965 1280
rect 46924 1240 49612 1280
rect 49652 1240 49661 1280
rect 36067 1156 36076 1196
rect 36116 1156 38284 1196
rect 38324 1156 39628 1196
rect 39668 1156 39677 1196
rect 46924 1112 46964 1240
rect 47395 1156 47404 1196
rect 47444 1156 49900 1196
rect 49940 1156 52492 1196
rect 52532 1156 52684 1196
rect 52724 1156 52733 1196
rect 23875 1072 23884 1112
rect 23924 1072 25324 1112
rect 25364 1072 25373 1112
rect 35779 1072 35788 1112
rect 35828 1072 37900 1112
rect 37940 1072 37949 1112
rect 42403 1072 42412 1112
rect 42452 1072 44428 1112
rect 44468 1072 45964 1112
rect 46004 1072 46924 1112
rect 46964 1072 46973 1112
rect 88684 1028 89057 1041
rect 39523 988 39532 1028
rect 39572 988 44716 1028
rect 44756 988 47308 1028
rect 47348 988 47500 1028
rect 47540 988 47549 1028
rect 79843 988 79852 1028
rect 79892 988 80620 1028
rect 80660 988 81964 1028
rect 82004 1001 89057 1028
rect 89097 1001 89106 1041
rect 82004 988 88724 1001
rect 82051 904 82060 944
rect 82100 904 94233 944
rect 94273 904 94282 944
rect 38371 820 38380 860
rect 38420 820 89260 860
rect 89300 820 89309 860
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 81859 736 81868 776
rect 81908 736 90777 776
rect 90817 736 90826 776
rect 30787 652 30796 692
rect 30836 652 90988 692
rect 91028 652 91037 692
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 4780 35848 4820 35888
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 20812 34504 20852 34544
rect 50188 34504 50228 34544
rect 42124 34420 42164 34460
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 50188 33748 50228 33788
rect 22924 33412 22964 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 17452 33076 17492 33116
rect 68812 33076 68852 33116
rect 17452 32656 17492 32696
rect 69100 32656 69140 32696
rect 61996 32572 62036 32612
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 4972 32236 5012 32276
rect 66220 32236 66260 32276
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 69292 31648 69332 31688
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 69196 31060 69236 31100
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 97321 30472 97361 30512
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 7852 30052 7892 30092
rect 22924 30052 22964 30092
rect 3532 29464 3572 29504
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 4204 26188 4244 26228
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 4972 24424 5012 24464
rect 3532 24340 3572 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 4204 23248 4244 23288
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 4204 21736 4244 21776
rect 6412 21484 6452 21524
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 76972 17200 77012 17240
rect 82924 17116 82964 17156
rect 91084 17116 91124 17156
rect 91084 16780 91124 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 6412 14428 6452 14468
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 4780 13168 4820 13208
rect 6604 13000 6644 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 99940 11461 99980 11501
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 1804 11152 1844 11192
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 99921 8968 99961 9008
rect 83500 8800 83540 8840
rect 99940 8773 99980 8813
rect 1708 8464 1748 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 99940 6253 99980 6293
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 26860 5860 26900 5900
rect 72748 5776 72788 5816
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 6604 5188 6644 5228
rect 6412 5104 6452 5144
rect 73036 5020 73076 5060
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 63340 3760 63380 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 33964 3592 34004 3632
rect 37228 3592 37268 3632
rect 68812 3340 68852 3380
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 55756 2836 55796 2876
rect 69292 2752 69332 2792
rect 7852 2584 7892 2624
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 69100 1996 69140 2036
rect 69196 1912 69236 1952
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 4780 35888 4820 35897
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3532 29504 3572 29513
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3532 24380 3572 29464
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3532 24331 3572 24340
rect 4204 26228 4244 26237
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 4204 23288 4244 26188
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4204 21776 4244 23248
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 4204 21727 4244 21736
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4780 13208 4820 35848
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 20812 34544 20852 34555
rect 20812 34469 20852 34504
rect 50188 34544 50228 34553
rect 20811 34460 20853 34469
rect 20811 34420 20812 34460
rect 20852 34420 20853 34460
rect 20811 34411 20853 34420
rect 42123 34460 42165 34469
rect 42123 34420 42124 34460
rect 42164 34420 42165 34460
rect 42123 34411 42165 34420
rect 42124 34326 42164 34411
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 50188 33788 50228 34504
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 50188 33739 50228 33748
rect 22924 33452 22964 33461
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 17452 33116 17492 33125
rect 17452 32696 17492 33076
rect 17452 32647 17492 32656
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 4972 32276 5012 32285
rect 4972 24464 5012 32236
rect 6411 30512 6453 30521
rect 6411 30472 6412 30512
rect 6452 30472 6453 30512
rect 6411 30463 6453 30472
rect 4972 24415 5012 24424
rect 6412 21524 6452 30463
rect 6412 21475 6452 21484
rect 7852 30092 7892 30101
rect 4780 13159 4820 13168
rect 6412 14468 6452 14477
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 1804 11192 1844 11201
rect 1708 8504 1748 8513
rect 1708 5657 1748 8464
rect 1804 5741 1844 11152
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 1803 5732 1845 5741
rect 1803 5692 1804 5732
rect 1844 5692 1845 5732
rect 1803 5683 1845 5692
rect 1707 5648 1749 5657
rect 1707 5608 1708 5648
rect 1748 5608 1749 5648
rect 1707 5599 1749 5608
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 6412 5144 6452 14428
rect 6604 13040 6644 13049
rect 6604 5228 6644 13000
rect 6604 5179 6644 5188
rect 6412 5095 6452 5104
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 7852 2624 7892 30052
rect 22924 30092 22964 33412
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 68812 33116 68852 33125
rect 61996 32612 62036 32621
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 22924 30043 22964 30052
rect 61996 28757 62036 32572
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 66220 32276 66260 32285
rect 61995 28748 62037 28757
rect 61995 28708 61996 28748
rect 62036 28708 62037 28748
rect 61995 28699 62037 28708
rect 66220 28589 66260 32236
rect 66219 28580 66261 28589
rect 66219 28540 66220 28580
rect 66260 28540 66261 28580
rect 66219 28531 66261 28540
rect 26859 6068 26901 6077
rect 26859 6028 26860 6068
rect 26900 6028 26901 6068
rect 26859 6019 26901 6028
rect 26860 5900 26900 6019
rect 26860 5851 26900 5860
rect 55755 5060 55797 5069
rect 55755 5020 55756 5060
rect 55796 5020 55797 5060
rect 55755 5011 55797 5020
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 33964 3632 34004 3641
rect 33964 3473 34004 3592
rect 37227 3632 37269 3641
rect 37227 3592 37228 3632
rect 37268 3592 37269 3632
rect 37227 3583 37269 3592
rect 37228 3498 37268 3583
rect 33963 3464 34005 3473
rect 33963 3424 33964 3464
rect 34004 3424 34005 3464
rect 33963 3415 34005 3424
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 55756 2876 55796 5011
rect 63339 4472 63381 4481
rect 63339 4432 63340 4472
rect 63380 4432 63381 4472
rect 63339 4423 63381 4432
rect 63340 3800 63380 4423
rect 63340 3751 63380 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 68812 3380 68852 33076
rect 68812 3331 68852 3340
rect 69100 32696 69140 32705
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 55756 2827 55796 2836
rect 7852 2575 7892 2584
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 69100 2036 69140 32656
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 69292 31688 69332 31697
rect 69100 1987 69140 1996
rect 69196 31100 69236 31109
rect 69196 1952 69236 31060
rect 69292 2792 69332 31648
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 97320 30512 97362 30521
rect 97320 30472 97321 30512
rect 97361 30472 97362 30512
rect 97320 30463 97362 30472
rect 97321 30378 97361 30463
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 76972 17240 77012 17249
rect 73035 8924 73077 8933
rect 73035 8884 73036 8924
rect 73076 8884 73077 8924
rect 73035 8875 73077 8884
rect 72747 6068 72789 6077
rect 72747 6028 72748 6068
rect 72788 6028 72789 6068
rect 72747 6019 72789 6028
rect 72748 5816 72788 6019
rect 72748 5767 72788 5776
rect 73036 5060 73076 8875
rect 76972 5657 77012 17200
rect 82924 17156 82964 17165
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 82924 5741 82964 17116
rect 91084 17156 91124 17165
rect 91084 16820 91124 17116
rect 91084 16771 91124 16780
rect 99940 11501 99980 11510
rect 99940 11201 99980 11461
rect 95691 11192 95733 11201
rect 95691 11152 95692 11192
rect 95732 11152 95733 11192
rect 95691 11143 95733 11152
rect 99939 11192 99981 11201
rect 99939 11152 99940 11192
rect 99980 11152 99981 11192
rect 99939 11143 99981 11152
rect 83499 8840 83541 8849
rect 83499 8800 83500 8840
rect 83540 8800 83541 8840
rect 83499 8791 83541 8800
rect 83500 8706 83540 8791
rect 93579 6068 93621 6077
rect 93579 6028 93580 6068
rect 93620 6028 93621 6068
rect 93579 6019 93621 6028
rect 82923 5732 82965 5741
rect 82923 5692 82924 5732
rect 82964 5692 82965 5732
rect 82923 5683 82965 5692
rect 76971 5648 77013 5657
rect 76971 5608 76972 5648
rect 77012 5608 77013 5648
rect 76971 5599 77013 5608
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 73036 5011 73076 5020
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 93580 3473 93620 6019
rect 95692 3557 95732 11143
rect 99920 9008 99962 9017
rect 99920 8968 99921 9008
rect 99961 8968 99962 9008
rect 99920 8959 99962 8968
rect 99921 8874 99961 8959
rect 99940 8813 99980 8822
rect 99940 8765 99980 8773
rect 99928 8756 99980 8765
rect 99928 8716 99929 8756
rect 99969 8716 99980 8756
rect 99928 8707 99970 8716
rect 99929 8689 99969 8707
rect 99940 6293 99980 6302
rect 99940 6077 99980 6253
rect 99939 6068 99981 6077
rect 99939 6028 99940 6068
rect 99980 6028 99981 6068
rect 99939 6019 99981 6028
rect 95691 3548 95733 3557
rect 95691 3508 95692 3548
rect 95732 3508 95733 3548
rect 95691 3499 95733 3508
rect 93579 3464 93621 3473
rect 93579 3424 93580 3464
rect 93620 3424 93621 3464
rect 93579 3415 93621 3424
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 69292 2743 69332 2752
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 69196 1903 69236 1912
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 20812 34420 20852 34460
rect 42124 34420 42164 34460
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 6412 30472 6452 30512
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 1804 5692 1844 5732
rect 1708 5608 1748 5648
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 61996 28708 62036 28748
rect 66220 28540 66260 28580
rect 26860 6028 26900 6068
rect 55756 5020 55796 5060
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 37228 3592 37268 3632
rect 33964 3424 34004 3464
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63340 4432 63380 4472
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 97321 30472 97361 30512
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 73036 8884 73076 8924
rect 72748 6028 72788 6068
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 95692 11152 95732 11192
rect 99940 11152 99980 11192
rect 83500 8800 83540 8840
rect 93580 6028 93620 6068
rect 82924 5692 82964 5732
rect 76972 5608 77012 5648
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 99921 8968 99961 9008
rect 99929 8716 99969 8756
rect 99940 6028 99980 6068
rect 95692 3508 95732 3548
rect 93580 3424 93620 3464
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal5 >>
rect 4343 38576 4390 38618
rect 4514 38576 4558 38618
rect 4682 38576 4729 38618
rect 4343 38536 4352 38576
rect 4514 38536 4516 38576
rect 4556 38536 4558 38576
rect 4720 38536 4729 38576
rect 4343 38494 4390 38536
rect 4514 38494 4558 38536
rect 4682 38494 4729 38536
rect 19463 38576 19510 38618
rect 19634 38576 19678 38618
rect 19802 38576 19849 38618
rect 19463 38536 19472 38576
rect 19634 38536 19636 38576
rect 19676 38536 19678 38576
rect 19840 38536 19849 38576
rect 19463 38494 19510 38536
rect 19634 38494 19678 38536
rect 19802 38494 19849 38536
rect 34583 38576 34630 38618
rect 34754 38576 34798 38618
rect 34922 38576 34969 38618
rect 34583 38536 34592 38576
rect 34754 38536 34756 38576
rect 34796 38536 34798 38576
rect 34960 38536 34969 38576
rect 34583 38494 34630 38536
rect 34754 38494 34798 38536
rect 34922 38494 34969 38536
rect 49703 38576 49750 38618
rect 49874 38576 49918 38618
rect 50042 38576 50089 38618
rect 49703 38536 49712 38576
rect 49874 38536 49876 38576
rect 49916 38536 49918 38576
rect 50080 38536 50089 38576
rect 49703 38494 49750 38536
rect 49874 38494 49918 38536
rect 50042 38494 50089 38536
rect 64823 38576 64870 38618
rect 64994 38576 65038 38618
rect 65162 38576 65209 38618
rect 64823 38536 64832 38576
rect 64994 38536 64996 38576
rect 65036 38536 65038 38576
rect 65200 38536 65209 38576
rect 64823 38494 64870 38536
rect 64994 38494 65038 38536
rect 65162 38494 65209 38536
rect 79943 38576 79990 38618
rect 80114 38576 80158 38618
rect 80282 38576 80329 38618
rect 79943 38536 79952 38576
rect 80114 38536 80116 38576
rect 80156 38536 80158 38576
rect 80320 38536 80329 38576
rect 79943 38494 79990 38536
rect 80114 38494 80158 38536
rect 80282 38494 80329 38536
rect 3103 37820 3150 37862
rect 3274 37820 3318 37862
rect 3442 37820 3489 37862
rect 3103 37780 3112 37820
rect 3274 37780 3276 37820
rect 3316 37780 3318 37820
rect 3480 37780 3489 37820
rect 3103 37738 3150 37780
rect 3274 37738 3318 37780
rect 3442 37738 3489 37780
rect 18223 37820 18270 37862
rect 18394 37820 18438 37862
rect 18562 37820 18609 37862
rect 18223 37780 18232 37820
rect 18394 37780 18396 37820
rect 18436 37780 18438 37820
rect 18600 37780 18609 37820
rect 18223 37738 18270 37780
rect 18394 37738 18438 37780
rect 18562 37738 18609 37780
rect 33343 37820 33390 37862
rect 33514 37820 33558 37862
rect 33682 37820 33729 37862
rect 33343 37780 33352 37820
rect 33514 37780 33516 37820
rect 33556 37780 33558 37820
rect 33720 37780 33729 37820
rect 33343 37738 33390 37780
rect 33514 37738 33558 37780
rect 33682 37738 33729 37780
rect 48463 37820 48510 37862
rect 48634 37820 48678 37862
rect 48802 37820 48849 37862
rect 48463 37780 48472 37820
rect 48634 37780 48636 37820
rect 48676 37780 48678 37820
rect 48840 37780 48849 37820
rect 48463 37738 48510 37780
rect 48634 37738 48678 37780
rect 48802 37738 48849 37780
rect 63583 37820 63630 37862
rect 63754 37820 63798 37862
rect 63922 37820 63969 37862
rect 63583 37780 63592 37820
rect 63754 37780 63756 37820
rect 63796 37780 63798 37820
rect 63960 37780 63969 37820
rect 63583 37738 63630 37780
rect 63754 37738 63798 37780
rect 63922 37738 63969 37780
rect 78703 37820 78750 37862
rect 78874 37820 78918 37862
rect 79042 37820 79089 37862
rect 78703 37780 78712 37820
rect 78874 37780 78876 37820
rect 78916 37780 78918 37820
rect 79080 37780 79089 37820
rect 78703 37738 78750 37780
rect 78874 37738 78918 37780
rect 79042 37738 79089 37780
rect 4343 37064 4390 37106
rect 4514 37064 4558 37106
rect 4682 37064 4729 37106
rect 4343 37024 4352 37064
rect 4514 37024 4516 37064
rect 4556 37024 4558 37064
rect 4720 37024 4729 37064
rect 4343 36982 4390 37024
rect 4514 36982 4558 37024
rect 4682 36982 4729 37024
rect 19463 37064 19510 37106
rect 19634 37064 19678 37106
rect 19802 37064 19849 37106
rect 19463 37024 19472 37064
rect 19634 37024 19636 37064
rect 19676 37024 19678 37064
rect 19840 37024 19849 37064
rect 19463 36982 19510 37024
rect 19634 36982 19678 37024
rect 19802 36982 19849 37024
rect 34583 37064 34630 37106
rect 34754 37064 34798 37106
rect 34922 37064 34969 37106
rect 34583 37024 34592 37064
rect 34754 37024 34756 37064
rect 34796 37024 34798 37064
rect 34960 37024 34969 37064
rect 34583 36982 34630 37024
rect 34754 36982 34798 37024
rect 34922 36982 34969 37024
rect 49703 37064 49750 37106
rect 49874 37064 49918 37106
rect 50042 37064 50089 37106
rect 49703 37024 49712 37064
rect 49874 37024 49876 37064
rect 49916 37024 49918 37064
rect 50080 37024 50089 37064
rect 49703 36982 49750 37024
rect 49874 36982 49918 37024
rect 50042 36982 50089 37024
rect 64823 37064 64870 37106
rect 64994 37064 65038 37106
rect 65162 37064 65209 37106
rect 64823 37024 64832 37064
rect 64994 37024 64996 37064
rect 65036 37024 65038 37064
rect 65200 37024 65209 37064
rect 64823 36982 64870 37024
rect 64994 36982 65038 37024
rect 65162 36982 65209 37024
rect 79943 37064 79990 37106
rect 80114 37064 80158 37106
rect 80282 37064 80329 37106
rect 79943 37024 79952 37064
rect 80114 37024 80116 37064
rect 80156 37024 80158 37064
rect 80320 37024 80329 37064
rect 79943 36982 79990 37024
rect 80114 36982 80158 37024
rect 80282 36982 80329 37024
rect 3103 36308 3150 36350
rect 3274 36308 3318 36350
rect 3442 36308 3489 36350
rect 3103 36268 3112 36308
rect 3274 36268 3276 36308
rect 3316 36268 3318 36308
rect 3480 36268 3489 36308
rect 3103 36226 3150 36268
rect 3274 36226 3318 36268
rect 3442 36226 3489 36268
rect 18223 36308 18270 36350
rect 18394 36308 18438 36350
rect 18562 36308 18609 36350
rect 18223 36268 18232 36308
rect 18394 36268 18396 36308
rect 18436 36268 18438 36308
rect 18600 36268 18609 36308
rect 18223 36226 18270 36268
rect 18394 36226 18438 36268
rect 18562 36226 18609 36268
rect 33343 36308 33390 36350
rect 33514 36308 33558 36350
rect 33682 36308 33729 36350
rect 33343 36268 33352 36308
rect 33514 36268 33516 36308
rect 33556 36268 33558 36308
rect 33720 36268 33729 36308
rect 33343 36226 33390 36268
rect 33514 36226 33558 36268
rect 33682 36226 33729 36268
rect 48463 36308 48510 36350
rect 48634 36308 48678 36350
rect 48802 36308 48849 36350
rect 48463 36268 48472 36308
rect 48634 36268 48636 36308
rect 48676 36268 48678 36308
rect 48840 36268 48849 36308
rect 48463 36226 48510 36268
rect 48634 36226 48678 36268
rect 48802 36226 48849 36268
rect 63583 36308 63630 36350
rect 63754 36308 63798 36350
rect 63922 36308 63969 36350
rect 63583 36268 63592 36308
rect 63754 36268 63756 36308
rect 63796 36268 63798 36308
rect 63960 36268 63969 36308
rect 63583 36226 63630 36268
rect 63754 36226 63798 36268
rect 63922 36226 63969 36268
rect 78703 36308 78750 36350
rect 78874 36308 78918 36350
rect 79042 36308 79089 36350
rect 78703 36268 78712 36308
rect 78874 36268 78876 36308
rect 78916 36268 78918 36308
rect 79080 36268 79089 36308
rect 78703 36226 78750 36268
rect 78874 36226 78918 36268
rect 79042 36226 79089 36268
rect 4343 35552 4390 35594
rect 4514 35552 4558 35594
rect 4682 35552 4729 35594
rect 4343 35512 4352 35552
rect 4514 35512 4516 35552
rect 4556 35512 4558 35552
rect 4720 35512 4729 35552
rect 4343 35470 4390 35512
rect 4514 35470 4558 35512
rect 4682 35470 4729 35512
rect 19463 35552 19510 35594
rect 19634 35552 19678 35594
rect 19802 35552 19849 35594
rect 19463 35512 19472 35552
rect 19634 35512 19636 35552
rect 19676 35512 19678 35552
rect 19840 35512 19849 35552
rect 19463 35470 19510 35512
rect 19634 35470 19678 35512
rect 19802 35470 19849 35512
rect 34583 35552 34630 35594
rect 34754 35552 34798 35594
rect 34922 35552 34969 35594
rect 34583 35512 34592 35552
rect 34754 35512 34756 35552
rect 34796 35512 34798 35552
rect 34960 35512 34969 35552
rect 34583 35470 34630 35512
rect 34754 35470 34798 35512
rect 34922 35470 34969 35512
rect 49703 35552 49750 35594
rect 49874 35552 49918 35594
rect 50042 35552 50089 35594
rect 49703 35512 49712 35552
rect 49874 35512 49876 35552
rect 49916 35512 49918 35552
rect 50080 35512 50089 35552
rect 49703 35470 49750 35512
rect 49874 35470 49918 35512
rect 50042 35470 50089 35512
rect 64823 35552 64870 35594
rect 64994 35552 65038 35594
rect 65162 35552 65209 35594
rect 64823 35512 64832 35552
rect 64994 35512 64996 35552
rect 65036 35512 65038 35552
rect 65200 35512 65209 35552
rect 64823 35470 64870 35512
rect 64994 35470 65038 35512
rect 65162 35470 65209 35512
rect 79943 35552 79990 35594
rect 80114 35552 80158 35594
rect 80282 35552 80329 35594
rect 79943 35512 79952 35552
rect 80114 35512 80116 35552
rect 80156 35512 80158 35552
rect 80320 35512 80329 35552
rect 79943 35470 79990 35512
rect 80114 35470 80158 35512
rect 80282 35470 80329 35512
rect 3103 34796 3150 34838
rect 3274 34796 3318 34838
rect 3442 34796 3489 34838
rect 3103 34756 3112 34796
rect 3274 34756 3276 34796
rect 3316 34756 3318 34796
rect 3480 34756 3489 34796
rect 3103 34714 3150 34756
rect 3274 34714 3318 34756
rect 3442 34714 3489 34756
rect 18223 34796 18270 34838
rect 18394 34796 18438 34838
rect 18562 34796 18609 34838
rect 18223 34756 18232 34796
rect 18394 34756 18396 34796
rect 18436 34756 18438 34796
rect 18600 34756 18609 34796
rect 18223 34714 18270 34756
rect 18394 34714 18438 34756
rect 18562 34714 18609 34756
rect 33343 34796 33390 34838
rect 33514 34796 33558 34838
rect 33682 34796 33729 34838
rect 33343 34756 33352 34796
rect 33514 34756 33516 34796
rect 33556 34756 33558 34796
rect 33720 34756 33729 34796
rect 33343 34714 33390 34756
rect 33514 34714 33558 34756
rect 33682 34714 33729 34756
rect 48463 34796 48510 34838
rect 48634 34796 48678 34838
rect 48802 34796 48849 34838
rect 48463 34756 48472 34796
rect 48634 34756 48636 34796
rect 48676 34756 48678 34796
rect 48840 34756 48849 34796
rect 48463 34714 48510 34756
rect 48634 34714 48678 34756
rect 48802 34714 48849 34756
rect 63583 34796 63630 34838
rect 63754 34796 63798 34838
rect 63922 34796 63969 34838
rect 63583 34756 63592 34796
rect 63754 34756 63756 34796
rect 63796 34756 63798 34796
rect 63960 34756 63969 34796
rect 63583 34714 63630 34756
rect 63754 34714 63798 34756
rect 63922 34714 63969 34756
rect 78703 34796 78750 34838
rect 78874 34796 78918 34838
rect 79042 34796 79089 34838
rect 78703 34756 78712 34796
rect 78874 34756 78876 34796
rect 78916 34756 78918 34796
rect 79080 34756 79089 34796
rect 78703 34714 78750 34756
rect 78874 34714 78918 34756
rect 79042 34714 79089 34756
rect 20803 34420 20812 34460
rect 20852 34420 42124 34460
rect 42164 34420 42173 34460
rect 4343 34040 4390 34082
rect 4514 34040 4558 34082
rect 4682 34040 4729 34082
rect 4343 34000 4352 34040
rect 4514 34000 4516 34040
rect 4556 34000 4558 34040
rect 4720 34000 4729 34040
rect 4343 33958 4390 34000
rect 4514 33958 4558 34000
rect 4682 33958 4729 34000
rect 19463 34040 19510 34082
rect 19634 34040 19678 34082
rect 19802 34040 19849 34082
rect 19463 34000 19472 34040
rect 19634 34000 19636 34040
rect 19676 34000 19678 34040
rect 19840 34000 19849 34040
rect 19463 33958 19510 34000
rect 19634 33958 19678 34000
rect 19802 33958 19849 34000
rect 34583 34040 34630 34082
rect 34754 34040 34798 34082
rect 34922 34040 34969 34082
rect 34583 34000 34592 34040
rect 34754 34000 34756 34040
rect 34796 34000 34798 34040
rect 34960 34000 34969 34040
rect 34583 33958 34630 34000
rect 34754 33958 34798 34000
rect 34922 33958 34969 34000
rect 49703 34040 49750 34082
rect 49874 34040 49918 34082
rect 50042 34040 50089 34082
rect 49703 34000 49712 34040
rect 49874 34000 49876 34040
rect 49916 34000 49918 34040
rect 50080 34000 50089 34040
rect 49703 33958 49750 34000
rect 49874 33958 49918 34000
rect 50042 33958 50089 34000
rect 64823 34040 64870 34082
rect 64994 34040 65038 34082
rect 65162 34040 65209 34082
rect 64823 34000 64832 34040
rect 64994 34000 64996 34040
rect 65036 34000 65038 34040
rect 65200 34000 65209 34040
rect 64823 33958 64870 34000
rect 64994 33958 65038 34000
rect 65162 33958 65209 34000
rect 79943 34040 79990 34082
rect 80114 34040 80158 34082
rect 80282 34040 80329 34082
rect 79943 34000 79952 34040
rect 80114 34000 80116 34040
rect 80156 34000 80158 34040
rect 80320 34000 80329 34040
rect 79943 33958 79990 34000
rect 80114 33958 80158 34000
rect 80282 33958 80329 34000
rect 93796 33822 94236 33896
rect 93796 33698 93870 33822
rect 93994 33698 94038 33822
rect 94162 33698 94236 33822
rect 93796 33654 94236 33698
rect 93796 33530 93870 33654
rect 93994 33530 94038 33654
rect 94162 33530 94236 33654
rect 93796 33456 94236 33530
rect 3103 33284 3150 33326
rect 3274 33284 3318 33326
rect 3442 33284 3489 33326
rect 3103 33244 3112 33284
rect 3274 33244 3276 33284
rect 3316 33244 3318 33284
rect 3480 33244 3489 33284
rect 3103 33202 3150 33244
rect 3274 33202 3318 33244
rect 3442 33202 3489 33244
rect 18223 33284 18270 33326
rect 18394 33284 18438 33326
rect 18562 33284 18609 33326
rect 18223 33244 18232 33284
rect 18394 33244 18396 33284
rect 18436 33244 18438 33284
rect 18600 33244 18609 33284
rect 18223 33202 18270 33244
rect 18394 33202 18438 33244
rect 18562 33202 18609 33244
rect 33343 33284 33390 33326
rect 33514 33284 33558 33326
rect 33682 33284 33729 33326
rect 33343 33244 33352 33284
rect 33514 33244 33516 33284
rect 33556 33244 33558 33284
rect 33720 33244 33729 33284
rect 33343 33202 33390 33244
rect 33514 33202 33558 33244
rect 33682 33202 33729 33244
rect 48463 33284 48510 33326
rect 48634 33284 48678 33326
rect 48802 33284 48849 33326
rect 48463 33244 48472 33284
rect 48634 33244 48636 33284
rect 48676 33244 48678 33284
rect 48840 33244 48849 33284
rect 48463 33202 48510 33244
rect 48634 33202 48678 33244
rect 48802 33202 48849 33244
rect 63583 33284 63630 33326
rect 63754 33284 63798 33326
rect 63922 33284 63969 33326
rect 63583 33244 63592 33284
rect 63754 33244 63756 33284
rect 63796 33244 63798 33284
rect 63960 33244 63969 33284
rect 63583 33202 63630 33244
rect 63754 33202 63798 33244
rect 63922 33202 63969 33244
rect 78703 33284 78750 33326
rect 78874 33284 78918 33326
rect 79042 33284 79089 33326
rect 78703 33244 78712 33284
rect 78874 33244 78876 33284
rect 78916 33244 78918 33284
rect 79080 33244 79089 33284
rect 78703 33202 78750 33244
rect 78874 33202 78918 33244
rect 79042 33202 79089 33244
rect 4343 32528 4390 32570
rect 4514 32528 4558 32570
rect 4682 32528 4729 32570
rect 4343 32488 4352 32528
rect 4514 32488 4516 32528
rect 4556 32488 4558 32528
rect 4720 32488 4729 32528
rect 4343 32446 4390 32488
rect 4514 32446 4558 32488
rect 4682 32446 4729 32488
rect 19463 32528 19510 32570
rect 19634 32528 19678 32570
rect 19802 32528 19849 32570
rect 19463 32488 19472 32528
rect 19634 32488 19636 32528
rect 19676 32488 19678 32528
rect 19840 32488 19849 32528
rect 19463 32446 19510 32488
rect 19634 32446 19678 32488
rect 19802 32446 19849 32488
rect 34583 32528 34630 32570
rect 34754 32528 34798 32570
rect 34922 32528 34969 32570
rect 34583 32488 34592 32528
rect 34754 32488 34756 32528
rect 34796 32488 34798 32528
rect 34960 32488 34969 32528
rect 34583 32446 34630 32488
rect 34754 32446 34798 32488
rect 34922 32446 34969 32488
rect 49703 32528 49750 32570
rect 49874 32528 49918 32570
rect 50042 32528 50089 32570
rect 49703 32488 49712 32528
rect 49874 32488 49876 32528
rect 49916 32488 49918 32528
rect 50080 32488 50089 32528
rect 49703 32446 49750 32488
rect 49874 32446 49918 32488
rect 50042 32446 50089 32488
rect 64823 32528 64870 32570
rect 64994 32528 65038 32570
rect 65162 32528 65209 32570
rect 64823 32488 64832 32528
rect 64994 32488 64996 32528
rect 65036 32488 65038 32528
rect 65200 32488 65209 32528
rect 64823 32446 64870 32488
rect 64994 32446 65038 32488
rect 65162 32446 65209 32488
rect 79943 32528 79990 32570
rect 80114 32528 80158 32570
rect 80282 32528 80329 32570
rect 79943 32488 79952 32528
rect 80114 32488 80116 32528
rect 80156 32488 80158 32528
rect 80320 32488 80329 32528
rect 79943 32446 79990 32488
rect 80114 32446 80158 32488
rect 80282 32446 80329 32488
rect 3103 31772 3150 31814
rect 3274 31772 3318 31814
rect 3442 31772 3489 31814
rect 3103 31732 3112 31772
rect 3274 31732 3276 31772
rect 3316 31732 3318 31772
rect 3480 31732 3489 31772
rect 3103 31690 3150 31732
rect 3274 31690 3318 31732
rect 3442 31690 3489 31732
rect 78703 31772 78750 31814
rect 78874 31772 78918 31814
rect 79042 31772 79089 31814
rect 78703 31732 78712 31772
rect 78874 31732 78876 31772
rect 78916 31732 78918 31772
rect 79080 31732 79089 31772
rect 78703 31690 78750 31732
rect 78874 31690 78918 31732
rect 79042 31690 79089 31732
rect 4343 31016 4390 31058
rect 4514 31016 4558 31058
rect 4682 31016 4729 31058
rect 4343 30976 4352 31016
rect 4514 30976 4516 31016
rect 4556 30976 4558 31016
rect 4720 30976 4729 31016
rect 4343 30934 4390 30976
rect 4514 30934 4558 30976
rect 4682 30934 4729 30976
rect 79943 31016 79990 31058
rect 80114 31016 80158 31058
rect 80282 31016 80329 31058
rect 79943 30976 79952 31016
rect 80114 30976 80116 31016
rect 80156 30976 80158 31016
rect 80320 30976 80329 31016
rect 79943 30934 79990 30976
rect 80114 30934 80158 30976
rect 80282 30934 80329 30976
rect 6403 30472 6412 30512
rect 6452 30472 97321 30512
rect 97361 30472 97370 30512
rect 3103 30260 3150 30302
rect 3274 30260 3318 30302
rect 3442 30260 3489 30302
rect 3103 30220 3112 30260
rect 3274 30220 3276 30260
rect 3316 30220 3318 30260
rect 3480 30220 3489 30260
rect 3103 30178 3150 30220
rect 3274 30178 3318 30220
rect 3442 30178 3489 30220
rect 78703 30260 78750 30302
rect 78874 30260 78918 30302
rect 79042 30260 79089 30302
rect 78703 30220 78712 30260
rect 78874 30220 78876 30260
rect 78916 30220 78918 30260
rect 79080 30220 79089 30260
rect 78703 30178 78750 30220
rect 78874 30178 78918 30220
rect 79042 30178 79089 30220
rect 4343 29504 4390 29546
rect 4514 29504 4558 29546
rect 4682 29504 4729 29546
rect 4343 29464 4352 29504
rect 4514 29464 4516 29504
rect 4556 29464 4558 29504
rect 4720 29464 4729 29504
rect 4343 29422 4390 29464
rect 4514 29422 4558 29464
rect 4682 29422 4729 29464
rect 79943 29504 79990 29546
rect 80114 29504 80158 29546
rect 80282 29504 80329 29546
rect 79943 29464 79952 29504
rect 80114 29464 80116 29504
rect 80156 29464 80158 29504
rect 80320 29464 80329 29504
rect 79943 29422 79990 29464
rect 80114 29422 80158 29464
rect 80282 29422 80329 29464
rect 95036 29062 95476 29136
rect 95036 28938 95110 29062
rect 95234 28938 95278 29062
rect 95402 28938 95476 29062
rect 95036 28894 95476 28938
rect 3103 28748 3150 28790
rect 3274 28748 3318 28790
rect 3442 28748 3489 28790
rect 3103 28708 3112 28748
rect 3274 28708 3276 28748
rect 3316 28708 3318 28748
rect 3480 28708 3489 28748
rect 61987 28708 61996 28748
rect 62036 28708 66386 28748
rect 3103 28666 3150 28708
rect 3274 28666 3318 28708
rect 3442 28666 3489 28708
rect 78703 28748 78750 28790
rect 78874 28748 78918 28790
rect 79042 28748 79089 28790
rect 78703 28708 78712 28748
rect 78874 28708 78876 28748
rect 78916 28708 78918 28748
rect 79080 28708 79089 28748
rect 78703 28666 78750 28708
rect 78874 28666 78918 28708
rect 79042 28666 79089 28708
rect 95036 28770 95110 28894
rect 95234 28770 95278 28894
rect 95402 28770 95476 28894
rect 95036 28696 95476 28770
rect 66211 28540 66220 28580
rect 66260 28540 67298 28580
rect 4343 27992 4390 28034
rect 4514 27992 4558 28034
rect 4682 27992 4729 28034
rect 4343 27952 4352 27992
rect 4514 27952 4516 27992
rect 4556 27952 4558 27992
rect 4720 27952 4729 27992
rect 4343 27910 4390 27952
rect 4514 27910 4558 27952
rect 4682 27910 4729 27952
rect 79943 27992 79990 28034
rect 80114 27992 80158 28034
rect 80282 27992 80329 28034
rect 79943 27952 79952 27992
rect 80114 27952 80116 27992
rect 80156 27952 80158 27992
rect 80320 27952 80329 27992
rect 79943 27910 79990 27952
rect 80114 27910 80158 27952
rect 80282 27910 80329 27952
rect 93796 27822 94236 27896
rect 93796 27698 93870 27822
rect 93994 27698 94038 27822
rect 94162 27698 94236 27822
rect 18196 27622 18636 27696
rect 18196 27498 18270 27622
rect 18394 27498 18438 27622
rect 18562 27498 18636 27622
rect 18196 27454 18636 27498
rect 18196 27330 18270 27454
rect 18394 27330 18438 27454
rect 18562 27330 18636 27454
rect 3103 27236 3150 27278
rect 3274 27236 3318 27278
rect 3442 27236 3489 27278
rect 18196 27256 18636 27330
rect 33316 27622 33756 27696
rect 33316 27498 33390 27622
rect 33514 27498 33558 27622
rect 33682 27498 33756 27622
rect 33316 27454 33756 27498
rect 33316 27330 33390 27454
rect 33514 27330 33558 27454
rect 33682 27330 33756 27454
rect 33316 27256 33756 27330
rect 48436 27622 48876 27696
rect 48436 27498 48510 27622
rect 48634 27498 48678 27622
rect 48802 27498 48876 27622
rect 48436 27454 48876 27498
rect 48436 27330 48510 27454
rect 48634 27330 48678 27454
rect 48802 27330 48876 27454
rect 48436 27256 48876 27330
rect 63556 27622 63996 27696
rect 63556 27498 63630 27622
rect 63754 27498 63798 27622
rect 63922 27498 63996 27622
rect 63556 27454 63996 27498
rect 93796 27654 94236 27698
rect 93796 27530 93870 27654
rect 93994 27530 94038 27654
rect 94162 27530 94236 27654
rect 93796 27456 94236 27530
rect 63556 27330 63630 27454
rect 63754 27330 63798 27454
rect 63922 27330 63996 27454
rect 63556 27256 63996 27330
rect 3103 27196 3112 27236
rect 3274 27196 3276 27236
rect 3316 27196 3318 27236
rect 3480 27196 3489 27236
rect 3103 27154 3150 27196
rect 3274 27154 3318 27196
rect 3442 27154 3489 27196
rect 78703 27236 78750 27278
rect 78874 27236 78918 27278
rect 79042 27236 79089 27278
rect 78703 27196 78712 27236
rect 78874 27196 78876 27236
rect 78916 27196 78918 27236
rect 79080 27196 79089 27236
rect 78703 27154 78750 27196
rect 78874 27154 78918 27196
rect 79042 27154 79089 27196
rect 4343 26480 4390 26522
rect 4514 26480 4558 26522
rect 4682 26480 4729 26522
rect 4343 26440 4352 26480
rect 4514 26440 4516 26480
rect 4556 26440 4558 26480
rect 4720 26440 4729 26480
rect 4343 26398 4390 26440
rect 4514 26398 4558 26440
rect 4682 26398 4729 26440
rect 79943 26480 79990 26522
rect 80114 26480 80158 26522
rect 80282 26480 80329 26522
rect 79943 26440 79952 26480
rect 80114 26440 80116 26480
rect 80156 26440 80158 26480
rect 80320 26440 80329 26480
rect 79943 26398 79990 26440
rect 80114 26398 80158 26440
rect 80282 26398 80329 26440
rect 3103 25724 3150 25766
rect 3274 25724 3318 25766
rect 3442 25724 3489 25766
rect 3103 25684 3112 25724
rect 3274 25684 3276 25724
rect 3316 25684 3318 25724
rect 3480 25684 3489 25724
rect 3103 25642 3150 25684
rect 3274 25642 3318 25684
rect 3442 25642 3489 25684
rect 78703 25724 78750 25766
rect 78874 25724 78918 25766
rect 79042 25724 79089 25766
rect 78703 25684 78712 25724
rect 78874 25684 78876 25724
rect 78916 25684 78918 25724
rect 79080 25684 79089 25724
rect 78703 25642 78750 25684
rect 78874 25642 78918 25684
rect 79042 25642 79089 25684
rect 4343 24968 4390 25010
rect 4514 24968 4558 25010
rect 4682 24968 4729 25010
rect 4343 24928 4352 24968
rect 4514 24928 4516 24968
rect 4556 24928 4558 24968
rect 4720 24928 4729 24968
rect 4343 24886 4390 24928
rect 4514 24886 4558 24928
rect 4682 24886 4729 24928
rect 79943 24968 79990 25010
rect 80114 24968 80158 25010
rect 80282 24968 80329 25010
rect 79943 24928 79952 24968
rect 80114 24928 80116 24968
rect 80156 24928 80158 24968
rect 80320 24928 80329 24968
rect 79943 24886 79990 24928
rect 80114 24886 80158 24928
rect 80282 24886 80329 24928
rect 3103 24212 3150 24254
rect 3274 24212 3318 24254
rect 3442 24212 3489 24254
rect 3103 24172 3112 24212
rect 3274 24172 3276 24212
rect 3316 24172 3318 24212
rect 3480 24172 3489 24212
rect 3103 24130 3150 24172
rect 3274 24130 3318 24172
rect 3442 24130 3489 24172
rect 78703 24212 78750 24254
rect 78874 24212 78918 24254
rect 79042 24212 79089 24254
rect 78703 24172 78712 24212
rect 78874 24172 78876 24212
rect 78916 24172 78918 24212
rect 79080 24172 79089 24212
rect 78703 24130 78750 24172
rect 78874 24130 78918 24172
rect 79042 24130 79089 24172
rect 4343 23456 4390 23498
rect 4514 23456 4558 23498
rect 4682 23456 4729 23498
rect 4343 23416 4352 23456
rect 4514 23416 4516 23456
rect 4556 23416 4558 23456
rect 4720 23416 4729 23456
rect 4343 23374 4390 23416
rect 4514 23374 4558 23416
rect 4682 23374 4729 23416
rect 79943 23456 79990 23498
rect 80114 23456 80158 23498
rect 80282 23456 80329 23498
rect 79943 23416 79952 23456
rect 80114 23416 80116 23456
rect 80156 23416 80158 23456
rect 80320 23416 80329 23456
rect 79943 23374 79990 23416
rect 80114 23374 80158 23416
rect 80282 23374 80329 23416
rect 19436 22862 19876 22936
rect 3103 22700 3150 22742
rect 3274 22700 3318 22742
rect 3442 22700 3489 22742
rect 3103 22660 3112 22700
rect 3274 22660 3276 22700
rect 3316 22660 3318 22700
rect 3480 22660 3489 22700
rect 3103 22618 3150 22660
rect 3274 22618 3318 22660
rect 3442 22618 3489 22660
rect 19436 22738 19510 22862
rect 19634 22738 19678 22862
rect 19802 22738 19876 22862
rect 19436 22694 19876 22738
rect 19436 22570 19510 22694
rect 19634 22570 19678 22694
rect 19802 22570 19876 22694
rect 19436 22496 19876 22570
rect 34556 22862 34996 22936
rect 34556 22738 34630 22862
rect 34754 22738 34798 22862
rect 34922 22738 34996 22862
rect 34556 22694 34996 22738
rect 34556 22570 34630 22694
rect 34754 22570 34798 22694
rect 34922 22570 34996 22694
rect 34556 22496 34996 22570
rect 49676 22862 50116 22936
rect 49676 22738 49750 22862
rect 49874 22738 49918 22862
rect 50042 22738 50116 22862
rect 49676 22694 50116 22738
rect 49676 22570 49750 22694
rect 49874 22570 49918 22694
rect 50042 22570 50116 22694
rect 49676 22496 50116 22570
rect 64796 22862 65236 22936
rect 64796 22738 64870 22862
rect 64994 22738 65038 22862
rect 65162 22738 65236 22862
rect 64796 22694 65236 22738
rect 64796 22570 64870 22694
rect 64994 22570 65038 22694
rect 65162 22570 65236 22694
rect 78703 22700 78750 22742
rect 78874 22700 78918 22742
rect 79042 22700 79089 22742
rect 78703 22660 78712 22700
rect 78874 22660 78876 22700
rect 78916 22660 78918 22700
rect 79080 22660 79089 22700
rect 78703 22618 78750 22660
rect 78874 22618 78918 22660
rect 79042 22618 79089 22660
rect 64796 22496 65236 22570
rect 4343 21944 4390 21986
rect 4514 21944 4558 21986
rect 4682 21944 4729 21986
rect 4343 21904 4352 21944
rect 4514 21904 4516 21944
rect 4556 21904 4558 21944
rect 4720 21904 4729 21944
rect 4343 21862 4390 21904
rect 4514 21862 4558 21904
rect 4682 21862 4729 21904
rect 79943 21944 79990 21986
rect 80114 21944 80158 21986
rect 80282 21944 80329 21986
rect 79943 21904 79952 21944
rect 80114 21904 80116 21944
rect 80156 21904 80158 21944
rect 80320 21904 80329 21944
rect 79943 21862 79990 21904
rect 80114 21862 80158 21904
rect 80282 21862 80329 21904
rect 95063 21944 95110 21986
rect 95234 21944 95278 21986
rect 95402 21944 95449 21986
rect 95063 21904 95072 21944
rect 95234 21904 95236 21944
rect 95276 21904 95278 21944
rect 95440 21904 95449 21944
rect 95063 21862 95110 21904
rect 95234 21862 95278 21904
rect 95402 21862 95449 21904
rect 18196 21622 18636 21696
rect 18196 21498 18270 21622
rect 18394 21498 18438 21622
rect 18562 21498 18636 21622
rect 18196 21454 18636 21498
rect 18196 21330 18270 21454
rect 18394 21330 18438 21454
rect 18562 21330 18636 21454
rect 18196 21256 18636 21330
rect 33316 21622 33756 21696
rect 33316 21498 33390 21622
rect 33514 21498 33558 21622
rect 33682 21498 33756 21622
rect 33316 21454 33756 21498
rect 33316 21330 33390 21454
rect 33514 21330 33558 21454
rect 33682 21330 33756 21454
rect 33316 21256 33756 21330
rect 48436 21622 48876 21696
rect 48436 21498 48510 21622
rect 48634 21498 48678 21622
rect 48802 21498 48876 21622
rect 48436 21454 48876 21498
rect 48436 21330 48510 21454
rect 48634 21330 48678 21454
rect 48802 21330 48876 21454
rect 48436 21256 48876 21330
rect 63556 21622 63996 21696
rect 63556 21498 63630 21622
rect 63754 21498 63798 21622
rect 63922 21498 63996 21622
rect 63556 21454 63996 21498
rect 63556 21330 63630 21454
rect 63754 21330 63798 21454
rect 63922 21330 63996 21454
rect 63556 21256 63996 21330
rect 3103 21188 3150 21230
rect 3274 21188 3318 21230
rect 3442 21188 3489 21230
rect 3103 21148 3112 21188
rect 3274 21148 3276 21188
rect 3316 21148 3318 21188
rect 3480 21148 3489 21188
rect 3103 21106 3150 21148
rect 3274 21106 3318 21148
rect 3442 21106 3489 21148
rect 78703 21188 78750 21230
rect 78874 21188 78918 21230
rect 79042 21188 79089 21230
rect 78703 21148 78712 21188
rect 78874 21148 78876 21188
rect 78916 21148 78918 21188
rect 79080 21148 79089 21188
rect 78703 21106 78750 21148
rect 78874 21106 78918 21148
rect 79042 21106 79089 21148
rect 93823 21188 93870 21230
rect 93994 21188 94038 21230
rect 94162 21188 94209 21230
rect 93823 21148 93832 21188
rect 93994 21148 93996 21188
rect 94036 21148 94038 21188
rect 94200 21148 94209 21188
rect 93823 21106 93870 21148
rect 93994 21106 94038 21148
rect 94162 21106 94209 21148
rect 4343 20432 4390 20474
rect 4514 20432 4558 20474
rect 4682 20432 4729 20474
rect 4343 20392 4352 20432
rect 4514 20392 4516 20432
rect 4556 20392 4558 20432
rect 4720 20392 4729 20432
rect 4343 20350 4390 20392
rect 4514 20350 4558 20392
rect 4682 20350 4729 20392
rect 79943 20432 79990 20474
rect 80114 20432 80158 20474
rect 80282 20432 80329 20474
rect 79943 20392 79952 20432
rect 80114 20392 80116 20432
rect 80156 20392 80158 20432
rect 80320 20392 80329 20432
rect 79943 20350 79990 20392
rect 80114 20350 80158 20392
rect 80282 20350 80329 20392
rect 95063 20432 95110 20474
rect 95234 20432 95278 20474
rect 95402 20432 95449 20474
rect 95063 20392 95072 20432
rect 95234 20392 95236 20432
rect 95276 20392 95278 20432
rect 95440 20392 95449 20432
rect 95063 20350 95110 20392
rect 95234 20350 95278 20392
rect 95402 20350 95449 20392
rect 3103 19676 3150 19718
rect 3274 19676 3318 19718
rect 3442 19676 3489 19718
rect 3103 19636 3112 19676
rect 3274 19636 3276 19676
rect 3316 19636 3318 19676
rect 3480 19636 3489 19676
rect 3103 19594 3150 19636
rect 3274 19594 3318 19636
rect 3442 19594 3489 19636
rect 78703 19676 78750 19718
rect 78874 19676 78918 19718
rect 79042 19676 79089 19718
rect 78703 19636 78712 19676
rect 78874 19636 78876 19676
rect 78916 19636 78918 19676
rect 79080 19636 79089 19676
rect 78703 19594 78750 19636
rect 78874 19594 78918 19636
rect 79042 19594 79089 19636
rect 93823 19676 93870 19718
rect 93994 19676 94038 19718
rect 94162 19676 94209 19718
rect 93823 19636 93832 19676
rect 93994 19636 93996 19676
rect 94036 19636 94038 19676
rect 94200 19636 94209 19676
rect 93823 19594 93870 19636
rect 93994 19594 94038 19636
rect 94162 19594 94209 19636
rect 4343 18920 4390 18962
rect 4514 18920 4558 18962
rect 4682 18920 4729 18962
rect 4343 18880 4352 18920
rect 4514 18880 4516 18920
rect 4556 18880 4558 18920
rect 4720 18880 4729 18920
rect 4343 18838 4390 18880
rect 4514 18838 4558 18880
rect 4682 18838 4729 18880
rect 79943 18920 79990 18962
rect 80114 18920 80158 18962
rect 80282 18920 80329 18962
rect 79943 18880 79952 18920
rect 80114 18880 80116 18920
rect 80156 18880 80158 18920
rect 80320 18880 80329 18920
rect 79943 18838 79990 18880
rect 80114 18838 80158 18880
rect 80282 18838 80329 18880
rect 3103 18164 3150 18206
rect 3274 18164 3318 18206
rect 3442 18164 3489 18206
rect 3103 18124 3112 18164
rect 3274 18124 3276 18164
rect 3316 18124 3318 18164
rect 3480 18124 3489 18164
rect 3103 18082 3150 18124
rect 3274 18082 3318 18124
rect 3442 18082 3489 18124
rect 78703 18164 78750 18206
rect 78874 18164 78918 18206
rect 79042 18164 79089 18206
rect 78703 18124 78712 18164
rect 78874 18124 78876 18164
rect 78916 18124 78918 18164
rect 79080 18124 79089 18164
rect 78703 18082 78750 18124
rect 78874 18082 78918 18124
rect 79042 18082 79089 18124
rect 4343 17408 4390 17450
rect 4514 17408 4558 17450
rect 4682 17408 4729 17450
rect 4343 17368 4352 17408
rect 4514 17368 4516 17408
rect 4556 17368 4558 17408
rect 4720 17368 4729 17408
rect 4343 17326 4390 17368
rect 4514 17326 4558 17368
rect 4682 17326 4729 17368
rect 79943 17408 79990 17450
rect 80114 17408 80158 17450
rect 80282 17408 80329 17450
rect 79943 17368 79952 17408
rect 80114 17368 80116 17408
rect 80156 17368 80158 17408
rect 80320 17368 80329 17408
rect 79943 17326 79990 17368
rect 80114 17326 80158 17368
rect 80282 17326 80329 17368
rect 19436 16862 19876 16936
rect 19436 16738 19510 16862
rect 19634 16738 19678 16862
rect 19802 16738 19876 16862
rect 19436 16694 19876 16738
rect 3103 16652 3150 16694
rect 3274 16652 3318 16694
rect 3442 16652 3489 16694
rect 3103 16612 3112 16652
rect 3274 16612 3276 16652
rect 3316 16612 3318 16652
rect 3480 16612 3489 16652
rect 3103 16570 3150 16612
rect 3274 16570 3318 16612
rect 3442 16570 3489 16612
rect 19436 16570 19510 16694
rect 19634 16570 19678 16694
rect 19802 16570 19876 16694
rect 19436 16496 19876 16570
rect 34556 16862 34996 16936
rect 34556 16738 34630 16862
rect 34754 16738 34798 16862
rect 34922 16738 34996 16862
rect 34556 16694 34996 16738
rect 34556 16570 34630 16694
rect 34754 16570 34798 16694
rect 34922 16570 34996 16694
rect 34556 16496 34996 16570
rect 49676 16862 50116 16936
rect 49676 16738 49750 16862
rect 49874 16738 49918 16862
rect 50042 16738 50116 16862
rect 49676 16694 50116 16738
rect 49676 16570 49750 16694
rect 49874 16570 49918 16694
rect 50042 16570 50116 16694
rect 49676 16496 50116 16570
rect 64796 16862 65236 16936
rect 64796 16738 64870 16862
rect 64994 16738 65038 16862
rect 65162 16738 65236 16862
rect 64796 16694 65236 16738
rect 64796 16570 64870 16694
rect 64994 16570 65038 16694
rect 65162 16570 65236 16694
rect 78703 16652 78750 16694
rect 78874 16652 78918 16694
rect 79042 16652 79089 16694
rect 78703 16612 78712 16652
rect 78874 16612 78876 16652
rect 78916 16612 78918 16652
rect 79080 16612 79089 16652
rect 78703 16570 78750 16612
rect 78874 16570 78918 16612
rect 79042 16570 79089 16612
rect 64796 16496 65236 16570
rect 4343 15896 4390 15938
rect 4514 15896 4558 15938
rect 4682 15896 4729 15938
rect 4343 15856 4352 15896
rect 4514 15856 4516 15896
rect 4556 15856 4558 15896
rect 4720 15856 4729 15896
rect 4343 15814 4390 15856
rect 4514 15814 4558 15856
rect 4682 15814 4729 15856
rect 79943 15896 79990 15938
rect 80114 15896 80158 15938
rect 80282 15896 80329 15938
rect 79943 15856 79952 15896
rect 80114 15856 80116 15896
rect 80156 15856 80158 15896
rect 80320 15856 80329 15896
rect 79943 15814 79990 15856
rect 80114 15814 80158 15856
rect 80282 15814 80329 15856
rect 18196 15622 18636 15696
rect 18196 15498 18270 15622
rect 18394 15498 18438 15622
rect 18562 15498 18636 15622
rect 18196 15454 18636 15498
rect 18196 15330 18270 15454
rect 18394 15330 18438 15454
rect 18562 15330 18636 15454
rect 18196 15256 18636 15330
rect 33316 15622 33756 15696
rect 33316 15498 33390 15622
rect 33514 15498 33558 15622
rect 33682 15498 33756 15622
rect 33316 15454 33756 15498
rect 33316 15330 33390 15454
rect 33514 15330 33558 15454
rect 33682 15330 33756 15454
rect 33316 15256 33756 15330
rect 48436 15622 48876 15696
rect 48436 15498 48510 15622
rect 48634 15498 48678 15622
rect 48802 15498 48876 15622
rect 48436 15454 48876 15498
rect 48436 15330 48510 15454
rect 48634 15330 48678 15454
rect 48802 15330 48876 15454
rect 48436 15256 48876 15330
rect 63556 15622 63996 15696
rect 63556 15498 63630 15622
rect 63754 15498 63798 15622
rect 63922 15498 63996 15622
rect 63556 15454 63996 15498
rect 63556 15330 63630 15454
rect 63754 15330 63798 15454
rect 63922 15330 63996 15454
rect 63556 15256 63996 15330
rect 3103 15140 3150 15182
rect 3274 15140 3318 15182
rect 3442 15140 3489 15182
rect 3103 15100 3112 15140
rect 3274 15100 3276 15140
rect 3316 15100 3318 15140
rect 3480 15100 3489 15140
rect 3103 15058 3150 15100
rect 3274 15058 3318 15100
rect 3442 15058 3489 15100
rect 78703 15140 78750 15182
rect 78874 15140 78918 15182
rect 79042 15140 79089 15182
rect 78703 15100 78712 15140
rect 78874 15100 78876 15140
rect 78916 15100 78918 15140
rect 79080 15100 79089 15140
rect 78703 15058 78750 15100
rect 78874 15058 78918 15100
rect 79042 15058 79089 15100
rect 4343 14384 4390 14426
rect 4514 14384 4558 14426
rect 4682 14384 4729 14426
rect 4343 14344 4352 14384
rect 4514 14344 4516 14384
rect 4556 14344 4558 14384
rect 4720 14344 4729 14384
rect 4343 14302 4390 14344
rect 4514 14302 4558 14344
rect 4682 14302 4729 14344
rect 79943 14384 79990 14426
rect 80114 14384 80158 14426
rect 80282 14384 80329 14426
rect 79943 14344 79952 14384
rect 80114 14344 80116 14384
rect 80156 14344 80158 14384
rect 80320 14344 80329 14384
rect 79943 14302 79990 14344
rect 80114 14302 80158 14344
rect 80282 14302 80329 14344
rect 3103 13628 3150 13670
rect 3274 13628 3318 13670
rect 3442 13628 3489 13670
rect 3103 13588 3112 13628
rect 3274 13588 3276 13628
rect 3316 13588 3318 13628
rect 3480 13588 3489 13628
rect 3103 13546 3150 13588
rect 3274 13546 3318 13588
rect 3442 13546 3489 13588
rect 78703 13628 78750 13670
rect 78874 13628 78918 13670
rect 79042 13628 79089 13670
rect 78703 13588 78712 13628
rect 78874 13588 78876 13628
rect 78916 13588 78918 13628
rect 79080 13588 79089 13628
rect 78703 13546 78750 13588
rect 78874 13546 78918 13588
rect 79042 13546 79089 13588
rect 4343 12872 4390 12914
rect 4514 12872 4558 12914
rect 4682 12872 4729 12914
rect 4343 12832 4352 12872
rect 4514 12832 4516 12872
rect 4556 12832 4558 12872
rect 4720 12832 4729 12872
rect 4343 12790 4390 12832
rect 4514 12790 4558 12832
rect 4682 12790 4729 12832
rect 79943 12872 79990 12914
rect 80114 12872 80158 12914
rect 80282 12872 80329 12914
rect 79943 12832 79952 12872
rect 80114 12832 80116 12872
rect 80156 12832 80158 12872
rect 80320 12832 80329 12872
rect 79943 12790 79990 12832
rect 80114 12790 80158 12832
rect 80282 12790 80329 12832
rect 3103 12116 3150 12158
rect 3274 12116 3318 12158
rect 3442 12116 3489 12158
rect 3103 12076 3112 12116
rect 3274 12076 3276 12116
rect 3316 12076 3318 12116
rect 3480 12076 3489 12116
rect 3103 12034 3150 12076
rect 3274 12034 3318 12076
rect 3442 12034 3489 12076
rect 78703 12116 78750 12158
rect 78874 12116 78918 12158
rect 79042 12116 79089 12158
rect 78703 12076 78712 12116
rect 78874 12076 78876 12116
rect 78916 12076 78918 12116
rect 79080 12076 79089 12116
rect 78703 12034 78750 12076
rect 78874 12034 78918 12076
rect 79042 12034 79089 12076
rect 95036 11862 95476 11936
rect 95036 11738 95110 11862
rect 95234 11738 95278 11862
rect 95402 11738 95476 11862
rect 95036 11694 95476 11738
rect 95036 11570 95110 11694
rect 95234 11570 95278 11694
rect 95402 11570 95476 11694
rect 95036 11496 95476 11570
rect 4343 11360 4390 11402
rect 4514 11360 4558 11402
rect 4682 11360 4729 11402
rect 4343 11320 4352 11360
rect 4514 11320 4516 11360
rect 4556 11320 4558 11360
rect 4720 11320 4729 11360
rect 4343 11278 4390 11320
rect 4514 11278 4558 11320
rect 4682 11278 4729 11320
rect 79943 11360 79990 11402
rect 80114 11360 80158 11402
rect 80282 11360 80329 11402
rect 79943 11320 79952 11360
rect 80114 11320 80116 11360
rect 80156 11320 80158 11360
rect 80320 11320 80329 11360
rect 79943 11278 79990 11320
rect 80114 11278 80158 11320
rect 80282 11278 80329 11320
rect 95683 11152 95692 11192
rect 95732 11152 99940 11192
rect 99980 11152 99989 11192
rect 19436 10862 19876 10936
rect 19436 10738 19510 10862
rect 19634 10738 19678 10862
rect 19802 10738 19876 10862
rect 19436 10694 19876 10738
rect 3103 10604 3150 10646
rect 3274 10604 3318 10646
rect 3442 10604 3489 10646
rect 3103 10564 3112 10604
rect 3274 10564 3276 10604
rect 3316 10564 3318 10604
rect 3480 10564 3489 10604
rect 3103 10522 3150 10564
rect 3274 10522 3318 10564
rect 3442 10522 3489 10564
rect 19436 10570 19510 10694
rect 19634 10570 19678 10694
rect 19802 10570 19876 10694
rect 19436 10496 19876 10570
rect 34556 10862 34996 10936
rect 34556 10738 34630 10862
rect 34754 10738 34798 10862
rect 34922 10738 34996 10862
rect 34556 10694 34996 10738
rect 34556 10570 34630 10694
rect 34754 10570 34798 10694
rect 34922 10570 34996 10694
rect 34556 10496 34996 10570
rect 49676 10862 50116 10936
rect 49676 10738 49750 10862
rect 49874 10738 49918 10862
rect 50042 10738 50116 10862
rect 49676 10694 50116 10738
rect 49676 10570 49750 10694
rect 49874 10570 49918 10694
rect 50042 10570 50116 10694
rect 49676 10496 50116 10570
rect 64796 10862 65236 10936
rect 64796 10738 64870 10862
rect 64994 10738 65038 10862
rect 65162 10738 65236 10862
rect 64796 10694 65236 10738
rect 64796 10570 64870 10694
rect 64994 10570 65038 10694
rect 65162 10570 65236 10694
rect 64796 10496 65236 10570
rect 78703 10604 78750 10646
rect 78874 10604 78918 10646
rect 79042 10604 79089 10646
rect 78703 10564 78712 10604
rect 78874 10564 78876 10604
rect 78916 10564 78918 10604
rect 79080 10564 79089 10604
rect 78703 10522 78750 10564
rect 78874 10522 78918 10564
rect 79042 10522 79089 10564
rect 93796 10622 94236 10696
rect 93796 10498 93870 10622
rect 93994 10498 94038 10622
rect 94162 10498 94236 10622
rect 93796 10454 94236 10498
rect 93796 10330 93870 10454
rect 93994 10330 94038 10454
rect 94162 10330 94236 10454
rect 93796 10256 94236 10330
rect 4343 9848 4390 9890
rect 4514 9848 4558 9890
rect 4682 9848 4729 9890
rect 4343 9808 4352 9848
rect 4514 9808 4516 9848
rect 4556 9808 4558 9848
rect 4720 9808 4729 9848
rect 4343 9766 4390 9808
rect 4514 9766 4558 9808
rect 4682 9766 4729 9808
rect 79943 9848 79990 9890
rect 80114 9848 80158 9890
rect 80282 9848 80329 9890
rect 79943 9808 79952 9848
rect 80114 9808 80116 9848
rect 80156 9808 80158 9848
rect 80320 9808 80329 9848
rect 79943 9766 79990 9808
rect 80114 9766 80158 9808
rect 80282 9766 80329 9808
rect 18196 9622 18636 9696
rect 18196 9498 18270 9622
rect 18394 9498 18438 9622
rect 18562 9498 18636 9622
rect 18196 9454 18636 9498
rect 18196 9330 18270 9454
rect 18394 9330 18438 9454
rect 18562 9330 18636 9454
rect 18196 9256 18636 9330
rect 33316 9622 33756 9696
rect 33316 9498 33390 9622
rect 33514 9498 33558 9622
rect 33682 9498 33756 9622
rect 33316 9454 33756 9498
rect 33316 9330 33390 9454
rect 33514 9330 33558 9454
rect 33682 9330 33756 9454
rect 33316 9256 33756 9330
rect 48436 9622 48876 9696
rect 48436 9498 48510 9622
rect 48634 9498 48678 9622
rect 48802 9498 48876 9622
rect 48436 9454 48876 9498
rect 48436 9330 48510 9454
rect 48634 9330 48678 9454
rect 48802 9330 48876 9454
rect 48436 9256 48876 9330
rect 63556 9622 63996 9696
rect 63556 9498 63630 9622
rect 63754 9498 63798 9622
rect 63922 9498 63996 9622
rect 63556 9454 63996 9498
rect 63556 9330 63630 9454
rect 63754 9330 63798 9454
rect 63922 9330 63996 9454
rect 63556 9256 63996 9330
rect 3103 9092 3150 9134
rect 3274 9092 3318 9134
rect 3442 9092 3489 9134
rect 3103 9052 3112 9092
rect 3274 9052 3276 9092
rect 3316 9052 3318 9092
rect 3480 9052 3489 9092
rect 3103 9010 3150 9052
rect 3274 9010 3318 9052
rect 3442 9010 3489 9052
rect 78703 9092 78750 9134
rect 78874 9092 78918 9134
rect 79042 9092 79089 9134
rect 78703 9052 78712 9092
rect 78874 9052 78876 9092
rect 78916 9052 78918 9092
rect 79080 9052 79089 9092
rect 78703 9010 78750 9052
rect 78874 9010 78918 9052
rect 79042 9010 79089 9052
rect 87820 8968 99921 9008
rect 99961 8968 99970 9008
rect 87820 8924 87860 8968
rect 73027 8884 73036 8924
rect 73076 8884 87860 8924
rect 83491 8800 83500 8840
rect 83540 8800 87860 8840
rect 87820 8756 87860 8800
rect 87820 8716 99929 8756
rect 99969 8716 99978 8756
rect 4343 8336 4390 8378
rect 4514 8336 4558 8378
rect 4682 8336 4729 8378
rect 4343 8296 4352 8336
rect 4514 8296 4516 8336
rect 4556 8296 4558 8336
rect 4720 8296 4729 8336
rect 4343 8254 4390 8296
rect 4514 8254 4558 8296
rect 4682 8254 4729 8296
rect 79943 8336 79990 8378
rect 80114 8336 80158 8378
rect 80282 8336 80329 8378
rect 79943 8296 79952 8336
rect 80114 8296 80116 8336
rect 80156 8296 80158 8336
rect 80320 8296 80329 8336
rect 79943 8254 79990 8296
rect 80114 8254 80158 8296
rect 80282 8254 80329 8296
rect 3103 7580 3150 7622
rect 3274 7580 3318 7622
rect 3442 7580 3489 7622
rect 3103 7540 3112 7580
rect 3274 7540 3276 7580
rect 3316 7540 3318 7580
rect 3480 7540 3489 7580
rect 3103 7498 3150 7540
rect 3274 7498 3318 7540
rect 3442 7498 3489 7540
rect 78703 7580 78750 7622
rect 78874 7580 78918 7622
rect 79042 7580 79089 7622
rect 78703 7540 78712 7580
rect 78874 7540 78876 7580
rect 78916 7540 78918 7580
rect 79080 7540 79089 7580
rect 78703 7498 78750 7540
rect 78874 7498 78918 7540
rect 79042 7498 79089 7540
rect 4343 6824 4390 6866
rect 4514 6824 4558 6866
rect 4682 6824 4729 6866
rect 4343 6784 4352 6824
rect 4514 6784 4516 6824
rect 4556 6784 4558 6824
rect 4720 6784 4729 6824
rect 4343 6742 4390 6784
rect 4514 6742 4558 6784
rect 4682 6742 4729 6784
rect 79943 6824 79990 6866
rect 80114 6824 80158 6866
rect 80282 6824 80329 6866
rect 79943 6784 79952 6824
rect 80114 6784 80116 6824
rect 80156 6784 80158 6824
rect 80320 6784 80329 6824
rect 79943 6742 79990 6784
rect 80114 6742 80158 6784
rect 80282 6742 80329 6784
rect 3103 6068 3150 6110
rect 3274 6068 3318 6110
rect 3442 6068 3489 6110
rect 78703 6068 78750 6110
rect 78874 6068 78918 6110
rect 79042 6068 79089 6110
rect 3103 6028 3112 6068
rect 3274 6028 3276 6068
rect 3316 6028 3318 6068
rect 3480 6028 3489 6068
rect 26851 6028 26860 6068
rect 26900 6028 72748 6068
rect 72788 6028 72797 6068
rect 78703 6028 78712 6068
rect 78874 6028 78876 6068
rect 78916 6028 78918 6068
rect 79080 6028 79089 6068
rect 93571 6028 93580 6068
rect 93620 6028 99940 6068
rect 99980 6028 99989 6068
rect 3103 5986 3150 6028
rect 3274 5986 3318 6028
rect 3442 5986 3489 6028
rect 78703 5986 78750 6028
rect 78874 5986 78918 6028
rect 79042 5986 79089 6028
rect 95036 5862 95476 5936
rect 95036 5738 95110 5862
rect 95234 5738 95278 5862
rect 95402 5738 95476 5862
rect 1795 5692 1804 5732
rect 1844 5692 82924 5732
rect 82964 5692 82973 5732
rect 95036 5694 95476 5738
rect 1699 5608 1708 5648
rect 1748 5608 76972 5648
rect 77012 5608 77021 5648
rect 95036 5570 95110 5694
rect 95234 5570 95278 5694
rect 95402 5570 95476 5694
rect 95036 5496 95476 5570
rect 4343 5312 4390 5354
rect 4514 5312 4558 5354
rect 4682 5312 4729 5354
rect 4343 5272 4352 5312
rect 4514 5272 4516 5312
rect 4556 5272 4558 5312
rect 4720 5272 4729 5312
rect 4343 5230 4390 5272
rect 4514 5230 4558 5272
rect 4682 5230 4729 5272
rect 79943 5312 79990 5354
rect 80114 5312 80158 5354
rect 80282 5312 80329 5354
rect 79943 5272 79952 5312
rect 80114 5272 80116 5312
rect 80156 5272 80158 5312
rect 80320 5272 80329 5312
rect 79943 5230 79990 5272
rect 80114 5230 80158 5272
rect 80282 5230 80329 5272
rect 55747 5020 55756 5060
rect 55796 5020 66386 5060
rect 93796 4622 94236 4696
rect 3103 4556 3150 4598
rect 3274 4556 3318 4598
rect 3442 4556 3489 4598
rect 3103 4516 3112 4556
rect 3274 4516 3276 4556
rect 3316 4516 3318 4556
rect 3480 4516 3489 4556
rect 3103 4474 3150 4516
rect 3274 4474 3318 4516
rect 3442 4474 3489 4516
rect 78703 4556 78750 4598
rect 78874 4556 78918 4598
rect 79042 4556 79089 4598
rect 78703 4516 78712 4556
rect 78874 4516 78876 4556
rect 78916 4516 78918 4556
rect 79080 4516 79089 4556
rect 63331 4432 63340 4472
rect 63380 4432 67298 4472
rect 78703 4474 78750 4516
rect 78874 4474 78918 4516
rect 79042 4474 79089 4516
rect 93796 4498 93870 4622
rect 93994 4498 94038 4622
rect 94162 4498 94236 4622
rect 93796 4454 94236 4498
rect 93796 4330 93870 4454
rect 93994 4330 94038 4454
rect 94162 4330 94236 4454
rect 93796 4256 94236 4330
rect 4343 3800 4390 3842
rect 4514 3800 4558 3842
rect 4682 3800 4729 3842
rect 4343 3760 4352 3800
rect 4514 3760 4516 3800
rect 4556 3760 4558 3800
rect 4720 3760 4729 3800
rect 4343 3718 4390 3760
rect 4514 3718 4558 3760
rect 4682 3718 4729 3760
rect 19463 3800 19510 3842
rect 19634 3800 19678 3842
rect 19802 3800 19849 3842
rect 19463 3760 19472 3800
rect 19634 3760 19636 3800
rect 19676 3760 19678 3800
rect 19840 3760 19849 3800
rect 19463 3718 19510 3760
rect 19634 3718 19678 3760
rect 19802 3718 19849 3760
rect 34583 3800 34630 3842
rect 34754 3800 34798 3842
rect 34922 3800 34969 3842
rect 34583 3760 34592 3800
rect 34754 3760 34756 3800
rect 34796 3760 34798 3800
rect 34960 3760 34969 3800
rect 34583 3718 34630 3760
rect 34754 3718 34798 3760
rect 34922 3718 34969 3760
rect 49703 3800 49750 3842
rect 49874 3800 49918 3842
rect 50042 3800 50089 3842
rect 49703 3760 49712 3800
rect 49874 3760 49876 3800
rect 49916 3760 49918 3800
rect 50080 3760 50089 3800
rect 49703 3718 49750 3760
rect 49874 3718 49918 3760
rect 50042 3718 50089 3760
rect 64823 3800 64870 3842
rect 64994 3800 65038 3842
rect 65162 3800 65209 3842
rect 64823 3760 64832 3800
rect 64994 3760 64996 3800
rect 65036 3760 65038 3800
rect 65200 3760 65209 3800
rect 64823 3718 64870 3760
rect 64994 3718 65038 3760
rect 65162 3718 65209 3760
rect 79943 3800 79990 3842
rect 80114 3800 80158 3842
rect 80282 3800 80329 3842
rect 79943 3760 79952 3800
rect 80114 3760 80116 3800
rect 80156 3760 80158 3800
rect 80320 3760 80329 3800
rect 79943 3718 79990 3760
rect 80114 3718 80158 3760
rect 80282 3718 80329 3760
rect 37219 3592 37228 3632
rect 37268 3592 43220 3632
rect 43180 3548 43220 3592
rect 43180 3508 95692 3548
rect 95732 3508 95741 3548
rect 33955 3424 33964 3464
rect 34004 3424 93580 3464
rect 93620 3424 93629 3464
rect 3103 3044 3150 3086
rect 3274 3044 3318 3086
rect 3442 3044 3489 3086
rect 3103 3004 3112 3044
rect 3274 3004 3276 3044
rect 3316 3004 3318 3044
rect 3480 3004 3489 3044
rect 3103 2962 3150 3004
rect 3274 2962 3318 3004
rect 3442 2962 3489 3004
rect 18223 3044 18270 3086
rect 18394 3044 18438 3086
rect 18562 3044 18609 3086
rect 18223 3004 18232 3044
rect 18394 3004 18396 3044
rect 18436 3004 18438 3044
rect 18600 3004 18609 3044
rect 18223 2962 18270 3004
rect 18394 2962 18438 3004
rect 18562 2962 18609 3004
rect 33343 3044 33390 3086
rect 33514 3044 33558 3086
rect 33682 3044 33729 3086
rect 33343 3004 33352 3044
rect 33514 3004 33516 3044
rect 33556 3004 33558 3044
rect 33720 3004 33729 3044
rect 33343 2962 33390 3004
rect 33514 2962 33558 3004
rect 33682 2962 33729 3004
rect 48463 3044 48510 3086
rect 48634 3044 48678 3086
rect 48802 3044 48849 3086
rect 48463 3004 48472 3044
rect 48634 3004 48636 3044
rect 48676 3004 48678 3044
rect 48840 3004 48849 3044
rect 48463 2962 48510 3004
rect 48634 2962 48678 3004
rect 48802 2962 48849 3004
rect 63583 3044 63630 3086
rect 63754 3044 63798 3086
rect 63922 3044 63969 3086
rect 63583 3004 63592 3044
rect 63754 3004 63756 3044
rect 63796 3004 63798 3044
rect 63960 3004 63969 3044
rect 63583 2962 63630 3004
rect 63754 2962 63798 3004
rect 63922 2962 63969 3004
rect 78703 3044 78750 3086
rect 78874 3044 78918 3086
rect 79042 3044 79089 3086
rect 78703 3004 78712 3044
rect 78874 3004 78876 3044
rect 78916 3004 78918 3044
rect 79080 3004 79089 3044
rect 78703 2962 78750 3004
rect 78874 2962 78918 3004
rect 79042 2962 79089 3004
rect 4343 2288 4390 2330
rect 4514 2288 4558 2330
rect 4682 2288 4729 2330
rect 4343 2248 4352 2288
rect 4514 2248 4516 2288
rect 4556 2248 4558 2288
rect 4720 2248 4729 2288
rect 4343 2206 4390 2248
rect 4514 2206 4558 2248
rect 4682 2206 4729 2248
rect 19463 2288 19510 2330
rect 19634 2288 19678 2330
rect 19802 2288 19849 2330
rect 19463 2248 19472 2288
rect 19634 2248 19636 2288
rect 19676 2248 19678 2288
rect 19840 2248 19849 2288
rect 19463 2206 19510 2248
rect 19634 2206 19678 2248
rect 19802 2206 19849 2248
rect 34583 2288 34630 2330
rect 34754 2288 34798 2330
rect 34922 2288 34969 2330
rect 34583 2248 34592 2288
rect 34754 2248 34756 2288
rect 34796 2248 34798 2288
rect 34960 2248 34969 2288
rect 34583 2206 34630 2248
rect 34754 2206 34798 2248
rect 34922 2206 34969 2248
rect 49703 2288 49750 2330
rect 49874 2288 49918 2330
rect 50042 2288 50089 2330
rect 49703 2248 49712 2288
rect 49874 2248 49876 2288
rect 49916 2248 49918 2288
rect 50080 2248 50089 2288
rect 49703 2206 49750 2248
rect 49874 2206 49918 2248
rect 50042 2206 50089 2248
rect 64823 2288 64870 2330
rect 64994 2288 65038 2330
rect 65162 2288 65209 2330
rect 64823 2248 64832 2288
rect 64994 2248 64996 2288
rect 65036 2248 65038 2288
rect 65200 2248 65209 2288
rect 64823 2206 64870 2248
rect 64994 2206 65038 2248
rect 65162 2206 65209 2248
rect 79943 2288 79990 2330
rect 80114 2288 80158 2330
rect 80282 2288 80329 2330
rect 79943 2248 79952 2288
rect 80114 2248 80116 2288
rect 80156 2248 80158 2288
rect 80320 2248 80329 2288
rect 79943 2206 79990 2248
rect 80114 2206 80158 2248
rect 80282 2206 80329 2248
rect 3103 1532 3150 1574
rect 3274 1532 3318 1574
rect 3442 1532 3489 1574
rect 3103 1492 3112 1532
rect 3274 1492 3276 1532
rect 3316 1492 3318 1532
rect 3480 1492 3489 1532
rect 3103 1450 3150 1492
rect 3274 1450 3318 1492
rect 3442 1450 3489 1492
rect 18223 1532 18270 1574
rect 18394 1532 18438 1574
rect 18562 1532 18609 1574
rect 18223 1492 18232 1532
rect 18394 1492 18396 1532
rect 18436 1492 18438 1532
rect 18600 1492 18609 1532
rect 18223 1450 18270 1492
rect 18394 1450 18438 1492
rect 18562 1450 18609 1492
rect 33343 1532 33390 1574
rect 33514 1532 33558 1574
rect 33682 1532 33729 1574
rect 33343 1492 33352 1532
rect 33514 1492 33516 1532
rect 33556 1492 33558 1532
rect 33720 1492 33729 1532
rect 33343 1450 33390 1492
rect 33514 1450 33558 1492
rect 33682 1450 33729 1492
rect 48463 1532 48510 1574
rect 48634 1532 48678 1574
rect 48802 1532 48849 1574
rect 48463 1492 48472 1532
rect 48634 1492 48636 1532
rect 48676 1492 48678 1532
rect 48840 1492 48849 1532
rect 48463 1450 48510 1492
rect 48634 1450 48678 1492
rect 48802 1450 48849 1492
rect 63583 1532 63630 1574
rect 63754 1532 63798 1574
rect 63922 1532 63969 1574
rect 63583 1492 63592 1532
rect 63754 1492 63756 1532
rect 63796 1492 63798 1532
rect 63960 1492 63969 1532
rect 63583 1450 63630 1492
rect 63754 1450 63798 1492
rect 63922 1450 63969 1492
rect 78703 1532 78750 1574
rect 78874 1532 78918 1574
rect 79042 1532 79089 1574
rect 78703 1492 78712 1532
rect 78874 1492 78876 1532
rect 78916 1492 78918 1532
rect 79080 1492 79089 1532
rect 78703 1450 78750 1492
rect 78874 1450 78918 1492
rect 79042 1450 79089 1492
rect 4343 776 4390 818
rect 4514 776 4558 818
rect 4682 776 4729 818
rect 4343 736 4352 776
rect 4514 736 4516 776
rect 4556 736 4558 776
rect 4720 736 4729 776
rect 4343 694 4390 736
rect 4514 694 4558 736
rect 4682 694 4729 736
rect 19463 776 19510 818
rect 19634 776 19678 818
rect 19802 776 19849 818
rect 19463 736 19472 776
rect 19634 736 19636 776
rect 19676 736 19678 776
rect 19840 736 19849 776
rect 19463 694 19510 736
rect 19634 694 19678 736
rect 19802 694 19849 736
rect 34583 776 34630 818
rect 34754 776 34798 818
rect 34922 776 34969 818
rect 34583 736 34592 776
rect 34754 736 34756 776
rect 34796 736 34798 776
rect 34960 736 34969 776
rect 34583 694 34630 736
rect 34754 694 34798 736
rect 34922 694 34969 736
rect 49703 776 49750 818
rect 49874 776 49918 818
rect 50042 776 50089 818
rect 49703 736 49712 776
rect 49874 736 49876 776
rect 49916 736 49918 776
rect 50080 736 50089 776
rect 49703 694 49750 736
rect 49874 694 49918 736
rect 50042 694 50089 736
rect 64823 776 64870 818
rect 64994 776 65038 818
rect 65162 776 65209 818
rect 64823 736 64832 776
rect 64994 736 64996 776
rect 65036 736 65038 776
rect 65200 736 65209 776
rect 64823 694 64870 736
rect 64994 694 65038 736
rect 65162 694 65209 736
rect 79943 776 79990 818
rect 80114 776 80158 818
rect 80282 776 80329 818
rect 79943 736 79952 776
rect 80114 736 80116 776
rect 80156 736 80158 776
rect 80320 736 80329 776
rect 79943 694 79990 736
rect 80114 694 80158 736
rect 80282 694 80329 736
<< via5 >>
rect 4390 38576 4514 38618
rect 4558 38576 4682 38618
rect 4390 38536 4392 38576
rect 4392 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4514 38576
rect 4558 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4680 38576
rect 4680 38536 4682 38576
rect 4390 38494 4514 38536
rect 4558 38494 4682 38536
rect 19510 38576 19634 38618
rect 19678 38576 19802 38618
rect 19510 38536 19512 38576
rect 19512 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19634 38576
rect 19678 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19800 38576
rect 19800 38536 19802 38576
rect 19510 38494 19634 38536
rect 19678 38494 19802 38536
rect 34630 38576 34754 38618
rect 34798 38576 34922 38618
rect 34630 38536 34632 38576
rect 34632 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34754 38576
rect 34798 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34920 38576
rect 34920 38536 34922 38576
rect 34630 38494 34754 38536
rect 34798 38494 34922 38536
rect 49750 38576 49874 38618
rect 49918 38576 50042 38618
rect 49750 38536 49752 38576
rect 49752 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49874 38576
rect 49918 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50040 38576
rect 50040 38536 50042 38576
rect 49750 38494 49874 38536
rect 49918 38494 50042 38536
rect 64870 38576 64994 38618
rect 65038 38576 65162 38618
rect 64870 38536 64872 38576
rect 64872 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64994 38576
rect 65038 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65160 38576
rect 65160 38536 65162 38576
rect 64870 38494 64994 38536
rect 65038 38494 65162 38536
rect 79990 38576 80114 38618
rect 80158 38576 80282 38618
rect 79990 38536 79992 38576
rect 79992 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80114 38576
rect 80158 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80280 38576
rect 80280 38536 80282 38576
rect 79990 38494 80114 38536
rect 80158 38494 80282 38536
rect 3150 37820 3274 37862
rect 3318 37820 3442 37862
rect 3150 37780 3152 37820
rect 3152 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3274 37820
rect 3318 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3440 37820
rect 3440 37780 3442 37820
rect 3150 37738 3274 37780
rect 3318 37738 3442 37780
rect 18270 37820 18394 37862
rect 18438 37820 18562 37862
rect 18270 37780 18272 37820
rect 18272 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18394 37820
rect 18438 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18560 37820
rect 18560 37780 18562 37820
rect 18270 37738 18394 37780
rect 18438 37738 18562 37780
rect 33390 37820 33514 37862
rect 33558 37820 33682 37862
rect 33390 37780 33392 37820
rect 33392 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33514 37820
rect 33558 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33680 37820
rect 33680 37780 33682 37820
rect 33390 37738 33514 37780
rect 33558 37738 33682 37780
rect 48510 37820 48634 37862
rect 48678 37820 48802 37862
rect 48510 37780 48512 37820
rect 48512 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48634 37820
rect 48678 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48800 37820
rect 48800 37780 48802 37820
rect 48510 37738 48634 37780
rect 48678 37738 48802 37780
rect 63630 37820 63754 37862
rect 63798 37820 63922 37862
rect 63630 37780 63632 37820
rect 63632 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63754 37820
rect 63798 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63920 37820
rect 63920 37780 63922 37820
rect 63630 37738 63754 37780
rect 63798 37738 63922 37780
rect 78750 37820 78874 37862
rect 78918 37820 79042 37862
rect 78750 37780 78752 37820
rect 78752 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78874 37820
rect 78918 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79040 37820
rect 79040 37780 79042 37820
rect 78750 37738 78874 37780
rect 78918 37738 79042 37780
rect 4390 37064 4514 37106
rect 4558 37064 4682 37106
rect 4390 37024 4392 37064
rect 4392 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4514 37064
rect 4558 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4680 37064
rect 4680 37024 4682 37064
rect 4390 36982 4514 37024
rect 4558 36982 4682 37024
rect 19510 37064 19634 37106
rect 19678 37064 19802 37106
rect 19510 37024 19512 37064
rect 19512 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19634 37064
rect 19678 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19800 37064
rect 19800 37024 19802 37064
rect 19510 36982 19634 37024
rect 19678 36982 19802 37024
rect 34630 37064 34754 37106
rect 34798 37064 34922 37106
rect 34630 37024 34632 37064
rect 34632 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34754 37064
rect 34798 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34920 37064
rect 34920 37024 34922 37064
rect 34630 36982 34754 37024
rect 34798 36982 34922 37024
rect 49750 37064 49874 37106
rect 49918 37064 50042 37106
rect 49750 37024 49752 37064
rect 49752 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49874 37064
rect 49918 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50040 37064
rect 50040 37024 50042 37064
rect 49750 36982 49874 37024
rect 49918 36982 50042 37024
rect 64870 37064 64994 37106
rect 65038 37064 65162 37106
rect 64870 37024 64872 37064
rect 64872 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64994 37064
rect 65038 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65160 37064
rect 65160 37024 65162 37064
rect 64870 36982 64994 37024
rect 65038 36982 65162 37024
rect 79990 37064 80114 37106
rect 80158 37064 80282 37106
rect 79990 37024 79992 37064
rect 79992 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80114 37064
rect 80158 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80280 37064
rect 80280 37024 80282 37064
rect 79990 36982 80114 37024
rect 80158 36982 80282 37024
rect 3150 36308 3274 36350
rect 3318 36308 3442 36350
rect 3150 36268 3152 36308
rect 3152 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3274 36308
rect 3318 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3440 36308
rect 3440 36268 3442 36308
rect 3150 36226 3274 36268
rect 3318 36226 3442 36268
rect 18270 36308 18394 36350
rect 18438 36308 18562 36350
rect 18270 36268 18272 36308
rect 18272 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18394 36308
rect 18438 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18560 36308
rect 18560 36268 18562 36308
rect 18270 36226 18394 36268
rect 18438 36226 18562 36268
rect 33390 36308 33514 36350
rect 33558 36308 33682 36350
rect 33390 36268 33392 36308
rect 33392 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33514 36308
rect 33558 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33680 36308
rect 33680 36268 33682 36308
rect 33390 36226 33514 36268
rect 33558 36226 33682 36268
rect 48510 36308 48634 36350
rect 48678 36308 48802 36350
rect 48510 36268 48512 36308
rect 48512 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48634 36308
rect 48678 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48800 36308
rect 48800 36268 48802 36308
rect 48510 36226 48634 36268
rect 48678 36226 48802 36268
rect 63630 36308 63754 36350
rect 63798 36308 63922 36350
rect 63630 36268 63632 36308
rect 63632 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63754 36308
rect 63798 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63920 36308
rect 63920 36268 63922 36308
rect 63630 36226 63754 36268
rect 63798 36226 63922 36268
rect 78750 36308 78874 36350
rect 78918 36308 79042 36350
rect 78750 36268 78752 36308
rect 78752 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78874 36308
rect 78918 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79040 36308
rect 79040 36268 79042 36308
rect 78750 36226 78874 36268
rect 78918 36226 79042 36268
rect 4390 35552 4514 35594
rect 4558 35552 4682 35594
rect 4390 35512 4392 35552
rect 4392 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4514 35552
rect 4558 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4680 35552
rect 4680 35512 4682 35552
rect 4390 35470 4514 35512
rect 4558 35470 4682 35512
rect 19510 35552 19634 35594
rect 19678 35552 19802 35594
rect 19510 35512 19512 35552
rect 19512 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19634 35552
rect 19678 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19800 35552
rect 19800 35512 19802 35552
rect 19510 35470 19634 35512
rect 19678 35470 19802 35512
rect 34630 35552 34754 35594
rect 34798 35552 34922 35594
rect 34630 35512 34632 35552
rect 34632 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34754 35552
rect 34798 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34920 35552
rect 34920 35512 34922 35552
rect 34630 35470 34754 35512
rect 34798 35470 34922 35512
rect 49750 35552 49874 35594
rect 49918 35552 50042 35594
rect 49750 35512 49752 35552
rect 49752 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49874 35552
rect 49918 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50040 35552
rect 50040 35512 50042 35552
rect 49750 35470 49874 35512
rect 49918 35470 50042 35512
rect 64870 35552 64994 35594
rect 65038 35552 65162 35594
rect 64870 35512 64872 35552
rect 64872 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64994 35552
rect 65038 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65160 35552
rect 65160 35512 65162 35552
rect 64870 35470 64994 35512
rect 65038 35470 65162 35512
rect 79990 35552 80114 35594
rect 80158 35552 80282 35594
rect 79990 35512 79992 35552
rect 79992 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80114 35552
rect 80158 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80280 35552
rect 80280 35512 80282 35552
rect 79990 35470 80114 35512
rect 80158 35470 80282 35512
rect 3150 34796 3274 34838
rect 3318 34796 3442 34838
rect 3150 34756 3152 34796
rect 3152 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3274 34796
rect 3318 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3440 34796
rect 3440 34756 3442 34796
rect 3150 34714 3274 34756
rect 3318 34714 3442 34756
rect 18270 34796 18394 34838
rect 18438 34796 18562 34838
rect 18270 34756 18272 34796
rect 18272 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18394 34796
rect 18438 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18560 34796
rect 18560 34756 18562 34796
rect 18270 34714 18394 34756
rect 18438 34714 18562 34756
rect 33390 34796 33514 34838
rect 33558 34796 33682 34838
rect 33390 34756 33392 34796
rect 33392 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33514 34796
rect 33558 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33680 34796
rect 33680 34756 33682 34796
rect 33390 34714 33514 34756
rect 33558 34714 33682 34756
rect 48510 34796 48634 34838
rect 48678 34796 48802 34838
rect 48510 34756 48512 34796
rect 48512 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48634 34796
rect 48678 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48800 34796
rect 48800 34756 48802 34796
rect 48510 34714 48634 34756
rect 48678 34714 48802 34756
rect 63630 34796 63754 34838
rect 63798 34796 63922 34838
rect 63630 34756 63632 34796
rect 63632 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63754 34796
rect 63798 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63920 34796
rect 63920 34756 63922 34796
rect 63630 34714 63754 34756
rect 63798 34714 63922 34756
rect 78750 34796 78874 34838
rect 78918 34796 79042 34838
rect 78750 34756 78752 34796
rect 78752 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78874 34796
rect 78918 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79040 34796
rect 79040 34756 79042 34796
rect 78750 34714 78874 34756
rect 78918 34714 79042 34756
rect 4390 34040 4514 34082
rect 4558 34040 4682 34082
rect 4390 34000 4392 34040
rect 4392 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4514 34040
rect 4558 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4680 34040
rect 4680 34000 4682 34040
rect 4390 33958 4514 34000
rect 4558 33958 4682 34000
rect 19510 34040 19634 34082
rect 19678 34040 19802 34082
rect 19510 34000 19512 34040
rect 19512 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19634 34040
rect 19678 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19800 34040
rect 19800 34000 19802 34040
rect 19510 33958 19634 34000
rect 19678 33958 19802 34000
rect 34630 34040 34754 34082
rect 34798 34040 34922 34082
rect 34630 34000 34632 34040
rect 34632 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34754 34040
rect 34798 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34920 34040
rect 34920 34000 34922 34040
rect 34630 33958 34754 34000
rect 34798 33958 34922 34000
rect 49750 34040 49874 34082
rect 49918 34040 50042 34082
rect 49750 34000 49752 34040
rect 49752 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49874 34040
rect 49918 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50040 34040
rect 50040 34000 50042 34040
rect 49750 33958 49874 34000
rect 49918 33958 50042 34000
rect 64870 34040 64994 34082
rect 65038 34040 65162 34082
rect 64870 34000 64872 34040
rect 64872 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64994 34040
rect 65038 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65160 34040
rect 65160 34000 65162 34040
rect 64870 33958 64994 34000
rect 65038 33958 65162 34000
rect 79990 34040 80114 34082
rect 80158 34040 80282 34082
rect 79990 34000 79992 34040
rect 79992 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80114 34040
rect 80158 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80280 34040
rect 80280 34000 80282 34040
rect 79990 33958 80114 34000
rect 80158 33958 80282 34000
rect 93870 33698 93994 33822
rect 94038 33698 94162 33822
rect 93870 33530 93994 33654
rect 94038 33530 94162 33654
rect 3150 33284 3274 33326
rect 3318 33284 3442 33326
rect 3150 33244 3152 33284
rect 3152 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3274 33284
rect 3318 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3440 33284
rect 3440 33244 3442 33284
rect 3150 33202 3274 33244
rect 3318 33202 3442 33244
rect 18270 33284 18394 33326
rect 18438 33284 18562 33326
rect 18270 33244 18272 33284
rect 18272 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18394 33284
rect 18438 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18560 33284
rect 18560 33244 18562 33284
rect 18270 33202 18394 33244
rect 18438 33202 18562 33244
rect 33390 33284 33514 33326
rect 33558 33284 33682 33326
rect 33390 33244 33392 33284
rect 33392 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33514 33284
rect 33558 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33680 33284
rect 33680 33244 33682 33284
rect 33390 33202 33514 33244
rect 33558 33202 33682 33244
rect 48510 33284 48634 33326
rect 48678 33284 48802 33326
rect 48510 33244 48512 33284
rect 48512 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48634 33284
rect 48678 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48800 33284
rect 48800 33244 48802 33284
rect 48510 33202 48634 33244
rect 48678 33202 48802 33244
rect 63630 33284 63754 33326
rect 63798 33284 63922 33326
rect 63630 33244 63632 33284
rect 63632 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63754 33284
rect 63798 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63920 33284
rect 63920 33244 63922 33284
rect 63630 33202 63754 33244
rect 63798 33202 63922 33244
rect 78750 33284 78874 33326
rect 78918 33284 79042 33326
rect 78750 33244 78752 33284
rect 78752 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78874 33284
rect 78918 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79040 33284
rect 79040 33244 79042 33284
rect 78750 33202 78874 33244
rect 78918 33202 79042 33244
rect 4390 32528 4514 32570
rect 4558 32528 4682 32570
rect 4390 32488 4392 32528
rect 4392 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4514 32528
rect 4558 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4680 32528
rect 4680 32488 4682 32528
rect 4390 32446 4514 32488
rect 4558 32446 4682 32488
rect 19510 32528 19634 32570
rect 19678 32528 19802 32570
rect 19510 32488 19512 32528
rect 19512 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19634 32528
rect 19678 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19800 32528
rect 19800 32488 19802 32528
rect 19510 32446 19634 32488
rect 19678 32446 19802 32488
rect 34630 32528 34754 32570
rect 34798 32528 34922 32570
rect 34630 32488 34632 32528
rect 34632 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34754 32528
rect 34798 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34920 32528
rect 34920 32488 34922 32528
rect 34630 32446 34754 32488
rect 34798 32446 34922 32488
rect 49750 32528 49874 32570
rect 49918 32528 50042 32570
rect 49750 32488 49752 32528
rect 49752 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49874 32528
rect 49918 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50040 32528
rect 50040 32488 50042 32528
rect 49750 32446 49874 32488
rect 49918 32446 50042 32488
rect 64870 32528 64994 32570
rect 65038 32528 65162 32570
rect 64870 32488 64872 32528
rect 64872 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64994 32528
rect 65038 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65160 32528
rect 65160 32488 65162 32528
rect 64870 32446 64994 32488
rect 65038 32446 65162 32488
rect 79990 32528 80114 32570
rect 80158 32528 80282 32570
rect 79990 32488 79992 32528
rect 79992 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80114 32528
rect 80158 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80280 32528
rect 80280 32488 80282 32528
rect 79990 32446 80114 32488
rect 80158 32446 80282 32488
rect 3150 31772 3274 31814
rect 3318 31772 3442 31814
rect 3150 31732 3152 31772
rect 3152 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3274 31772
rect 3318 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3440 31772
rect 3440 31732 3442 31772
rect 3150 31690 3274 31732
rect 3318 31690 3442 31732
rect 78750 31772 78874 31814
rect 78918 31772 79042 31814
rect 78750 31732 78752 31772
rect 78752 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78874 31772
rect 78918 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79040 31772
rect 79040 31732 79042 31772
rect 78750 31690 78874 31732
rect 78918 31690 79042 31732
rect 4390 31016 4514 31058
rect 4558 31016 4682 31058
rect 4390 30976 4392 31016
rect 4392 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4514 31016
rect 4558 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4680 31016
rect 4680 30976 4682 31016
rect 4390 30934 4514 30976
rect 4558 30934 4682 30976
rect 79990 31016 80114 31058
rect 80158 31016 80282 31058
rect 79990 30976 79992 31016
rect 79992 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80114 31016
rect 80158 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80280 31016
rect 80280 30976 80282 31016
rect 79990 30934 80114 30976
rect 80158 30934 80282 30976
rect 3150 30260 3274 30302
rect 3318 30260 3442 30302
rect 3150 30220 3152 30260
rect 3152 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3274 30260
rect 3318 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3440 30260
rect 3440 30220 3442 30260
rect 3150 30178 3274 30220
rect 3318 30178 3442 30220
rect 78750 30260 78874 30302
rect 78918 30260 79042 30302
rect 78750 30220 78752 30260
rect 78752 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78874 30260
rect 78918 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79040 30260
rect 79040 30220 79042 30260
rect 78750 30178 78874 30220
rect 78918 30178 79042 30220
rect 4390 29504 4514 29546
rect 4558 29504 4682 29546
rect 4390 29464 4392 29504
rect 4392 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4514 29504
rect 4558 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4680 29504
rect 4680 29464 4682 29504
rect 4390 29422 4514 29464
rect 4558 29422 4682 29464
rect 79990 29504 80114 29546
rect 80158 29504 80282 29546
rect 79990 29464 79992 29504
rect 79992 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80114 29504
rect 80158 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80280 29504
rect 80280 29464 80282 29504
rect 79990 29422 80114 29464
rect 80158 29422 80282 29464
rect 95110 28938 95234 29062
rect 95278 28938 95402 29062
rect 3150 28748 3274 28790
rect 3318 28748 3442 28790
rect 3150 28708 3152 28748
rect 3152 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3274 28748
rect 3318 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3440 28748
rect 3440 28708 3442 28748
rect 3150 28666 3274 28708
rect 3318 28666 3442 28708
rect 66386 28666 66510 28790
rect 78750 28748 78874 28790
rect 78918 28748 79042 28790
rect 78750 28708 78752 28748
rect 78752 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78874 28748
rect 78918 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79040 28748
rect 79040 28708 79042 28748
rect 78750 28666 78874 28708
rect 78918 28666 79042 28708
rect 95110 28770 95234 28894
rect 95278 28770 95402 28894
rect 67298 28498 67422 28622
rect 4390 27992 4514 28034
rect 4558 27992 4682 28034
rect 4390 27952 4392 27992
rect 4392 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4514 27992
rect 4558 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4680 27992
rect 4680 27952 4682 27992
rect 4390 27910 4514 27952
rect 4558 27910 4682 27952
rect 79990 27992 80114 28034
rect 80158 27992 80282 28034
rect 79990 27952 79992 27992
rect 79992 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80114 27992
rect 80158 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80280 27992
rect 80280 27952 80282 27992
rect 79990 27910 80114 27952
rect 80158 27910 80282 27952
rect 93870 27698 93994 27822
rect 94038 27698 94162 27822
rect 18270 27498 18394 27622
rect 18438 27498 18562 27622
rect 18270 27330 18394 27454
rect 18438 27330 18562 27454
rect 3150 27236 3274 27278
rect 3318 27236 3442 27278
rect 33390 27498 33514 27622
rect 33558 27498 33682 27622
rect 33390 27330 33514 27454
rect 33558 27330 33682 27454
rect 48510 27498 48634 27622
rect 48678 27498 48802 27622
rect 48510 27330 48634 27454
rect 48678 27330 48802 27454
rect 63630 27498 63754 27622
rect 63798 27498 63922 27622
rect 93870 27530 93994 27654
rect 94038 27530 94162 27654
rect 63630 27330 63754 27454
rect 63798 27330 63922 27454
rect 3150 27196 3152 27236
rect 3152 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3274 27236
rect 3318 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3440 27236
rect 3440 27196 3442 27236
rect 3150 27154 3274 27196
rect 3318 27154 3442 27196
rect 78750 27236 78874 27278
rect 78918 27236 79042 27278
rect 78750 27196 78752 27236
rect 78752 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78874 27236
rect 78918 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79040 27236
rect 79040 27196 79042 27236
rect 78750 27154 78874 27196
rect 78918 27154 79042 27196
rect 4390 26480 4514 26522
rect 4558 26480 4682 26522
rect 4390 26440 4392 26480
rect 4392 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4514 26480
rect 4558 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4680 26480
rect 4680 26440 4682 26480
rect 4390 26398 4514 26440
rect 4558 26398 4682 26440
rect 79990 26480 80114 26522
rect 80158 26480 80282 26522
rect 79990 26440 79992 26480
rect 79992 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80114 26480
rect 80158 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80280 26480
rect 80280 26440 80282 26480
rect 79990 26398 80114 26440
rect 80158 26398 80282 26440
rect 3150 25724 3274 25766
rect 3318 25724 3442 25766
rect 3150 25684 3152 25724
rect 3152 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3274 25724
rect 3318 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3440 25724
rect 3440 25684 3442 25724
rect 3150 25642 3274 25684
rect 3318 25642 3442 25684
rect 78750 25724 78874 25766
rect 78918 25724 79042 25766
rect 78750 25684 78752 25724
rect 78752 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78874 25724
rect 78918 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79040 25724
rect 79040 25684 79042 25724
rect 78750 25642 78874 25684
rect 78918 25642 79042 25684
rect 4390 24968 4514 25010
rect 4558 24968 4682 25010
rect 4390 24928 4392 24968
rect 4392 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4514 24968
rect 4558 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4680 24968
rect 4680 24928 4682 24968
rect 4390 24886 4514 24928
rect 4558 24886 4682 24928
rect 79990 24968 80114 25010
rect 80158 24968 80282 25010
rect 79990 24928 79992 24968
rect 79992 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80114 24968
rect 80158 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80280 24968
rect 80280 24928 80282 24968
rect 79990 24886 80114 24928
rect 80158 24886 80282 24928
rect 3150 24212 3274 24254
rect 3318 24212 3442 24254
rect 3150 24172 3152 24212
rect 3152 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3274 24212
rect 3318 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3440 24212
rect 3440 24172 3442 24212
rect 3150 24130 3274 24172
rect 3318 24130 3442 24172
rect 78750 24212 78874 24254
rect 78918 24212 79042 24254
rect 78750 24172 78752 24212
rect 78752 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78874 24212
rect 78918 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79040 24212
rect 79040 24172 79042 24212
rect 78750 24130 78874 24172
rect 78918 24130 79042 24172
rect 4390 23456 4514 23498
rect 4558 23456 4682 23498
rect 4390 23416 4392 23456
rect 4392 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4514 23456
rect 4558 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4680 23456
rect 4680 23416 4682 23456
rect 4390 23374 4514 23416
rect 4558 23374 4682 23416
rect 79990 23456 80114 23498
rect 80158 23456 80282 23498
rect 79990 23416 79992 23456
rect 79992 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80114 23456
rect 80158 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80280 23456
rect 80280 23416 80282 23456
rect 79990 23374 80114 23416
rect 80158 23374 80282 23416
rect 3150 22700 3274 22742
rect 3318 22700 3442 22742
rect 3150 22660 3152 22700
rect 3152 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3274 22700
rect 3318 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3440 22700
rect 3440 22660 3442 22700
rect 3150 22618 3274 22660
rect 3318 22618 3442 22660
rect 19510 22738 19634 22862
rect 19678 22738 19802 22862
rect 19510 22570 19634 22694
rect 19678 22570 19802 22694
rect 34630 22738 34754 22862
rect 34798 22738 34922 22862
rect 34630 22570 34754 22694
rect 34798 22570 34922 22694
rect 49750 22738 49874 22862
rect 49918 22738 50042 22862
rect 49750 22570 49874 22694
rect 49918 22570 50042 22694
rect 64870 22738 64994 22862
rect 65038 22738 65162 22862
rect 64870 22570 64994 22694
rect 65038 22570 65162 22694
rect 78750 22700 78874 22742
rect 78918 22700 79042 22742
rect 78750 22660 78752 22700
rect 78752 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78874 22700
rect 78918 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79040 22700
rect 79040 22660 79042 22700
rect 78750 22618 78874 22660
rect 78918 22618 79042 22660
rect 4390 21944 4514 21986
rect 4558 21944 4682 21986
rect 4390 21904 4392 21944
rect 4392 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4514 21944
rect 4558 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4680 21944
rect 4680 21904 4682 21944
rect 4390 21862 4514 21904
rect 4558 21862 4682 21904
rect 79990 21944 80114 21986
rect 80158 21944 80282 21986
rect 79990 21904 79992 21944
rect 79992 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80114 21944
rect 80158 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80280 21944
rect 80280 21904 80282 21944
rect 79990 21862 80114 21904
rect 80158 21862 80282 21904
rect 95110 21944 95234 21986
rect 95278 21944 95402 21986
rect 95110 21904 95112 21944
rect 95112 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95234 21944
rect 95278 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95400 21944
rect 95400 21904 95402 21944
rect 95110 21862 95234 21904
rect 95278 21862 95402 21904
rect 18270 21498 18394 21622
rect 18438 21498 18562 21622
rect 18270 21330 18394 21454
rect 18438 21330 18562 21454
rect 33390 21498 33514 21622
rect 33558 21498 33682 21622
rect 33390 21330 33514 21454
rect 33558 21330 33682 21454
rect 48510 21498 48634 21622
rect 48678 21498 48802 21622
rect 48510 21330 48634 21454
rect 48678 21330 48802 21454
rect 63630 21498 63754 21622
rect 63798 21498 63922 21622
rect 63630 21330 63754 21454
rect 63798 21330 63922 21454
rect 3150 21188 3274 21230
rect 3318 21188 3442 21230
rect 3150 21148 3152 21188
rect 3152 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3274 21188
rect 3318 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3440 21188
rect 3440 21148 3442 21188
rect 3150 21106 3274 21148
rect 3318 21106 3442 21148
rect 78750 21188 78874 21230
rect 78918 21188 79042 21230
rect 78750 21148 78752 21188
rect 78752 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78874 21188
rect 78918 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79040 21188
rect 79040 21148 79042 21188
rect 78750 21106 78874 21148
rect 78918 21106 79042 21148
rect 93870 21188 93994 21230
rect 94038 21188 94162 21230
rect 93870 21148 93872 21188
rect 93872 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93994 21188
rect 94038 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94160 21188
rect 94160 21148 94162 21188
rect 93870 21106 93994 21148
rect 94038 21106 94162 21148
rect 4390 20432 4514 20474
rect 4558 20432 4682 20474
rect 4390 20392 4392 20432
rect 4392 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4514 20432
rect 4558 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4680 20432
rect 4680 20392 4682 20432
rect 4390 20350 4514 20392
rect 4558 20350 4682 20392
rect 79990 20432 80114 20474
rect 80158 20432 80282 20474
rect 79990 20392 79992 20432
rect 79992 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80114 20432
rect 80158 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80280 20432
rect 80280 20392 80282 20432
rect 79990 20350 80114 20392
rect 80158 20350 80282 20392
rect 95110 20432 95234 20474
rect 95278 20432 95402 20474
rect 95110 20392 95112 20432
rect 95112 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95234 20432
rect 95278 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95400 20432
rect 95400 20392 95402 20432
rect 95110 20350 95234 20392
rect 95278 20350 95402 20392
rect 3150 19676 3274 19718
rect 3318 19676 3442 19718
rect 3150 19636 3152 19676
rect 3152 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3274 19676
rect 3318 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3440 19676
rect 3440 19636 3442 19676
rect 3150 19594 3274 19636
rect 3318 19594 3442 19636
rect 78750 19676 78874 19718
rect 78918 19676 79042 19718
rect 78750 19636 78752 19676
rect 78752 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78874 19676
rect 78918 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79040 19676
rect 79040 19636 79042 19676
rect 78750 19594 78874 19636
rect 78918 19594 79042 19636
rect 93870 19676 93994 19718
rect 94038 19676 94162 19718
rect 93870 19636 93872 19676
rect 93872 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93994 19676
rect 94038 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94160 19676
rect 94160 19636 94162 19676
rect 93870 19594 93994 19636
rect 94038 19594 94162 19636
rect 4390 18920 4514 18962
rect 4558 18920 4682 18962
rect 4390 18880 4392 18920
rect 4392 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4514 18920
rect 4558 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4680 18920
rect 4680 18880 4682 18920
rect 4390 18838 4514 18880
rect 4558 18838 4682 18880
rect 79990 18920 80114 18962
rect 80158 18920 80282 18962
rect 79990 18880 79992 18920
rect 79992 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80114 18920
rect 80158 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80280 18920
rect 80280 18880 80282 18920
rect 79990 18838 80114 18880
rect 80158 18838 80282 18880
rect 3150 18164 3274 18206
rect 3318 18164 3442 18206
rect 3150 18124 3152 18164
rect 3152 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3274 18164
rect 3318 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3440 18164
rect 3440 18124 3442 18164
rect 3150 18082 3274 18124
rect 3318 18082 3442 18124
rect 78750 18164 78874 18206
rect 78918 18164 79042 18206
rect 78750 18124 78752 18164
rect 78752 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78874 18164
rect 78918 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79040 18164
rect 79040 18124 79042 18164
rect 78750 18082 78874 18124
rect 78918 18082 79042 18124
rect 4390 17408 4514 17450
rect 4558 17408 4682 17450
rect 4390 17368 4392 17408
rect 4392 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4514 17408
rect 4558 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4680 17408
rect 4680 17368 4682 17408
rect 4390 17326 4514 17368
rect 4558 17326 4682 17368
rect 79990 17408 80114 17450
rect 80158 17408 80282 17450
rect 79990 17368 79992 17408
rect 79992 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80114 17408
rect 80158 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80280 17408
rect 80280 17368 80282 17408
rect 79990 17326 80114 17368
rect 80158 17326 80282 17368
rect 19510 16738 19634 16862
rect 19678 16738 19802 16862
rect 3150 16652 3274 16694
rect 3318 16652 3442 16694
rect 3150 16612 3152 16652
rect 3152 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3274 16652
rect 3318 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3440 16652
rect 3440 16612 3442 16652
rect 3150 16570 3274 16612
rect 3318 16570 3442 16612
rect 19510 16570 19634 16694
rect 19678 16570 19802 16694
rect 34630 16738 34754 16862
rect 34798 16738 34922 16862
rect 34630 16570 34754 16694
rect 34798 16570 34922 16694
rect 49750 16738 49874 16862
rect 49918 16738 50042 16862
rect 49750 16570 49874 16694
rect 49918 16570 50042 16694
rect 64870 16738 64994 16862
rect 65038 16738 65162 16862
rect 64870 16570 64994 16694
rect 65038 16570 65162 16694
rect 78750 16652 78874 16694
rect 78918 16652 79042 16694
rect 78750 16612 78752 16652
rect 78752 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78874 16652
rect 78918 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79040 16652
rect 79040 16612 79042 16652
rect 78750 16570 78874 16612
rect 78918 16570 79042 16612
rect 4390 15896 4514 15938
rect 4558 15896 4682 15938
rect 4390 15856 4392 15896
rect 4392 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4514 15896
rect 4558 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4680 15896
rect 4680 15856 4682 15896
rect 4390 15814 4514 15856
rect 4558 15814 4682 15856
rect 79990 15896 80114 15938
rect 80158 15896 80282 15938
rect 79990 15856 79992 15896
rect 79992 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80114 15896
rect 80158 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80280 15896
rect 80280 15856 80282 15896
rect 79990 15814 80114 15856
rect 80158 15814 80282 15856
rect 18270 15498 18394 15622
rect 18438 15498 18562 15622
rect 18270 15330 18394 15454
rect 18438 15330 18562 15454
rect 33390 15498 33514 15622
rect 33558 15498 33682 15622
rect 33390 15330 33514 15454
rect 33558 15330 33682 15454
rect 48510 15498 48634 15622
rect 48678 15498 48802 15622
rect 48510 15330 48634 15454
rect 48678 15330 48802 15454
rect 63630 15498 63754 15622
rect 63798 15498 63922 15622
rect 63630 15330 63754 15454
rect 63798 15330 63922 15454
rect 3150 15140 3274 15182
rect 3318 15140 3442 15182
rect 3150 15100 3152 15140
rect 3152 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3274 15140
rect 3318 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3440 15140
rect 3440 15100 3442 15140
rect 3150 15058 3274 15100
rect 3318 15058 3442 15100
rect 78750 15140 78874 15182
rect 78918 15140 79042 15182
rect 78750 15100 78752 15140
rect 78752 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78874 15140
rect 78918 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79040 15140
rect 79040 15100 79042 15140
rect 78750 15058 78874 15100
rect 78918 15058 79042 15100
rect 4390 14384 4514 14426
rect 4558 14384 4682 14426
rect 4390 14344 4392 14384
rect 4392 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4514 14384
rect 4558 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4680 14384
rect 4680 14344 4682 14384
rect 4390 14302 4514 14344
rect 4558 14302 4682 14344
rect 79990 14384 80114 14426
rect 80158 14384 80282 14426
rect 79990 14344 79992 14384
rect 79992 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80114 14384
rect 80158 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80280 14384
rect 80280 14344 80282 14384
rect 79990 14302 80114 14344
rect 80158 14302 80282 14344
rect 3150 13628 3274 13670
rect 3318 13628 3442 13670
rect 3150 13588 3152 13628
rect 3152 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3274 13628
rect 3318 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3440 13628
rect 3440 13588 3442 13628
rect 3150 13546 3274 13588
rect 3318 13546 3442 13588
rect 78750 13628 78874 13670
rect 78918 13628 79042 13670
rect 78750 13588 78752 13628
rect 78752 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78874 13628
rect 78918 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79040 13628
rect 79040 13588 79042 13628
rect 78750 13546 78874 13588
rect 78918 13546 79042 13588
rect 4390 12872 4514 12914
rect 4558 12872 4682 12914
rect 4390 12832 4392 12872
rect 4392 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4514 12872
rect 4558 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4680 12872
rect 4680 12832 4682 12872
rect 4390 12790 4514 12832
rect 4558 12790 4682 12832
rect 79990 12872 80114 12914
rect 80158 12872 80282 12914
rect 79990 12832 79992 12872
rect 79992 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80114 12872
rect 80158 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80280 12872
rect 80280 12832 80282 12872
rect 79990 12790 80114 12832
rect 80158 12790 80282 12832
rect 3150 12116 3274 12158
rect 3318 12116 3442 12158
rect 3150 12076 3152 12116
rect 3152 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3274 12116
rect 3318 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3440 12116
rect 3440 12076 3442 12116
rect 3150 12034 3274 12076
rect 3318 12034 3442 12076
rect 78750 12116 78874 12158
rect 78918 12116 79042 12158
rect 78750 12076 78752 12116
rect 78752 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78874 12116
rect 78918 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79040 12116
rect 79040 12076 79042 12116
rect 78750 12034 78874 12076
rect 78918 12034 79042 12076
rect 95110 11738 95234 11862
rect 95278 11738 95402 11862
rect 95110 11570 95234 11694
rect 95278 11570 95402 11694
rect 4390 11360 4514 11402
rect 4558 11360 4682 11402
rect 4390 11320 4392 11360
rect 4392 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4514 11360
rect 4558 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4680 11360
rect 4680 11320 4682 11360
rect 4390 11278 4514 11320
rect 4558 11278 4682 11320
rect 79990 11360 80114 11402
rect 80158 11360 80282 11402
rect 79990 11320 79992 11360
rect 79992 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80114 11360
rect 80158 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80280 11360
rect 80280 11320 80282 11360
rect 79990 11278 80114 11320
rect 80158 11278 80282 11320
rect 19510 10738 19634 10862
rect 19678 10738 19802 10862
rect 3150 10604 3274 10646
rect 3318 10604 3442 10646
rect 3150 10564 3152 10604
rect 3152 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3274 10604
rect 3318 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3440 10604
rect 3440 10564 3442 10604
rect 3150 10522 3274 10564
rect 3318 10522 3442 10564
rect 19510 10570 19634 10694
rect 19678 10570 19802 10694
rect 34630 10738 34754 10862
rect 34798 10738 34922 10862
rect 34630 10570 34754 10694
rect 34798 10570 34922 10694
rect 49750 10738 49874 10862
rect 49918 10738 50042 10862
rect 49750 10570 49874 10694
rect 49918 10570 50042 10694
rect 64870 10738 64994 10862
rect 65038 10738 65162 10862
rect 64870 10570 64994 10694
rect 65038 10570 65162 10694
rect 78750 10604 78874 10646
rect 78918 10604 79042 10646
rect 78750 10564 78752 10604
rect 78752 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78874 10604
rect 78918 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79040 10604
rect 79040 10564 79042 10604
rect 78750 10522 78874 10564
rect 78918 10522 79042 10564
rect 93870 10498 93994 10622
rect 94038 10498 94162 10622
rect 93870 10330 93994 10454
rect 94038 10330 94162 10454
rect 4390 9848 4514 9890
rect 4558 9848 4682 9890
rect 4390 9808 4392 9848
rect 4392 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4514 9848
rect 4558 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4680 9848
rect 4680 9808 4682 9848
rect 4390 9766 4514 9808
rect 4558 9766 4682 9808
rect 79990 9848 80114 9890
rect 80158 9848 80282 9890
rect 79990 9808 79992 9848
rect 79992 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80114 9848
rect 80158 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80280 9848
rect 80280 9808 80282 9848
rect 79990 9766 80114 9808
rect 80158 9766 80282 9808
rect 18270 9498 18394 9622
rect 18438 9498 18562 9622
rect 18270 9330 18394 9454
rect 18438 9330 18562 9454
rect 33390 9498 33514 9622
rect 33558 9498 33682 9622
rect 33390 9330 33514 9454
rect 33558 9330 33682 9454
rect 48510 9498 48634 9622
rect 48678 9498 48802 9622
rect 48510 9330 48634 9454
rect 48678 9330 48802 9454
rect 63630 9498 63754 9622
rect 63798 9498 63922 9622
rect 63630 9330 63754 9454
rect 63798 9330 63922 9454
rect 3150 9092 3274 9134
rect 3318 9092 3442 9134
rect 3150 9052 3152 9092
rect 3152 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3274 9092
rect 3318 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3440 9092
rect 3440 9052 3442 9092
rect 3150 9010 3274 9052
rect 3318 9010 3442 9052
rect 78750 9092 78874 9134
rect 78918 9092 79042 9134
rect 78750 9052 78752 9092
rect 78752 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78874 9092
rect 78918 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79040 9092
rect 79040 9052 79042 9092
rect 78750 9010 78874 9052
rect 78918 9010 79042 9052
rect 4390 8336 4514 8378
rect 4558 8336 4682 8378
rect 4390 8296 4392 8336
rect 4392 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4514 8336
rect 4558 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4680 8336
rect 4680 8296 4682 8336
rect 4390 8254 4514 8296
rect 4558 8254 4682 8296
rect 79990 8336 80114 8378
rect 80158 8336 80282 8378
rect 79990 8296 79992 8336
rect 79992 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80114 8336
rect 80158 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80280 8336
rect 80280 8296 80282 8336
rect 79990 8254 80114 8296
rect 80158 8254 80282 8296
rect 3150 7580 3274 7622
rect 3318 7580 3442 7622
rect 3150 7540 3152 7580
rect 3152 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3274 7580
rect 3318 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3440 7580
rect 3440 7540 3442 7580
rect 3150 7498 3274 7540
rect 3318 7498 3442 7540
rect 78750 7580 78874 7622
rect 78918 7580 79042 7622
rect 78750 7540 78752 7580
rect 78752 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78874 7580
rect 78918 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79040 7580
rect 79040 7540 79042 7580
rect 78750 7498 78874 7540
rect 78918 7498 79042 7540
rect 4390 6824 4514 6866
rect 4558 6824 4682 6866
rect 4390 6784 4392 6824
rect 4392 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4514 6824
rect 4558 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4680 6824
rect 4680 6784 4682 6824
rect 4390 6742 4514 6784
rect 4558 6742 4682 6784
rect 79990 6824 80114 6866
rect 80158 6824 80282 6866
rect 79990 6784 79992 6824
rect 79992 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80114 6824
rect 80158 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80280 6824
rect 80280 6784 80282 6824
rect 79990 6742 80114 6784
rect 80158 6742 80282 6784
rect 3150 6068 3274 6110
rect 3318 6068 3442 6110
rect 78750 6068 78874 6110
rect 78918 6068 79042 6110
rect 3150 6028 3152 6068
rect 3152 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3274 6068
rect 3318 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3440 6068
rect 3440 6028 3442 6068
rect 78750 6028 78752 6068
rect 78752 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78874 6068
rect 78918 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79040 6068
rect 79040 6028 79042 6068
rect 3150 5986 3274 6028
rect 3318 5986 3442 6028
rect 78750 5986 78874 6028
rect 78918 5986 79042 6028
rect 95110 5738 95234 5862
rect 95278 5738 95402 5862
rect 95110 5570 95234 5694
rect 95278 5570 95402 5694
rect 4390 5312 4514 5354
rect 4558 5312 4682 5354
rect 4390 5272 4392 5312
rect 4392 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4514 5312
rect 4558 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4680 5312
rect 4680 5272 4682 5312
rect 4390 5230 4514 5272
rect 4558 5230 4682 5272
rect 79990 5312 80114 5354
rect 80158 5312 80282 5354
rect 79990 5272 79992 5312
rect 79992 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80114 5312
rect 80158 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80280 5312
rect 80280 5272 80282 5312
rect 79990 5230 80114 5272
rect 80158 5230 80282 5272
rect 66386 4978 66510 5102
rect 3150 4556 3274 4598
rect 3318 4556 3442 4598
rect 3150 4516 3152 4556
rect 3152 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3274 4556
rect 3318 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3440 4556
rect 3440 4516 3442 4556
rect 3150 4474 3274 4516
rect 3318 4474 3442 4516
rect 78750 4556 78874 4598
rect 78918 4556 79042 4598
rect 78750 4516 78752 4556
rect 78752 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78874 4556
rect 78918 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79040 4556
rect 79040 4516 79042 4556
rect 67298 4390 67422 4514
rect 78750 4474 78874 4516
rect 78918 4474 79042 4516
rect 93870 4498 93994 4622
rect 94038 4498 94162 4622
rect 93870 4330 93994 4454
rect 94038 4330 94162 4454
rect 4390 3800 4514 3842
rect 4558 3800 4682 3842
rect 4390 3760 4392 3800
rect 4392 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4514 3800
rect 4558 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4680 3800
rect 4680 3760 4682 3800
rect 4390 3718 4514 3760
rect 4558 3718 4682 3760
rect 19510 3800 19634 3842
rect 19678 3800 19802 3842
rect 19510 3760 19512 3800
rect 19512 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19634 3800
rect 19678 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19800 3800
rect 19800 3760 19802 3800
rect 19510 3718 19634 3760
rect 19678 3718 19802 3760
rect 34630 3800 34754 3842
rect 34798 3800 34922 3842
rect 34630 3760 34632 3800
rect 34632 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34754 3800
rect 34798 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34920 3800
rect 34920 3760 34922 3800
rect 34630 3718 34754 3760
rect 34798 3718 34922 3760
rect 49750 3800 49874 3842
rect 49918 3800 50042 3842
rect 49750 3760 49752 3800
rect 49752 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49874 3800
rect 49918 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50040 3800
rect 50040 3760 50042 3800
rect 49750 3718 49874 3760
rect 49918 3718 50042 3760
rect 64870 3800 64994 3842
rect 65038 3800 65162 3842
rect 64870 3760 64872 3800
rect 64872 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64994 3800
rect 65038 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65160 3800
rect 65160 3760 65162 3800
rect 64870 3718 64994 3760
rect 65038 3718 65162 3760
rect 79990 3800 80114 3842
rect 80158 3800 80282 3842
rect 79990 3760 79992 3800
rect 79992 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80114 3800
rect 80158 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80280 3800
rect 80280 3760 80282 3800
rect 79990 3718 80114 3760
rect 80158 3718 80282 3760
rect 3150 3044 3274 3086
rect 3318 3044 3442 3086
rect 3150 3004 3152 3044
rect 3152 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3274 3044
rect 3318 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3440 3044
rect 3440 3004 3442 3044
rect 3150 2962 3274 3004
rect 3318 2962 3442 3004
rect 18270 3044 18394 3086
rect 18438 3044 18562 3086
rect 18270 3004 18272 3044
rect 18272 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18394 3044
rect 18438 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18560 3044
rect 18560 3004 18562 3044
rect 18270 2962 18394 3004
rect 18438 2962 18562 3004
rect 33390 3044 33514 3086
rect 33558 3044 33682 3086
rect 33390 3004 33392 3044
rect 33392 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33514 3044
rect 33558 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33680 3044
rect 33680 3004 33682 3044
rect 33390 2962 33514 3004
rect 33558 2962 33682 3004
rect 48510 3044 48634 3086
rect 48678 3044 48802 3086
rect 48510 3004 48512 3044
rect 48512 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48634 3044
rect 48678 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48800 3044
rect 48800 3004 48802 3044
rect 48510 2962 48634 3004
rect 48678 2962 48802 3004
rect 63630 3044 63754 3086
rect 63798 3044 63922 3086
rect 63630 3004 63632 3044
rect 63632 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63754 3044
rect 63798 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63920 3044
rect 63920 3004 63922 3044
rect 63630 2962 63754 3004
rect 63798 2962 63922 3004
rect 78750 3044 78874 3086
rect 78918 3044 79042 3086
rect 78750 3004 78752 3044
rect 78752 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78874 3044
rect 78918 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79040 3044
rect 79040 3004 79042 3044
rect 78750 2962 78874 3004
rect 78918 2962 79042 3004
rect 4390 2288 4514 2330
rect 4558 2288 4682 2330
rect 4390 2248 4392 2288
rect 4392 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4514 2288
rect 4558 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4680 2288
rect 4680 2248 4682 2288
rect 4390 2206 4514 2248
rect 4558 2206 4682 2248
rect 19510 2288 19634 2330
rect 19678 2288 19802 2330
rect 19510 2248 19512 2288
rect 19512 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19634 2288
rect 19678 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19800 2288
rect 19800 2248 19802 2288
rect 19510 2206 19634 2248
rect 19678 2206 19802 2248
rect 34630 2288 34754 2330
rect 34798 2288 34922 2330
rect 34630 2248 34632 2288
rect 34632 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34754 2288
rect 34798 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34920 2288
rect 34920 2248 34922 2288
rect 34630 2206 34754 2248
rect 34798 2206 34922 2248
rect 49750 2288 49874 2330
rect 49918 2288 50042 2330
rect 49750 2248 49752 2288
rect 49752 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49874 2288
rect 49918 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50040 2288
rect 50040 2248 50042 2288
rect 49750 2206 49874 2248
rect 49918 2206 50042 2248
rect 64870 2288 64994 2330
rect 65038 2288 65162 2330
rect 64870 2248 64872 2288
rect 64872 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64994 2288
rect 65038 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65160 2288
rect 65160 2248 65162 2288
rect 64870 2206 64994 2248
rect 65038 2206 65162 2248
rect 79990 2288 80114 2330
rect 80158 2288 80282 2330
rect 79990 2248 79992 2288
rect 79992 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80114 2288
rect 80158 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80280 2288
rect 80280 2248 80282 2288
rect 79990 2206 80114 2248
rect 80158 2206 80282 2248
rect 3150 1532 3274 1574
rect 3318 1532 3442 1574
rect 3150 1492 3152 1532
rect 3152 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3274 1532
rect 3318 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3440 1532
rect 3440 1492 3442 1532
rect 3150 1450 3274 1492
rect 3318 1450 3442 1492
rect 18270 1532 18394 1574
rect 18438 1532 18562 1574
rect 18270 1492 18272 1532
rect 18272 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18394 1532
rect 18438 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18560 1532
rect 18560 1492 18562 1532
rect 18270 1450 18394 1492
rect 18438 1450 18562 1492
rect 33390 1532 33514 1574
rect 33558 1532 33682 1574
rect 33390 1492 33392 1532
rect 33392 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33514 1532
rect 33558 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33680 1532
rect 33680 1492 33682 1532
rect 33390 1450 33514 1492
rect 33558 1450 33682 1492
rect 48510 1532 48634 1574
rect 48678 1532 48802 1574
rect 48510 1492 48512 1532
rect 48512 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48634 1532
rect 48678 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48800 1532
rect 48800 1492 48802 1532
rect 48510 1450 48634 1492
rect 48678 1450 48802 1492
rect 63630 1532 63754 1574
rect 63798 1532 63922 1574
rect 63630 1492 63632 1532
rect 63632 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63754 1532
rect 63798 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63920 1532
rect 63920 1492 63922 1532
rect 63630 1450 63754 1492
rect 63798 1450 63922 1492
rect 78750 1532 78874 1574
rect 78918 1532 79042 1574
rect 78750 1492 78752 1532
rect 78752 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78874 1532
rect 78918 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79040 1532
rect 79040 1492 79042 1532
rect 78750 1450 78874 1492
rect 78918 1450 79042 1492
rect 4390 776 4514 818
rect 4558 776 4682 818
rect 4390 736 4392 776
rect 4392 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4514 776
rect 4558 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4680 776
rect 4680 736 4682 776
rect 4390 694 4514 736
rect 4558 694 4682 736
rect 19510 776 19634 818
rect 19678 776 19802 818
rect 19510 736 19512 776
rect 19512 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19634 776
rect 19678 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19800 776
rect 19800 736 19802 776
rect 19510 694 19634 736
rect 19678 694 19802 736
rect 34630 776 34754 818
rect 34798 776 34922 818
rect 34630 736 34632 776
rect 34632 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34754 776
rect 34798 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34920 776
rect 34920 736 34922 776
rect 34630 694 34754 736
rect 34798 694 34922 736
rect 49750 776 49874 818
rect 49918 776 50042 818
rect 49750 736 49752 776
rect 49752 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49874 776
rect 49918 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50040 776
rect 50040 736 50042 776
rect 49750 694 49874 736
rect 49918 694 50042 736
rect 64870 776 64994 818
rect 65038 776 65162 818
rect 64870 736 64872 776
rect 64872 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64994 776
rect 65038 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65160 776
rect 65160 736 65162 776
rect 64870 694 64994 736
rect 65038 694 65162 736
rect 79990 776 80114 818
rect 80158 776 80282 818
rect 79990 736 79992 776
rect 79992 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80114 776
rect 80158 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80280 776
rect 80280 736 80282 776
rect 79990 694 80114 736
rect 80158 694 80282 736
<< metal6 >>
rect 4316 38618 4756 38682
rect 3076 37862 3516 38600
rect 3076 37738 3150 37862
rect 3274 37738 3318 37862
rect 3442 37738 3516 37862
rect 3076 36350 3516 37738
rect 3076 36226 3150 36350
rect 3274 36226 3318 36350
rect 3442 36226 3516 36350
rect 3076 34838 3516 36226
rect 3076 34714 3150 34838
rect 3274 34714 3318 34838
rect 3442 34714 3516 34838
rect 3076 33326 3516 34714
rect 3076 33202 3150 33326
rect 3274 33202 3318 33326
rect 3442 33202 3516 33326
rect 3076 31814 3516 33202
rect 3076 31690 3150 31814
rect 3274 31690 3318 31814
rect 3442 31690 3516 31814
rect 3076 30302 3516 31690
rect 3076 30178 3150 30302
rect 3274 30178 3318 30302
rect 3442 30178 3516 30302
rect 3076 28790 3516 30178
rect 3076 28666 3150 28790
rect 3274 28666 3318 28790
rect 3442 28666 3516 28790
rect 3076 27278 3516 28666
rect 3076 27154 3150 27278
rect 3274 27154 3318 27278
rect 3442 27154 3516 27278
rect 3076 25766 3516 27154
rect 3076 25642 3150 25766
rect 3274 25642 3318 25766
rect 3442 25642 3516 25766
rect 3076 24254 3516 25642
rect 3076 24130 3150 24254
rect 3274 24130 3318 24254
rect 3442 24130 3516 24254
rect 3076 22742 3516 24130
rect 3076 22618 3150 22742
rect 3274 22618 3318 22742
rect 3442 22618 3516 22742
rect 3076 21230 3516 22618
rect 3076 21106 3150 21230
rect 3274 21106 3318 21230
rect 3442 21106 3516 21230
rect 3076 19718 3516 21106
rect 3076 19594 3150 19718
rect 3274 19594 3318 19718
rect 3442 19594 3516 19718
rect 3076 18206 3516 19594
rect 3076 18082 3150 18206
rect 3274 18082 3318 18206
rect 3442 18082 3516 18206
rect 3076 16694 3516 18082
rect 3076 16570 3150 16694
rect 3274 16570 3318 16694
rect 3442 16570 3516 16694
rect 3076 15182 3516 16570
rect 3076 15058 3150 15182
rect 3274 15058 3318 15182
rect 3442 15058 3516 15182
rect 3076 13670 3516 15058
rect 3076 13546 3150 13670
rect 3274 13546 3318 13670
rect 3442 13546 3516 13670
rect 3076 12158 3516 13546
rect 3076 12034 3150 12158
rect 3274 12034 3318 12158
rect 3442 12034 3516 12158
rect 3076 10646 3516 12034
rect 3076 10522 3150 10646
rect 3274 10522 3318 10646
rect 3442 10522 3516 10646
rect 3076 9134 3516 10522
rect 3076 9010 3150 9134
rect 3274 9010 3318 9134
rect 3442 9010 3516 9134
rect 3076 7622 3516 9010
rect 3076 7498 3150 7622
rect 3274 7498 3318 7622
rect 3442 7498 3516 7622
rect 3076 6110 3516 7498
rect 3076 5986 3150 6110
rect 3274 5986 3318 6110
rect 3442 5986 3516 6110
rect 3076 4598 3516 5986
rect 3076 4474 3150 4598
rect 3274 4474 3318 4598
rect 3442 4474 3516 4598
rect 3076 3086 3516 4474
rect 3076 2962 3150 3086
rect 3274 2962 3318 3086
rect 3442 2962 3516 3086
rect 3076 1574 3516 2962
rect 3076 1450 3150 1574
rect 3274 1450 3318 1574
rect 3442 1450 3516 1574
rect 3076 712 3516 1450
rect 4316 38494 4390 38618
rect 4514 38494 4558 38618
rect 4682 38494 4756 38618
rect 19436 38618 19876 38682
rect 4316 37106 4756 38494
rect 4316 36982 4390 37106
rect 4514 36982 4558 37106
rect 4682 36982 4756 37106
rect 4316 35594 4756 36982
rect 4316 35470 4390 35594
rect 4514 35470 4558 35594
rect 4682 35470 4756 35594
rect 4316 34082 4756 35470
rect 4316 33958 4390 34082
rect 4514 33958 4558 34082
rect 4682 33958 4756 34082
rect 4316 32570 4756 33958
rect 4316 32446 4390 32570
rect 4514 32446 4558 32570
rect 4682 32446 4756 32570
rect 4316 31058 4756 32446
rect 4316 30934 4390 31058
rect 4514 30934 4558 31058
rect 4682 30934 4756 31058
rect 4316 29546 4756 30934
rect 4316 29422 4390 29546
rect 4514 29422 4558 29546
rect 4682 29422 4756 29546
rect 4316 28034 4756 29422
rect 4316 27910 4390 28034
rect 4514 27910 4558 28034
rect 4682 27910 4756 28034
rect 4316 26522 4756 27910
rect 4316 26398 4390 26522
rect 4514 26398 4558 26522
rect 4682 26398 4756 26522
rect 4316 25010 4756 26398
rect 4316 24886 4390 25010
rect 4514 24886 4558 25010
rect 4682 24886 4756 25010
rect 4316 23498 4756 24886
rect 4316 23374 4390 23498
rect 4514 23374 4558 23498
rect 4682 23374 4756 23498
rect 4316 21986 4756 23374
rect 4316 21862 4390 21986
rect 4514 21862 4558 21986
rect 4682 21862 4756 21986
rect 4316 20474 4756 21862
rect 4316 20350 4390 20474
rect 4514 20350 4558 20474
rect 4682 20350 4756 20474
rect 4316 18962 4756 20350
rect 4316 18838 4390 18962
rect 4514 18838 4558 18962
rect 4682 18838 4756 18962
rect 4316 17450 4756 18838
rect 4316 17326 4390 17450
rect 4514 17326 4558 17450
rect 4682 17326 4756 17450
rect 4316 15938 4756 17326
rect 4316 15814 4390 15938
rect 4514 15814 4558 15938
rect 4682 15814 4756 15938
rect 4316 14426 4756 15814
rect 4316 14302 4390 14426
rect 4514 14302 4558 14426
rect 4682 14302 4756 14426
rect 4316 12914 4756 14302
rect 4316 12790 4390 12914
rect 4514 12790 4558 12914
rect 4682 12790 4756 12914
rect 4316 11402 4756 12790
rect 4316 11278 4390 11402
rect 4514 11278 4558 11402
rect 4682 11278 4756 11402
rect 4316 9890 4756 11278
rect 4316 9766 4390 9890
rect 4514 9766 4558 9890
rect 4682 9766 4756 9890
rect 4316 8378 4756 9766
rect 4316 8254 4390 8378
rect 4514 8254 4558 8378
rect 4682 8254 4756 8378
rect 4316 6866 4756 8254
rect 4316 6742 4390 6866
rect 4514 6742 4558 6866
rect 4682 6742 4756 6866
rect 4316 5354 4756 6742
rect 4316 5230 4390 5354
rect 4514 5230 4558 5354
rect 4682 5230 4756 5354
rect 4316 3842 4756 5230
rect 4316 3718 4390 3842
rect 4514 3718 4558 3842
rect 4682 3718 4756 3842
rect 4316 2330 4756 3718
rect 4316 2206 4390 2330
rect 4514 2206 4558 2330
rect 4682 2206 4756 2330
rect 4316 818 4756 2206
rect 4316 694 4390 818
rect 4514 694 4558 818
rect 4682 694 4756 818
rect 18196 37862 18636 38600
rect 18196 37738 18270 37862
rect 18394 37738 18438 37862
rect 18562 37738 18636 37862
rect 18196 36350 18636 37738
rect 18196 36226 18270 36350
rect 18394 36226 18438 36350
rect 18562 36226 18636 36350
rect 18196 34838 18636 36226
rect 18196 34714 18270 34838
rect 18394 34714 18438 34838
rect 18562 34714 18636 34838
rect 18196 33326 18636 34714
rect 18196 33202 18270 33326
rect 18394 33202 18438 33326
rect 18562 33202 18636 33326
rect 18196 27622 18636 33202
rect 18196 27498 18270 27622
rect 18394 27498 18438 27622
rect 18562 27498 18636 27622
rect 18196 27454 18636 27498
rect 18196 27330 18270 27454
rect 18394 27330 18438 27454
rect 18562 27330 18636 27454
rect 18196 21622 18636 27330
rect 18196 21498 18270 21622
rect 18394 21498 18438 21622
rect 18562 21498 18636 21622
rect 18196 21454 18636 21498
rect 18196 21330 18270 21454
rect 18394 21330 18438 21454
rect 18562 21330 18636 21454
rect 18196 15622 18636 21330
rect 18196 15498 18270 15622
rect 18394 15498 18438 15622
rect 18562 15498 18636 15622
rect 18196 15454 18636 15498
rect 18196 15330 18270 15454
rect 18394 15330 18438 15454
rect 18562 15330 18636 15454
rect 18196 9622 18636 15330
rect 18196 9498 18270 9622
rect 18394 9498 18438 9622
rect 18562 9498 18636 9622
rect 18196 9454 18636 9498
rect 18196 9330 18270 9454
rect 18394 9330 18438 9454
rect 18562 9330 18636 9454
rect 18196 3086 18636 9330
rect 18196 2962 18270 3086
rect 18394 2962 18438 3086
rect 18562 2962 18636 3086
rect 18196 1574 18636 2962
rect 18196 1450 18270 1574
rect 18394 1450 18438 1574
rect 18562 1450 18636 1574
rect 18196 712 18636 1450
rect 19436 38494 19510 38618
rect 19634 38494 19678 38618
rect 19802 38494 19876 38618
rect 34556 38618 34996 38682
rect 19436 37106 19876 38494
rect 19436 36982 19510 37106
rect 19634 36982 19678 37106
rect 19802 36982 19876 37106
rect 19436 35594 19876 36982
rect 19436 35470 19510 35594
rect 19634 35470 19678 35594
rect 19802 35470 19876 35594
rect 19436 34082 19876 35470
rect 19436 33958 19510 34082
rect 19634 33958 19678 34082
rect 19802 33958 19876 34082
rect 19436 32570 19876 33958
rect 19436 32446 19510 32570
rect 19634 32446 19678 32570
rect 19802 32446 19876 32570
rect 19436 22862 19876 32446
rect 19436 22738 19510 22862
rect 19634 22738 19678 22862
rect 19802 22738 19876 22862
rect 19436 22694 19876 22738
rect 19436 22570 19510 22694
rect 19634 22570 19678 22694
rect 19802 22570 19876 22694
rect 19436 16862 19876 22570
rect 19436 16738 19510 16862
rect 19634 16738 19678 16862
rect 19802 16738 19876 16862
rect 19436 16694 19876 16738
rect 19436 16570 19510 16694
rect 19634 16570 19678 16694
rect 19802 16570 19876 16694
rect 19436 10862 19876 16570
rect 19436 10738 19510 10862
rect 19634 10738 19678 10862
rect 19802 10738 19876 10862
rect 19436 10694 19876 10738
rect 19436 10570 19510 10694
rect 19634 10570 19678 10694
rect 19802 10570 19876 10694
rect 19436 3842 19876 10570
rect 19436 3718 19510 3842
rect 19634 3718 19678 3842
rect 19802 3718 19876 3842
rect 19436 2330 19876 3718
rect 19436 2206 19510 2330
rect 19634 2206 19678 2330
rect 19802 2206 19876 2330
rect 19436 818 19876 2206
rect 4316 630 4756 694
rect 19436 694 19510 818
rect 19634 694 19678 818
rect 19802 694 19876 818
rect 33316 37862 33756 38600
rect 33316 37738 33390 37862
rect 33514 37738 33558 37862
rect 33682 37738 33756 37862
rect 33316 36350 33756 37738
rect 33316 36226 33390 36350
rect 33514 36226 33558 36350
rect 33682 36226 33756 36350
rect 33316 34838 33756 36226
rect 33316 34714 33390 34838
rect 33514 34714 33558 34838
rect 33682 34714 33756 34838
rect 33316 33326 33756 34714
rect 33316 33202 33390 33326
rect 33514 33202 33558 33326
rect 33682 33202 33756 33326
rect 33316 27622 33756 33202
rect 33316 27498 33390 27622
rect 33514 27498 33558 27622
rect 33682 27498 33756 27622
rect 33316 27454 33756 27498
rect 33316 27330 33390 27454
rect 33514 27330 33558 27454
rect 33682 27330 33756 27454
rect 33316 21622 33756 27330
rect 33316 21498 33390 21622
rect 33514 21498 33558 21622
rect 33682 21498 33756 21622
rect 33316 21454 33756 21498
rect 33316 21330 33390 21454
rect 33514 21330 33558 21454
rect 33682 21330 33756 21454
rect 33316 15622 33756 21330
rect 33316 15498 33390 15622
rect 33514 15498 33558 15622
rect 33682 15498 33756 15622
rect 33316 15454 33756 15498
rect 33316 15330 33390 15454
rect 33514 15330 33558 15454
rect 33682 15330 33756 15454
rect 33316 9622 33756 15330
rect 33316 9498 33390 9622
rect 33514 9498 33558 9622
rect 33682 9498 33756 9622
rect 33316 9454 33756 9498
rect 33316 9330 33390 9454
rect 33514 9330 33558 9454
rect 33682 9330 33756 9454
rect 33316 3086 33756 9330
rect 33316 2962 33390 3086
rect 33514 2962 33558 3086
rect 33682 2962 33756 3086
rect 33316 1574 33756 2962
rect 33316 1450 33390 1574
rect 33514 1450 33558 1574
rect 33682 1450 33756 1574
rect 33316 712 33756 1450
rect 34556 38494 34630 38618
rect 34754 38494 34798 38618
rect 34922 38494 34996 38618
rect 49676 38618 50116 38682
rect 34556 37106 34996 38494
rect 34556 36982 34630 37106
rect 34754 36982 34798 37106
rect 34922 36982 34996 37106
rect 34556 35594 34996 36982
rect 34556 35470 34630 35594
rect 34754 35470 34798 35594
rect 34922 35470 34996 35594
rect 34556 34082 34996 35470
rect 34556 33958 34630 34082
rect 34754 33958 34798 34082
rect 34922 33958 34996 34082
rect 34556 32570 34996 33958
rect 34556 32446 34630 32570
rect 34754 32446 34798 32570
rect 34922 32446 34996 32570
rect 34556 22862 34996 32446
rect 34556 22738 34630 22862
rect 34754 22738 34798 22862
rect 34922 22738 34996 22862
rect 34556 22694 34996 22738
rect 34556 22570 34630 22694
rect 34754 22570 34798 22694
rect 34922 22570 34996 22694
rect 34556 16862 34996 22570
rect 34556 16738 34630 16862
rect 34754 16738 34798 16862
rect 34922 16738 34996 16862
rect 34556 16694 34996 16738
rect 34556 16570 34630 16694
rect 34754 16570 34798 16694
rect 34922 16570 34996 16694
rect 34556 10862 34996 16570
rect 34556 10738 34630 10862
rect 34754 10738 34798 10862
rect 34922 10738 34996 10862
rect 34556 10694 34996 10738
rect 34556 10570 34630 10694
rect 34754 10570 34798 10694
rect 34922 10570 34996 10694
rect 34556 3842 34996 10570
rect 34556 3718 34630 3842
rect 34754 3718 34798 3842
rect 34922 3718 34996 3842
rect 34556 2330 34996 3718
rect 34556 2206 34630 2330
rect 34754 2206 34798 2330
rect 34922 2206 34996 2330
rect 34556 818 34996 2206
rect 19436 630 19876 694
rect 34556 694 34630 818
rect 34754 694 34798 818
rect 34922 694 34996 818
rect 48436 37862 48876 38600
rect 48436 37738 48510 37862
rect 48634 37738 48678 37862
rect 48802 37738 48876 37862
rect 48436 36350 48876 37738
rect 48436 36226 48510 36350
rect 48634 36226 48678 36350
rect 48802 36226 48876 36350
rect 48436 34838 48876 36226
rect 48436 34714 48510 34838
rect 48634 34714 48678 34838
rect 48802 34714 48876 34838
rect 48436 33326 48876 34714
rect 48436 33202 48510 33326
rect 48634 33202 48678 33326
rect 48802 33202 48876 33326
rect 48436 27622 48876 33202
rect 48436 27498 48510 27622
rect 48634 27498 48678 27622
rect 48802 27498 48876 27622
rect 48436 27454 48876 27498
rect 48436 27330 48510 27454
rect 48634 27330 48678 27454
rect 48802 27330 48876 27454
rect 48436 21622 48876 27330
rect 48436 21498 48510 21622
rect 48634 21498 48678 21622
rect 48802 21498 48876 21622
rect 48436 21454 48876 21498
rect 48436 21330 48510 21454
rect 48634 21330 48678 21454
rect 48802 21330 48876 21454
rect 48436 15622 48876 21330
rect 48436 15498 48510 15622
rect 48634 15498 48678 15622
rect 48802 15498 48876 15622
rect 48436 15454 48876 15498
rect 48436 15330 48510 15454
rect 48634 15330 48678 15454
rect 48802 15330 48876 15454
rect 48436 9622 48876 15330
rect 48436 9498 48510 9622
rect 48634 9498 48678 9622
rect 48802 9498 48876 9622
rect 48436 9454 48876 9498
rect 48436 9330 48510 9454
rect 48634 9330 48678 9454
rect 48802 9330 48876 9454
rect 48436 3086 48876 9330
rect 48436 2962 48510 3086
rect 48634 2962 48678 3086
rect 48802 2962 48876 3086
rect 48436 1574 48876 2962
rect 48436 1450 48510 1574
rect 48634 1450 48678 1574
rect 48802 1450 48876 1574
rect 48436 712 48876 1450
rect 49676 38494 49750 38618
rect 49874 38494 49918 38618
rect 50042 38494 50116 38618
rect 64796 38618 65236 38682
rect 49676 37106 50116 38494
rect 49676 36982 49750 37106
rect 49874 36982 49918 37106
rect 50042 36982 50116 37106
rect 49676 35594 50116 36982
rect 49676 35470 49750 35594
rect 49874 35470 49918 35594
rect 50042 35470 50116 35594
rect 49676 34082 50116 35470
rect 49676 33958 49750 34082
rect 49874 33958 49918 34082
rect 50042 33958 50116 34082
rect 49676 32570 50116 33958
rect 49676 32446 49750 32570
rect 49874 32446 49918 32570
rect 50042 32446 50116 32570
rect 49676 22862 50116 32446
rect 49676 22738 49750 22862
rect 49874 22738 49918 22862
rect 50042 22738 50116 22862
rect 49676 22694 50116 22738
rect 49676 22570 49750 22694
rect 49874 22570 49918 22694
rect 50042 22570 50116 22694
rect 49676 16862 50116 22570
rect 49676 16738 49750 16862
rect 49874 16738 49918 16862
rect 50042 16738 50116 16862
rect 49676 16694 50116 16738
rect 49676 16570 49750 16694
rect 49874 16570 49918 16694
rect 50042 16570 50116 16694
rect 49676 10862 50116 16570
rect 49676 10738 49750 10862
rect 49874 10738 49918 10862
rect 50042 10738 50116 10862
rect 49676 10694 50116 10738
rect 49676 10570 49750 10694
rect 49874 10570 49918 10694
rect 50042 10570 50116 10694
rect 49676 3842 50116 10570
rect 49676 3718 49750 3842
rect 49874 3718 49918 3842
rect 50042 3718 50116 3842
rect 49676 2330 50116 3718
rect 49676 2206 49750 2330
rect 49874 2206 49918 2330
rect 50042 2206 50116 2330
rect 49676 818 50116 2206
rect 34556 630 34996 694
rect 49676 694 49750 818
rect 49874 694 49918 818
rect 50042 694 50116 818
rect 63556 37862 63996 38600
rect 63556 37738 63630 37862
rect 63754 37738 63798 37862
rect 63922 37738 63996 37862
rect 63556 36350 63996 37738
rect 63556 36226 63630 36350
rect 63754 36226 63798 36350
rect 63922 36226 63996 36350
rect 63556 34838 63996 36226
rect 63556 34714 63630 34838
rect 63754 34714 63798 34838
rect 63922 34714 63996 34838
rect 63556 33326 63996 34714
rect 63556 33202 63630 33326
rect 63754 33202 63798 33326
rect 63922 33202 63996 33326
rect 63556 27622 63996 33202
rect 63556 27498 63630 27622
rect 63754 27498 63798 27622
rect 63922 27498 63996 27622
rect 63556 27454 63996 27498
rect 63556 27330 63630 27454
rect 63754 27330 63798 27454
rect 63922 27330 63996 27454
rect 63556 21622 63996 27330
rect 63556 21498 63630 21622
rect 63754 21498 63798 21622
rect 63922 21498 63996 21622
rect 63556 21454 63996 21498
rect 63556 21330 63630 21454
rect 63754 21330 63798 21454
rect 63922 21330 63996 21454
rect 63556 15622 63996 21330
rect 63556 15498 63630 15622
rect 63754 15498 63798 15622
rect 63922 15498 63996 15622
rect 63556 15454 63996 15498
rect 63556 15330 63630 15454
rect 63754 15330 63798 15454
rect 63922 15330 63996 15454
rect 63556 9622 63996 15330
rect 63556 9498 63630 9622
rect 63754 9498 63798 9622
rect 63922 9498 63996 9622
rect 63556 9454 63996 9498
rect 63556 9330 63630 9454
rect 63754 9330 63798 9454
rect 63922 9330 63996 9454
rect 63556 3086 63996 9330
rect 63556 2962 63630 3086
rect 63754 2962 63798 3086
rect 63922 2962 63996 3086
rect 63556 1574 63996 2962
rect 63556 1450 63630 1574
rect 63754 1450 63798 1574
rect 63922 1450 63996 1574
rect 63556 712 63996 1450
rect 64796 38494 64870 38618
rect 64994 38494 65038 38618
rect 65162 38494 65236 38618
rect 79916 38618 80356 38682
rect 64796 37106 65236 38494
rect 64796 36982 64870 37106
rect 64994 36982 65038 37106
rect 65162 36982 65236 37106
rect 64796 35594 65236 36982
rect 64796 35470 64870 35594
rect 64994 35470 65038 35594
rect 65162 35470 65236 35594
rect 64796 34082 65236 35470
rect 64796 33958 64870 34082
rect 64994 33958 65038 34082
rect 65162 33958 65236 34082
rect 64796 32570 65236 33958
rect 64796 32446 64870 32570
rect 64994 32446 65038 32570
rect 65162 32446 65236 32570
rect 64796 22862 65236 32446
rect 78676 37862 79116 38600
rect 78676 37738 78750 37862
rect 78874 37738 78918 37862
rect 79042 37738 79116 37862
rect 78676 36350 79116 37738
rect 78676 36226 78750 36350
rect 78874 36226 78918 36350
rect 79042 36226 79116 36350
rect 78676 34838 79116 36226
rect 78676 34714 78750 34838
rect 78874 34714 78918 34838
rect 79042 34714 79116 34838
rect 78676 33326 79116 34714
rect 78676 33202 78750 33326
rect 78874 33202 78918 33326
rect 79042 33202 79116 33326
rect 78676 31814 79116 33202
rect 78676 31690 78750 31814
rect 78874 31690 78918 31814
rect 79042 31690 79116 31814
rect 78676 30302 79116 31690
rect 78676 30178 78750 30302
rect 78874 30178 78918 30302
rect 79042 30178 79116 30302
rect 64796 22738 64870 22862
rect 64994 22738 65038 22862
rect 65162 22738 65236 22862
rect 64796 22694 65236 22738
rect 64796 22570 64870 22694
rect 64994 22570 65038 22694
rect 65162 22570 65236 22694
rect 64796 16862 65236 22570
rect 64796 16738 64870 16862
rect 64994 16738 65038 16862
rect 65162 16738 65236 16862
rect 64796 16694 65236 16738
rect 64796 16570 64870 16694
rect 64994 16570 65038 16694
rect 65162 16570 65236 16694
rect 64796 10862 65236 16570
rect 64796 10738 64870 10862
rect 64994 10738 65038 10862
rect 65162 10738 65236 10862
rect 64796 10694 65236 10738
rect 64796 10570 64870 10694
rect 64994 10570 65038 10694
rect 65162 10570 65236 10694
rect 64796 3842 65236 10570
rect 66284 28790 66612 28892
rect 66284 28666 66386 28790
rect 66510 28666 66612 28790
rect 78676 28790 79116 30178
rect 66284 5102 66612 28666
rect 66284 4978 66386 5102
rect 66510 4978 66612 5102
rect 66284 4876 66612 4978
rect 67196 28622 67524 28724
rect 67196 28498 67298 28622
rect 67422 28498 67524 28622
rect 67196 4514 67524 28498
rect 67196 4390 67298 4514
rect 67422 4390 67524 4514
rect 67196 4288 67524 4390
rect 78676 28666 78750 28790
rect 78874 28666 78918 28790
rect 79042 28666 79116 28790
rect 78676 27278 79116 28666
rect 78676 27154 78750 27278
rect 78874 27154 78918 27278
rect 79042 27154 79116 27278
rect 78676 25766 79116 27154
rect 78676 25642 78750 25766
rect 78874 25642 78918 25766
rect 79042 25642 79116 25766
rect 78676 24254 79116 25642
rect 78676 24130 78750 24254
rect 78874 24130 78918 24254
rect 79042 24130 79116 24254
rect 78676 22742 79116 24130
rect 78676 22618 78750 22742
rect 78874 22618 78918 22742
rect 79042 22618 79116 22742
rect 78676 21230 79116 22618
rect 78676 21106 78750 21230
rect 78874 21106 78918 21230
rect 79042 21106 79116 21230
rect 78676 19718 79116 21106
rect 78676 19594 78750 19718
rect 78874 19594 78918 19718
rect 79042 19594 79116 19718
rect 78676 18206 79116 19594
rect 78676 18082 78750 18206
rect 78874 18082 78918 18206
rect 79042 18082 79116 18206
rect 78676 16694 79116 18082
rect 78676 16570 78750 16694
rect 78874 16570 78918 16694
rect 79042 16570 79116 16694
rect 78676 15182 79116 16570
rect 78676 15058 78750 15182
rect 78874 15058 78918 15182
rect 79042 15058 79116 15182
rect 78676 13670 79116 15058
rect 78676 13546 78750 13670
rect 78874 13546 78918 13670
rect 79042 13546 79116 13670
rect 78676 12158 79116 13546
rect 78676 12034 78750 12158
rect 78874 12034 78918 12158
rect 79042 12034 79116 12158
rect 78676 10646 79116 12034
rect 78676 10522 78750 10646
rect 78874 10522 78918 10646
rect 79042 10522 79116 10646
rect 78676 9134 79116 10522
rect 78676 9010 78750 9134
rect 78874 9010 78918 9134
rect 79042 9010 79116 9134
rect 78676 7622 79116 9010
rect 78676 7498 78750 7622
rect 78874 7498 78918 7622
rect 79042 7498 79116 7622
rect 78676 6110 79116 7498
rect 78676 5986 78750 6110
rect 78874 5986 78918 6110
rect 79042 5986 79116 6110
rect 78676 4598 79116 5986
rect 78676 4474 78750 4598
rect 78874 4474 78918 4598
rect 79042 4474 79116 4598
rect 64796 3718 64870 3842
rect 64994 3718 65038 3842
rect 65162 3718 65236 3842
rect 64796 2330 65236 3718
rect 64796 2206 64870 2330
rect 64994 2206 65038 2330
rect 65162 2206 65236 2330
rect 64796 818 65236 2206
rect 49676 630 50116 694
rect 64796 694 64870 818
rect 64994 694 65038 818
rect 65162 694 65236 818
rect 78676 3086 79116 4474
rect 78676 2962 78750 3086
rect 78874 2962 78918 3086
rect 79042 2962 79116 3086
rect 78676 1574 79116 2962
rect 78676 1450 78750 1574
rect 78874 1450 78918 1574
rect 79042 1450 79116 1574
rect 78676 712 79116 1450
rect 79916 38494 79990 38618
rect 80114 38494 80158 38618
rect 80282 38494 80356 38618
rect 79916 37106 80356 38494
rect 79916 36982 79990 37106
rect 80114 36982 80158 37106
rect 80282 36982 80356 37106
rect 79916 35594 80356 36982
rect 79916 35470 79990 35594
rect 80114 35470 80158 35594
rect 80282 35470 80356 35594
rect 79916 34082 80356 35470
rect 79916 33958 79990 34082
rect 80114 33958 80158 34082
rect 80282 33958 80356 34082
rect 79916 32570 80356 33958
rect 79916 32446 79990 32570
rect 80114 32446 80158 32570
rect 80282 32446 80356 32570
rect 79916 31058 80356 32446
rect 79916 30934 79990 31058
rect 80114 30934 80158 31058
rect 80282 30934 80356 31058
rect 79916 29546 80356 30934
rect 79916 29422 79990 29546
rect 80114 29422 80158 29546
rect 80282 29422 80356 29546
rect 79916 28034 80356 29422
rect 79916 27910 79990 28034
rect 80114 27910 80158 28034
rect 80282 27910 80356 28034
rect 79916 26522 80356 27910
rect 79916 26398 79990 26522
rect 80114 26398 80158 26522
rect 80282 26398 80356 26522
rect 79916 25010 80356 26398
rect 79916 24886 79990 25010
rect 80114 24886 80158 25010
rect 80282 24886 80356 25010
rect 79916 23498 80356 24886
rect 79916 23374 79990 23498
rect 80114 23374 80158 23498
rect 80282 23374 80356 23498
rect 79916 21986 80356 23374
rect 79916 21862 79990 21986
rect 80114 21862 80158 21986
rect 80282 21862 80356 21986
rect 79916 20474 80356 21862
rect 79916 20350 79990 20474
rect 80114 20350 80158 20474
rect 80282 20350 80356 20474
rect 79916 18962 80356 20350
rect 79916 18838 79990 18962
rect 80114 18838 80158 18962
rect 80282 18838 80356 18962
rect 79916 17450 80356 18838
rect 79916 17326 79990 17450
rect 80114 17326 80158 17450
rect 80282 17326 80356 17450
rect 79916 15938 80356 17326
rect 79916 15814 79990 15938
rect 80114 15814 80158 15938
rect 80282 15814 80356 15938
rect 79916 14426 80356 15814
rect 79916 14302 79990 14426
rect 80114 14302 80158 14426
rect 80282 14302 80356 14426
rect 79916 12914 80356 14302
rect 79916 12790 79990 12914
rect 80114 12790 80158 12914
rect 80282 12790 80356 12914
rect 79916 11402 80356 12790
rect 79916 11278 79990 11402
rect 80114 11278 80158 11402
rect 80282 11278 80356 11402
rect 79916 9890 80356 11278
rect 79916 9766 79990 9890
rect 80114 9766 80158 9890
rect 80282 9766 80356 9890
rect 79916 8378 80356 9766
rect 79916 8254 79990 8378
rect 80114 8254 80158 8378
rect 80282 8254 80356 8378
rect 79916 6866 80356 8254
rect 79916 6742 79990 6866
rect 80114 6742 80158 6866
rect 80282 6742 80356 6866
rect 79916 5354 80356 6742
rect 79916 5230 79990 5354
rect 80114 5230 80158 5354
rect 80282 5230 80356 5354
rect 79916 3842 80356 5230
rect 79916 3718 79990 3842
rect 80114 3718 80158 3842
rect 80282 3718 80356 3842
rect 79916 2330 80356 3718
rect 79916 2206 79990 2330
rect 80114 2206 80158 2330
rect 80282 2206 80356 2330
rect 79916 818 80356 2206
rect 64796 630 65236 694
rect 79916 694 79990 818
rect 80114 694 80158 818
rect 80282 694 80356 818
rect 93796 33822 94236 38600
rect 93796 33698 93870 33822
rect 93994 33698 94038 33822
rect 94162 33698 94236 33822
rect 93796 33654 94236 33698
rect 93796 33530 93870 33654
rect 93994 33530 94038 33654
rect 94162 33530 94236 33654
rect 93796 27822 94236 33530
rect 93796 27698 93870 27822
rect 93994 27698 94038 27822
rect 94162 27698 94236 27822
rect 93796 27654 94236 27698
rect 93796 27530 93870 27654
rect 93994 27530 94038 27654
rect 94162 27530 94236 27654
rect 93796 21230 94236 27530
rect 93796 21106 93870 21230
rect 93994 21106 94038 21230
rect 94162 21106 94236 21230
rect 93796 19718 94236 21106
rect 93796 19594 93870 19718
rect 93994 19594 94038 19718
rect 94162 19594 94236 19718
rect 93796 10622 94236 19594
rect 93796 10498 93870 10622
rect 93994 10498 94038 10622
rect 94162 10498 94236 10622
rect 93796 10454 94236 10498
rect 93796 10330 93870 10454
rect 93994 10330 94038 10454
rect 94162 10330 94236 10454
rect 93796 4622 94236 10330
rect 93796 4498 93870 4622
rect 93994 4498 94038 4622
rect 94162 4498 94236 4622
rect 93796 4454 94236 4498
rect 93796 4330 93870 4454
rect 93994 4330 94038 4454
rect 94162 4330 94236 4454
rect 93796 712 94236 4330
rect 95036 29062 95476 38600
rect 95036 28938 95110 29062
rect 95234 28938 95278 29062
rect 95402 28938 95476 29062
rect 95036 28894 95476 28938
rect 95036 28770 95110 28894
rect 95234 28770 95278 28894
rect 95402 28770 95476 28894
rect 95036 21986 95476 28770
rect 95036 21862 95110 21986
rect 95234 21862 95278 21986
rect 95402 21862 95476 21986
rect 95036 20474 95476 21862
rect 95036 20350 95110 20474
rect 95234 20350 95278 20474
rect 95402 20350 95476 20474
rect 95036 11862 95476 20350
rect 95036 11738 95110 11862
rect 95234 11738 95278 11862
rect 95402 11738 95476 11862
rect 95036 11694 95476 11738
rect 95036 11570 95110 11694
rect 95234 11570 95278 11694
rect 95402 11570 95476 11694
rect 95036 5862 95476 11570
rect 95036 5738 95110 5862
rect 95234 5738 95278 5862
rect 95402 5738 95476 5862
rect 95036 5694 95476 5738
rect 95036 5570 95110 5694
rect 95234 5570 95278 5694
rect 95402 5570 95476 5694
rect 95036 712 95476 5570
rect 79916 630 80356 694
use sg13g2_inv_1  _116_
timestamp 1676382929
transform -1 0 4704 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _117_
timestamp 1676382929
transform -1 0 4512 0 -1 24948
box -48 -56 336 834
use sg13g2_nor2b_1  _118_
timestamp 1685181386
transform -1 0 1248 0 -1 12852
box -54 -56 528 834
use sg13g2_and2_1  _119_
timestamp 1676901763
transform -1 0 1824 0 1 8316
box -48 -56 528 834
use sg13g2_and2_1  _120_
timestamp 1676901763
transform -1 0 1824 0 -1 11340
box -48 -56 528 834
use sg13g2_and2_1  _121_
timestamp 1676901763
transform -1 0 1440 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2_1  _122_
timestamp 1676627187
transform 1 0 1440 0 1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  _123_
timestamp 1685173987
transform 1 0 33888 0 -1 3780
box -48 -56 624 834
use sg13g2_inv_1  _124_
timestamp 1676382929
transform -1 0 1536 0 1 6804
box -48 -56 336 834
use sg13g2_a22oi_1  _125_
timestamp 1685173987
transform 1 0 30720 0 -1 3780
box -48 -56 624 834
use sg13g2_inv_1  _126_
timestamp 1676382929
transform -1 0 1824 0 1 6804
box -48 -56 336 834
use sg13g2_a22oi_1  _127_
timestamp 1685173987
transform -1 0 38304 0 -1 3780
box -48 -56 624 834
use sg13g2_inv_1  _128_
timestamp 1676382929
transform -1 0 2112 0 1 6804
box -48 -56 336 834
use sg13g2_a22oi_1  _129_
timestamp 1685173987
transform 1 0 36576 0 -1 3780
box -48 -56 624 834
use sg13g2_inv_1  _130_
timestamp 1676382929
transform -1 0 2112 0 1 12852
box -48 -56 336 834
use sg13g2_nand3b_1  _131_
timestamp 1676573470
transform 1 0 1248 0 -1 15876
box -48 -56 720 834
use sg13g2_a22oi_1  _132_
timestamp 1685173987
transform 1 0 37152 0 -1 3780
box -48 -56 624 834
use sg13g2_nand2_1  _133_
timestamp 1676557249
transform -1 0 2304 0 -1 15876
box -48 -56 432 834
use sg13g2_nor2b_1  _134_
timestamp 1685181386
transform 1 0 768 0 1 23436
box -54 -56 528 834
use sg13g2_nand2b_1  _135_
timestamp 1676567195
transform 1 0 1920 0 1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _136_
timestamp 1676627187
transform 1 0 4608 0 -1 26460
box -48 -56 432 834
use sg13g2_nor2b_1  _137_
timestamp 1685181386
transform 1 0 2304 0 1 26460
box -54 -56 528 834
use sg13g2_and2_1  _138_
timestamp 1676901763
transform 1 0 3744 0 -1 29484
box -48 -56 528 834
use sg13g2_nand4_1  _139_
timestamp 1685201930
transform -1 0 3744 0 -1 26460
box -48 -56 624 834
use sg13g2_inv_1  _140_
timestamp 1676382929
transform -1 0 2304 0 -1 24948
box -48 -56 336 834
use sg13g2_a21oi_1  _141_
timestamp 1683973020
transform 1 0 1632 0 1 24948
box -48 -56 528 834
use sg13g2_a21oi_1  _142_
timestamp 1683973020
transform -1 0 1824 0 1 26460
box -48 -56 528 834
use sg13g2_and2_1  _143_
timestamp 1676901763
transform 1 0 2688 0 -1 27972
box -48 -56 528 834
use sg13g2_and3_1  _144_
timestamp 1676971669
transform -1 0 2400 0 -1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _145_
timestamp 1683973020
transform 1 0 1824 0 -1 29484
box -48 -56 528 834
use sg13g2_nor2_1  _146_
timestamp 1676627187
transform -1 0 1824 0 -1 29484
box -48 -56 432 834
use sg13g2_nand4_1  _147_
timestamp 1685201930
transform -1 0 3168 0 -1 29484
box -48 -56 624 834
use sg13g2_o21ai_1  _148_
timestamp 1685175443
transform -1 0 2784 0 1 29484
box -48 -56 538 834
use sg13g2_inv_1  _149_
timestamp 1676382929
transform -1 0 2304 0 1 29484
box -48 -56 336 834
use sg13g2_and4_1  _150_
timestamp 1676985977
transform 1 0 3264 0 1 27972
box -48 -56 816 834
use sg13g2_a21oi_1  _151_
timestamp 1683973020
transform -1 0 3744 0 -1 29484
box -48 -56 528 834
use sg13g2_nand3_1  _152_
timestamp 1683988354
transform 1 0 3936 0 1 26460
box -48 -56 528 834
use sg13g2_and4_1  _153_
timestamp 1676985977
transform 1 0 3168 0 1 26460
box -48 -56 816 834
use sg13g2_nor2_1  _154_
timestamp 1676627187
transform -1 0 4416 0 1 27972
box -48 -56 432 834
use sg13g2_nor2_1  _155_
timestamp 1676627187
transform 1 0 4416 0 1 26460
box -48 -56 432 834
use sg13g2_nor3_1  _156_
timestamp 1676639442
transform -1 0 4224 0 -1 26460
box -48 -56 528 834
use sg13g2_nor2_1  _157_
timestamp 1676627187
transform -1 0 4608 0 -1 26460
box -48 -56 432 834
use sg13g2_nor2_1  _158_
timestamp 1676627187
transform 1 0 3840 0 -1 24948
box -48 -56 432 834
use sg13g2_xor2_1  _159_
timestamp 1677577977
transform -1 0 3840 0 -1 24948
box -48 -56 816 834
use sg13g2_mux2_1  _160_
timestamp 1677247768
transform 1 0 1056 0 1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  _161_
timestamp 1677247768
transform -1 0 28032 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _162_
timestamp 1677247768
transform -1 0 29856 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _163_
timestamp 1677247768
transform 1 0 30048 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _164_
timestamp 1677247768
transform 1 0 33600 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _165_
timestamp 1677247768
transform 1 0 40416 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _166_
timestamp 1677247768
transform 1 0 49152 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _167_
timestamp 1677247768
transform 1 0 51360 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _168_
timestamp 1677247768
transform -1 0 48096 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _169_
timestamp 1677247768
transform -1 0 46176 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _170_
timestamp 1677247768
transform -1 0 39072 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _171_
timestamp 1677247768
transform -1 0 33216 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _172_
timestamp 1677247768
transform 1 0 33600 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _173_
timestamp 1677247768
transform -1 0 33888 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _174_
timestamp 1677247768
transform 1 0 34464 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _175_
timestamp 1677247768
transform 1 0 45888 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _176_
timestamp 1677247768
transform 1 0 48480 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _177_
timestamp 1677247768
transform 1 0 51648 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _178_
timestamp 1677247768
transform 1 0 54432 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _179_
timestamp 1677247768
transform 1 0 51936 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _180_
timestamp 1677247768
transform 1 0 49440 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _181_
timestamp 1677247768
transform 1 0 46752 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _182_
timestamp 1677247768
transform 1 0 44256 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _183_
timestamp 1677247768
transform -1 0 39840 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _184_
timestamp 1677247768
transform -1 0 38496 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _185_
timestamp 1677247768
transform -1 0 36288 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _186_
timestamp 1677247768
transform 1 0 31104 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _187_
timestamp 1677247768
transform 1 0 29280 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _188_
timestamp 1677247768
transform 1 0 28224 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _189_
timestamp 1677247768
transform 1 0 26688 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _190_
timestamp 1677247768
transform 1 0 19488 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _191_
timestamp 1677247768
transform -1 0 20928 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _192_
timestamp 1677247768
transform 1 0 21600 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _193_
timestamp 1677247768
transform 1 0 21984 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _194_
timestamp 1677247768
transform 1 0 22944 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _195_
timestamp 1677247768
transform 1 0 24960 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _196_
timestamp 1677247768
transform 1 0 39456 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _197_
timestamp 1677247768
transform 1 0 41088 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _198_
timestamp 1677247768
transform 1 0 42240 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _199_
timestamp 1677247768
transform -1 0 5088 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _200_
timestamp 1677247768
transform -1 0 4800 0 1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  _201_
timestamp 1677247768
transform -1 0 5184 0 1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  _202_
timestamp 1677247768
transform 1 0 8736 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _203_
timestamp 1677247768
transform 1 0 13632 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _204_
timestamp 1677247768
transform 1 0 16800 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _205_
timestamp 1677247768
transform -1 0 16224 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _206_
timestamp 1677247768
transform -1 0 4896 0 -1 21924
box -48 -56 1008 834
use sg13g2_mux2_1  _207_
timestamp 1677247768
transform -1 0 4416 0 1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _208_
timestamp 1677247768
transform 1 0 1824 0 1 8316
box -48 -56 1008 834
use sg13g2_mux2_1  _209_
timestamp 1677247768
transform -1 0 2400 0 -1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  _210_
timestamp 1677247768
transform -1 0 2208 0 1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  _211_
timestamp 1677247768
transform -1 0 2208 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _212_
timestamp 1677247768
transform -1 0 2496 0 1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _213_
timestamp 1677247768
transform -1 0 2496 0 1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  _214_
timestamp 1677247768
transform -1 0 3360 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  _215_
timestamp 1677247768
transform -1 0 5856 0 1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  _216_
timestamp 1677247768
transform 1 0 17088 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _217_
timestamp 1677247768
transform 1 0 20544 0 -1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _218_
timestamp 1677247768
transform 1 0 21888 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _219_
timestamp 1677247768
transform -1 0 17760 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _220_
timestamp 1677247768
transform 1 0 12768 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _221_
timestamp 1677247768
transform -1 0 5088 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _222_
timestamp 1677247768
transform -1 0 4896 0 -1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  _223_
timestamp 1677247768
transform -1 0 4608 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  _224_
timestamp 1677247768
transform -1 0 4800 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _225_
timestamp 1677247768
transform -1 0 4512 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _226_
timestamp 1677247768
transform 1 0 75744 0 1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _227_
timestamp 1677247768
transform 1 0 78912 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _228_
timestamp 1677247768
transform -1 0 80832 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _229_
timestamp 1677247768
transform -1 0 80736 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  _230_
timestamp 1677247768
transform -1 0 80736 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _231_
timestamp 1677247768
transform 1 0 78432 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _232_
timestamp 1677247768
transform -1 0 80448 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _233_
timestamp 1677247768
transform -1 0 81024 0 1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _234_
timestamp 1677247768
transform -1 0 81312 0 1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _235_
timestamp 1677247768
transform 1 0 80832 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  _236_
timestamp 1677247768
transform -1 0 82272 0 1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  _237_
timestamp 1677247768
transform -1 0 82272 0 1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  _238_
timestamp 1677247768
transform -1 0 82464 0 -1 34020
box -48 -56 1008 834
use sg13g2_a21o_1  _239_
timestamp 1677175127
transform 1 0 1248 0 1 23436
box -48 -56 720 834
use sg13g2_dfrbpq_1  _240_
timestamp 1746535128
transform 1 0 576 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _241_
timestamp 1746535128
transform 1 0 672 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _242_
timestamp 1746535128
transform 1 0 1152 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _243_
timestamp 1746535128
transform 1 0 3360 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _244_
timestamp 1746535128
transform -1 0 5952 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _245_
timestamp 1746535128
transform 1 0 3360 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _246_
timestamp 1746535128
transform 1 0 2784 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _247_
timestamp 1746535128
transform 1 0 2304 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _248_
timestamp 1746535128
transform 1 0 27072 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _249_
timestamp 1746535128
transform 1 0 29280 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _250_
timestamp 1746535128
transform 1 0 31008 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _251_
timestamp 1746535128
transform 1 0 35232 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _252_
timestamp 1746535128
transform 1 0 41568 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _253_
timestamp 1746535128
transform 1 0 50016 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _254_
timestamp 1746535128
transform 1 0 51840 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _255_
timestamp 1746535128
transform 1 0 47424 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _256_
timestamp 1746535128
transform 1 0 44832 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _257_
timestamp 1746535128
transform 1 0 37824 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _258_
timestamp 1746535128
transform 1 0 32256 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _259_
timestamp 1746535128
transform 1 0 34272 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _260_
timestamp 1746535128
transform 1 0 32736 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _261_
timestamp 1746535128
transform 1 0 35712 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _262_
timestamp 1746535128
transform 1 0 46656 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _263_
timestamp 1746535128
transform 1 0 49536 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _264_
timestamp 1746535128
transform 1 0 52704 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _265_
timestamp 1746535128
transform 1 0 55296 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _266_
timestamp 1746535128
transform -1 0 55200 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _267_
timestamp 1746535128
transform -1 0 52608 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _268_
timestamp 1746535128
transform -1 0 50016 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _269_
timestamp 1746535128
transform -1 0 47424 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _270_
timestamp 1746535128
transform 1 0 38880 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _271_
timestamp 1746535128
transform 1 0 37632 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _272_
timestamp 1746535128
transform -1 0 37344 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _273_
timestamp 1746535128
transform 1 0 32064 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _274_
timestamp 1746535128
transform 1 0 30240 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _275_
timestamp 1746535128
transform 1 0 28704 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _276_
timestamp 1746535128
transform 1 0 27648 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _277_
timestamp 1746535128
transform -1 0 21120 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _278_
timestamp 1746535128
transform 1 0 20064 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _279_
timestamp 1746535128
transform 1 0 22560 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _280_
timestamp 1746535128
transform 1 0 22560 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _281_
timestamp 1746535128
transform 1 0 24000 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _282_
timestamp 1746535128
transform 1 0 25920 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _283_
timestamp 1746535128
transform 1 0 40416 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _284_
timestamp 1746535128
transform -1 0 44640 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _285_
timestamp 1746535128
transform -1 0 45792 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _286_
timestamp 1746535128
transform 1 0 3360 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _287_
timestamp 1746535128
transform 1 0 3360 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _288_
timestamp 1746535128
transform 1 0 3360 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _289_
timestamp 1746535128
transform 1 0 9792 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _290_
timestamp 1746535128
transform 1 0 13920 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _291_
timestamp 1746535128
transform 1 0 17952 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _292_
timestamp 1746535128
transform 1 0 15360 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _293_
timestamp 1746535128
transform 1 0 3360 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _294_
timestamp 1746535128
transform 1 0 3360 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _295_
timestamp 1746535128
transform 1 0 2784 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _296_
timestamp 1746535128
transform 1 0 768 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _297_
timestamp 1746535128
transform 1 0 1248 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _298_
timestamp 1746535128
transform 1 0 768 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _299_
timestamp 1746535128
transform 1 0 1920 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _300_
timestamp 1746535128
transform 1 0 768 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _301_
timestamp 1746535128
transform 1 0 2688 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _302_
timestamp 1746535128
transform 1 0 5280 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _303_
timestamp 1746535128
transform 1 0 18048 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _304_
timestamp 1746535128
transform 1 0 21216 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _305_
timestamp 1746535128
transform -1 0 25440 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _306_
timestamp 1746535128
transform 1 0 16800 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _307_
timestamp 1746535128
transform 1 0 13728 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _308_
timestamp 1746535128
transform 1 0 3360 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _309_
timestamp 1746535128
transform 1 0 3360 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _310_
timestamp 1746535128
transform 1 0 3360 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _311_
timestamp 1746535128
transform 1 0 3360 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _312_
timestamp 1746535128
transform 1 0 3360 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _313_
timestamp 1746535128
transform 1 0 76704 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _314_
timestamp 1746535128
transform 1 0 79392 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _315_
timestamp 1746535128
transform 1 0 79392 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _316_
timestamp 1746535128
transform 1 0 79392 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _317_
timestamp 1746535128
transform 1 0 79392 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _318_
timestamp 1746535128
transform 1 0 79392 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _319_
timestamp 1746535128
transform 1 0 79392 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _320_
timestamp 1746535128
transform 1 0 79392 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _321_
timestamp 1746535128
transform 1 0 79392 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _322_
timestamp 1746535128
transform 1 0 81792 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _323_
timestamp 1746535128
transform 1 0 80736 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _324_
timestamp 1746535128
transform 1 0 80736 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _325_
timestamp 1746535128
transform 1 0 80736 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _326_
timestamp 1746535128
transform 1 0 576 0 -1 23436
box -48 -56 2640 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 75456 0 1 12852
box -48 -56 336 834
use sg13g2_buf_16  clkbuf_0_clk_regs
timestamp 1676553496
transform 1 0 42528 0 1 32508
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_0_clk
timestamp 1676553496
transform -1 0 76416 0 -1 17388
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_0__f_clk
timestamp 1676553496
transform 1 0 72000 0 -1 2268
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_1__f_clk
timestamp 1676553496
transform -1 0 81984 0 -1 24948
box -48 -56 2448 834
use sg13g2_buf_8  clkbuf_4_0_0_clk_regs
timestamp 1676451365
transform -1 0 5952 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_1_0_clk_regs
timestamp 1676451365
transform -1 0 5952 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_2_0_clk_regs
timestamp 1676451365
transform -1 0 15360 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_3_0_clk_regs
timestamp 1676451365
transform -1 0 13632 0 1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_4_0_clk_regs
timestamp 1676451365
transform -1 0 34272 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_5_0_clk_regs
timestamp 1676451365
transform -1 0 38112 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_6_0_clk_regs
timestamp 1676451365
transform 1 0 21504 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_7_0_clk_regs
timestamp 1676451365
transform 1 0 25440 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_8_0_clk_regs
timestamp 1676451365
transform -1 0 49344 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_9_0_clk_regs
timestamp 1676451365
transform 1 0 50592 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_10_0_clk_regs
timestamp 1676451365
transform -1 0 50592 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_11_0_clk_regs
timestamp 1676451365
transform 1 0 50112 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_12_0_clk_regs
timestamp 1676451365
transform -1 0 70272 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_13_0_clk_regs
timestamp 1676451365
transform -1 0 66432 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_14_0_clk_regs
timestamp 1676451365
transform 1 0 78432 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_15_0_clk_regs
timestamp 1676451365
transform 1 0 82080 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_16  clkbuf_regs_0_clk
timestamp 1676553496
transform -1 0 44928 0 -1 3780
box -48 -56 2448 834
use sg13g2_inv_1  clkload0
timestamp 1676382929
transform -1 0 4704 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1676382929
transform 1 0 12096 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  clkload2
timestamp 1676382929
transform 1 0 36864 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  clkload3
timestamp 1676382929
transform -1 0 25632 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  clkload4
timestamp 1676382929
transform 1 0 52608 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  clkload5
timestamp 1676382929
transform -1 0 50400 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  clkload6
timestamp 1676382929
transform 1 0 64896 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  clkload7
timestamp 1676382929
transform -1 0 78432 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  clkload8
timestamp 1676382929
transform 1 0 81792 0 -1 30996
box -48 -56 336 834
use sg13g2_buf_16  delaybuf_0_clk
timestamp 1676553496
transform -1 0 39552 0 1 32508
box -48 -56 2448 834
use sg13g2_buf_1  fanout14
timestamp 1676381911
transform 1 0 1152 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout15
timestamp 1676381911
transform -1 0 1536 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout16
timestamp 1676381911
transform -1 0 2208 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout17
timestamp 1676381911
transform 1 0 4128 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout18
timestamp 1676381911
transform 1 0 14976 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout19
timestamp 1676381911
transform 1 0 21216 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout20
timestamp 1676381911
transform -1 0 32352 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  fanout21
timestamp 1676381911
transform 1 0 21504 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout22
timestamp 1676381911
transform 1 0 22848 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout23
timestamp 1676381911
transform 1 0 4512 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform -1 0 42528 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform -1 0 45696 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform -1 0 76512 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform 1 0 81216 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform -1 0 2880 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform -1 0 3360 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout30
timestamp 1676381911
transform 1 0 2592 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform 1 0 960 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout32
timestamp 1676381911
transform 1 0 1632 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform 1 0 1248 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform -1 0 23520 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform -1 0 32928 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform 1 0 21120 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform 1 0 20736 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform -1 0 45312 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform 1 0 42048 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform -1 0 77568 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform 1 0 82176 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform 1 0 1824 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_196
timestamp 1677579658
transform 1 0 19392 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_207
timestamp 1679581782
transform 1 0 20448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_214
timestamp 1679581782
transform 1 0 21120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_221
timestamp 1679581782
transform 1 0 21792 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_228
timestamp 1677579658
transform 1 0 22464 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_256
timestamp 1679581782
transform 1 0 25152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_263
timestamp 1679581782
transform 1 0 25824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_270
timestamp 1679581782
transform 1 0 26496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_277
timestamp 1679581782
transform 1 0 27168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_284
timestamp 1679581782
transform 1 0 27840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_291
timestamp 1679581782
transform 1 0 28512 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_298
timestamp 1677579658
transform 1 0 29184 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_357
timestamp 1679577901
transform 1 0 34848 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_361
timestamp 1677579658
transform 1 0 35232 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_372
timestamp 1679581782
transform 1 0 36288 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_379
timestamp 1679577901
transform 1 0 36960 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_383
timestamp 1677580104
transform 1 0 37344 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_395
timestamp 1679581782
transform 1 0 38496 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_402
timestamp 1677580104
transform 1 0 39168 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_404
timestamp 1677579658
transform 1 0 39360 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_442
timestamp 1679581782
transform 1 0 43008 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_449
timestamp 1679577901
transform 1 0 43680 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_453
timestamp 1677580104
transform 1 0 44064 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_465
timestamp 1679581782
transform 1 0 45216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_472
timestamp 1679581782
transform 1 0 45888 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_479
timestamp 1677580104
transform 1 0 46560 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_491
timestamp 1679581782
transform 1 0 47712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_498
timestamp 1679581782
transform 1 0 48384 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_505
timestamp 1679577901
transform 1 0 49056 0 1 756
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_519
timestamp 1679581782
transform 1 0 50400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_526
timestamp 1679581782
transform 1 0 51072 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_533
timestamp 1677580104
transform 1 0 51744 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_545
timestamp 1679581782
transform 1 0 52896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_552
timestamp 1679581782
transform 1 0 53568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_559
timestamp 1679581782
transform 1 0 54240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_566
timestamp 1679581782
transform 1 0 54912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_573
timestamp 1679581782
transform 1 0 55584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_580
timestamp 1679581782
transform 1 0 56256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_587
timestamp 1679581782
transform 1 0 56928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_594
timestamp 1679581782
transform 1 0 57600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_601
timestamp 1679581782
transform 1 0 58272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_608
timestamp 1679581782
transform 1 0 58944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_615
timestamp 1679581782
transform 1 0 59616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_622
timestamp 1679581782
transform 1 0 60288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_629
timestamp 1679581782
transform 1 0 60960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_636
timestamp 1679581782
transform 1 0 61632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_643
timestamp 1679581782
transform 1 0 62304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_650
timestamp 1679581782
transform 1 0 62976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_657
timestamp 1679581782
transform 1 0 63648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_664
timestamp 1679581782
transform 1 0 64320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_671
timestamp 1679581782
transform 1 0 64992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_678
timestamp 1679581782
transform 1 0 65664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_685
timestamp 1679581782
transform 1 0 66336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_692
timestamp 1679581782
transform 1 0 67008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_699
timestamp 1679581782
transform 1 0 67680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_706
timestamp 1679581782
transform 1 0 68352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_713
timestamp 1679581782
transform 1 0 69024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_720
timestamp 1679581782
transform 1 0 69696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_727
timestamp 1679581782
transform 1 0 70368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_734
timestamp 1679581782
transform 1 0 71040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_741
timestamp 1679581782
transform 1 0 71712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_748
timestamp 1679581782
transform 1 0 72384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_755
timestamp 1679581782
transform 1 0 73056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_762
timestamp 1679581782
transform 1 0 73728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_769
timestamp 1679581782
transform 1 0 74400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_776
timestamp 1679581782
transform 1 0 75072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_783
timestamp 1679581782
transform 1 0 75744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_790
timestamp 1679581782
transform 1 0 76416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_797
timestamp 1679581782
transform 1 0 77088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_804
timestamp 1679581782
transform 1 0 77760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_811
timestamp 1679581782
transform 1 0 78432 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_818
timestamp 1679577901
transform 1 0 79104 0 1 756
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_832
timestamp 1679581782
transform 1 0 80448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_839
timestamp 1679581782
transform 1 0 81120 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_846
timestamp 1677580104
transform 1 0 81792 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_182
timestamp 1679577901
transform 1 0 18048 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_186
timestamp 1677579658
transform 1 0 18432 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_214
timestamp 1679581782
transform 1 0 21120 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_221
timestamp 1677580104
transform 1 0 21792 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_243
timestamp 1677579658
transform 1 0 23904 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_271
timestamp 1677579658
transform 1 0 26592 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_309
timestamp 1679581782
transform 1 0 30240 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_316
timestamp 1677580104
transform 1 0 30912 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_355
timestamp 1677579658
transform 1 0 34656 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_383
timestamp 1677580104
transform 1 0 37344 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_385
timestamp 1677579658
transform 1 0 37536 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_420
timestamp 1677580104
transform 1 0 40896 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_459
timestamp 1677580104
transform 1 0 44640 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_569
timestamp 1679581782
transform 1 0 55200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_576
timestamp 1679581782
transform 1 0 55872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_583
timestamp 1679581782
transform 1 0 56544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_590
timestamp 1679581782
transform 1 0 57216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_597
timestamp 1679581782
transform 1 0 57888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_604
timestamp 1679581782
transform 1 0 58560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_611
timestamp 1679581782
transform 1 0 59232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_618
timestamp 1679581782
transform 1 0 59904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_625
timestamp 1679581782
transform 1 0 60576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_632
timestamp 1679581782
transform 1 0 61248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_639
timestamp 1679581782
transform 1 0 61920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_646
timestamp 1679581782
transform 1 0 62592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_653
timestamp 1679581782
transform 1 0 63264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_660
timestamp 1679581782
transform 1 0 63936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_667
timestamp 1679581782
transform 1 0 64608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_674
timestamp 1679581782
transform 1 0 65280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_681
timestamp 1679581782
transform 1 0 65952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_688
timestamp 1679581782
transform 1 0 66624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_695
timestamp 1679581782
transform 1 0 67296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_702
timestamp 1679581782
transform 1 0 67968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_709
timestamp 1679581782
transform 1 0 68640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_716
timestamp 1679581782
transform 1 0 69312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_723
timestamp 1679581782
transform 1 0 69984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_730
timestamp 1679581782
transform 1 0 70656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_737
timestamp 1679581782
transform 1 0 71328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_769
timestamp 1679581782
transform 1 0 74400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_776
timestamp 1679581782
transform 1 0 75072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_783
timestamp 1679581782
transform 1 0 75744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_790
timestamp 1679581782
transform 1 0 76416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_797
timestamp 1679581782
transform 1 0 77088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_804
timestamp 1679581782
transform 1 0 77760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_165
timestamp 1679577901
transform 1 0 16416 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_200
timestamp 1677580104
transform 1 0 19776 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_202
timestamp 1677579658
transform 1 0 19968 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_230
timestamp 1679577901
transform 1 0 22656 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_234
timestamp 1677579658
transform 1 0 23040 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_239
timestamp 1679581782
transform 1 0 23520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_246
timestamp 1679581782
transform 1 0 24192 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_253
timestamp 1677579658
transform 1 0 24864 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_291
timestamp 1677580104
transform 1 0 28512 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_320
timestamp 1679581782
transform 1 0 31296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_331
timestamp 1679577901
transform 1 0 32352 0 1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_2_362
timestamp 1679577901
transform 1 0 35328 0 1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_2_393
timestamp 1679577901
transform 1 0 38304 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_397
timestamp 1677580104
transform 1 0 38688 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_426
timestamp 1679581782
transform 1 0 41472 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_433
timestamp 1677579658
transform 1 0 42144 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_471
timestamp 1679581782
transform 1 0 45792 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_478
timestamp 1677580104
transform 1 0 46464 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_507
timestamp 1677580104
transform 1 0 49248 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_509
timestamp 1677579658
transform 1 0 49440 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_537
timestamp 1679577901
transform 1 0 52128 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_541
timestamp 1677580104
transform 1 0 52512 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_597
timestamp 1679581782
transform 1 0 57888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_604
timestamp 1679581782
transform 1 0 58560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_611
timestamp 1679581782
transform 1 0 59232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_618
timestamp 1679581782
transform 1 0 59904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_625
timestamp 1679581782
transform 1 0 60576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_632
timestamp 1679581782
transform 1 0 61248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_639
timestamp 1679581782
transform 1 0 61920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_646
timestamp 1679581782
transform 1 0 62592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_653
timestamp 1679581782
transform 1 0 63264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_660
timestamp 1679581782
transform 1 0 63936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_667
timestamp 1679581782
transform 1 0 64608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_674
timestamp 1679581782
transform 1 0 65280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_681
timestamp 1679581782
transform 1 0 65952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_688
timestamp 1679581782
transform 1 0 66624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_695
timestamp 1679581782
transform 1 0 67296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_702
timestamp 1679581782
transform 1 0 67968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_709
timestamp 1679581782
transform 1 0 68640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_716
timestamp 1679581782
transform 1 0 69312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_723
timestamp 1679581782
transform 1 0 69984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_730
timestamp 1679581782
transform 1 0 70656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_737
timestamp 1679581782
transform 1 0 71328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_744
timestamp 1679581782
transform 1 0 72000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_751
timestamp 1679581782
transform 1 0 72672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_758
timestamp 1679581782
transform 1 0 73344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_765
timestamp 1679581782
transform 1 0 74016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_772
timestamp 1679581782
transform 1 0 74688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_779
timestamp 1679581782
transform 1 0 75360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_786
timestamp 1679581782
transform 1 0 76032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_793
timestamp 1679581782
transform 1 0 76704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_800
timestamp 1679581782
transform 1 0 77376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_807
timestamp 1679581782
transform 1 0 78048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_814
timestamp 1679581782
transform 1 0 78720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_123
timestamp 1679577901
transform 1 0 12384 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_3_164
timestamp 1679577901
transform 1 0 16320 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_168
timestamp 1677579658
transform 1 0 16704 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_196
timestamp 1679577901
transform 1 0 19392 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_200
timestamp 1677580104
transform 1 0 19776 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_212
timestamp 1677580104
transform 1 0 20928 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_214
timestamp 1677579658
transform 1 0 21120 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_256
timestamp 1679581782
transform 1 0 25152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_263
timestamp 1679581782
transform 1 0 25824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_270
timestamp 1679581782
transform 1 0 26496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_277
timestamp 1679581782
transform 1 0 27168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_284
timestamp 1679577901
transform 1 0 27840 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679581782
transform 1 0 29184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679581782
transform 1 0 29856 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_312
timestamp 1677580104
transform 1 0 30528 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_320
timestamp 1679581782
transform 1 0 31296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_327
timestamp 1679577901
transform 1 0 31968 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_331
timestamp 1677580104
transform 1 0 32352 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_363
timestamp 1679581782
transform 1 0 35424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_370
timestamp 1679577901
transform 1 0 36096 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_374
timestamp 1677579658
transform 1 0 36480 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_393
timestamp 1679577901
transform 1 0 38304 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_397
timestamp 1677580104
transform 1 0 38688 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_409
timestamp 1679581782
transform 1 0 39840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_416
timestamp 1679581782
transform 1 0 40512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_423
timestamp 1679581782
transform 1 0 41184 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_430
timestamp 1677580104
transform 1 0 41856 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_432
timestamp 1677579658
transform 1 0 42048 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_466
timestamp 1679577901
transform 1 0 45312 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_470
timestamp 1677580104
transform 1 0 45696 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_482
timestamp 1679581782
transform 1 0 46848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_489
timestamp 1679581782
transform 1 0 47520 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_496
timestamp 1677580104
transform 1 0 48192 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_498
timestamp 1677579658
transform 1 0 48384 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_509
timestamp 1679581782
transform 1 0 49440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_516
timestamp 1679581782
transform 1 0 50112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_523
timestamp 1679581782
transform 1 0 50784 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_530
timestamp 1677580104
transform 1 0 51456 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_542
timestamp 1679581782
transform 1 0 52608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_549
timestamp 1679581782
transform 1 0 53280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_556
timestamp 1679577901
transform 1 0 53952 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_560
timestamp 1677579658
transform 1 0 54336 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_571
timestamp 1679581782
transform 1 0 55392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_578
timestamp 1679581782
transform 1 0 56064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_585
timestamp 1679581782
transform 1 0 56736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_592
timestamp 1679581782
transform 1 0 57408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_599
timestamp 1679581782
transform 1 0 58080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_606
timestamp 1679581782
transform 1 0 58752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_613
timestamp 1679581782
transform 1 0 59424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_620
timestamp 1679581782
transform 1 0 60096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_627
timestamp 1679581782
transform 1 0 60768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_634
timestamp 1679581782
transform 1 0 61440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_641
timestamp 1679581782
transform 1 0 62112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_648
timestamp 1679581782
transform 1 0 62784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_655
timestamp 1679581782
transform 1 0 63456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_662
timestamp 1679581782
transform 1 0 64128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_669
timestamp 1679581782
transform 1 0 64800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_676
timestamp 1679581782
transform 1 0 65472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_683
timestamp 1679581782
transform 1 0 66144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_690
timestamp 1679581782
transform 1 0 66816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_697
timestamp 1679581782
transform 1 0 67488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_704
timestamp 1679581782
transform 1 0 68160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_711
timestamp 1679581782
transform 1 0 68832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_718
timestamp 1679581782
transform 1 0 69504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_725
timestamp 1679581782
transform 1 0 70176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_732
timestamp 1679581782
transform 1 0 70848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_739
timestamp 1679581782
transform 1 0 71520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_746
timestamp 1679581782
transform 1 0 72192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_753
timestamp 1679581782
transform 1 0 72864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_760
timestamp 1679581782
transform 1 0 73536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_767
timestamp 1679581782
transform 1 0 74208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_774
timestamp 1679581782
transform 1 0 74880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_781
timestamp 1679581782
transform 1 0 75552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_788
timestamp 1679581782
transform 1 0 76224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_795
timestamp 1679581782
transform 1 0 76896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_802
timestamp 1679581782
transform 1 0 77568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679581782
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679581782
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_823
timestamp 1679581782
transform 1 0 79584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_830
timestamp 1679581782
transform 1 0 80256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_837
timestamp 1679581782
transform 1 0 80928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_844
timestamp 1679577901
transform 1 0 81600 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_53
timestamp 1677580104
transform 1 0 5664 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_55
timestamp 1677579658
transform 1 0 5856 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_765
timestamp 1679581782
transform 1 0 74016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_772
timestamp 1679581782
transform 1 0 74688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_779
timestamp 1679581782
transform 1 0 75360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_786
timestamp 1679581782
transform 1 0 76032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_793
timestamp 1679581782
transform 1 0 76704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_800
timestamp 1679581782
transform 1 0 77376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_807
timestamp 1679581782
transform 1 0 78048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_814
timestamp 1679581782
transform 1 0 78720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_32
timestamp 1679577901
transform 1 0 3648 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_36
timestamp 1677579658
transform 1 0 4032 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_47
timestamp 1679581782
transform 1 0 5088 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_54
timestamp 1677580104
transform 1 0 5760 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_765
timestamp 1679581782
transform 1 0 74016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_772
timestamp 1679581782
transform 1 0 74688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_779
timestamp 1679581782
transform 1 0 75360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_786
timestamp 1679581782
transform 1 0 76032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_793
timestamp 1679581782
transform 1 0 76704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_800
timestamp 1679581782
transform 1 0 77376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_807
timestamp 1679581782
transform 1 0 78048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_814
timestamp 1679581782
transform 1 0 78720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_821
timestamp 1679577901
transform 1 0 79392 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_835
timestamp 1679581782
transform 1 0 80736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_842
timestamp 1679577901
transform 1 0 81408 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_846
timestamp 1677580104
transform 1 0 81792 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_25
timestamp 1679577901
transform 1 0 2976 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_765
timestamp 1679581782
transform 1 0 74016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_772
timestamp 1679581782
transform 1 0 74688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_779
timestamp 1679581782
transform 1 0 75360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_786
timestamp 1679581782
transform 1 0 76032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_793
timestamp 1679581782
transform 1 0 76704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_800
timestamp 1679581782
transform 1 0 77376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_807
timestamp 1679581782
transform 1 0 78048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_814
timestamp 1679581782
transform 1 0 78720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_821
timestamp 1679581782
transform 1 0 79392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_838
timestamp 1679581782
transform 1 0 81024 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_845
timestamp 1677580104
transform 1 0 81696 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_847
timestamp 1677579658
transform 1 0 81888 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_765
timestamp 1679581782
transform 1 0 74016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_772
timestamp 1679581782
transform 1 0 74688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_779
timestamp 1679581782
transform 1 0 75360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_786
timestamp 1679581782
transform 1 0 76032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_793
timestamp 1679581782
transform 1 0 76704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_800
timestamp 1679581782
transform 1 0 77376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_807
timestamp 1679581782
transform 1 0 78048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_814
timestamp 1679581782
transform 1 0 78720 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_4
timestamp 1677580104
transform 1 0 960 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_6
timestamp 1677579658
transform 1 0 1152 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_16
timestamp 1679581782
transform 1 0 2112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_23
timestamp 1679581782
transform 1 0 2784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_40
timestamp 1679581782
transform 1 0 4416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_47
timestamp 1679581782
transform 1 0 5088 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_54
timestamp 1677580104
transform 1 0 5760 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_765
timestamp 1679581782
transform 1 0 74016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_772
timestamp 1679581782
transform 1 0 74688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_779
timestamp 1679581782
transform 1 0 75360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_786
timestamp 1679581782
transform 1 0 76032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_793
timestamp 1679581782
transform 1 0 76704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_800
timestamp 1679581782
transform 1 0 77376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_807
timestamp 1679581782
transform 1 0 78048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_814
timestamp 1679581782
transform 1 0 78720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_821
timestamp 1679581782
transform 1 0 79392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_828
timestamp 1679581782
transform 1 0 80064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_835
timestamp 1679581782
transform 1 0 80736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_842
timestamp 1679577901
transform 1 0 81408 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_846
timestamp 1677580104
transform 1 0 81792 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_25
timestamp 1679577901
transform 1 0 2976 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_765
timestamp 1679581782
transform 1 0 74016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_772
timestamp 1679581782
transform 1 0 74688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_779
timestamp 1679581782
transform 1 0 75360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_786
timestamp 1679581782
transform 1 0 76032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_793
timestamp 1679581782
transform 1 0 76704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_800
timestamp 1679581782
transform 1 0 77376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_807
timestamp 1679581782
transform 1 0 78048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_814
timestamp 1679581782
transform 1 0 78720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_821
timestamp 1679581782
transform 1 0 79392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_828
timestamp 1679581782
transform 1 0 80064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_835
timestamp 1679581782
transform 1 0 80736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_842
timestamp 1679577901
transform 1 0 81408 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_846
timestamp 1677580104
transform 1 0 81792 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_50
timestamp 1679577901
transform 1 0 5376 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_54
timestamp 1677580104
transform 1 0 5760 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_765
timestamp 1679581782
transform 1 0 74016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_772
timestamp 1679581782
transform 1 0 74688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_779
timestamp 1679581782
transform 1 0 75360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_786
timestamp 1679581782
transform 1 0 76032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_793
timestamp 1679581782
transform 1 0 76704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_800
timestamp 1679581782
transform 1 0 77376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_807
timestamp 1679581782
transform 1 0 78048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_814
timestamp 1679581782
transform 1 0 78720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_821
timestamp 1679581782
transform 1 0 79392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_828
timestamp 1679581782
transform 1 0 80064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_835
timestamp 1679581782
transform 1 0 80736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_842
timestamp 1679577901
transform 1 0 81408 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_846
timestamp 1677580104
transform 1 0 81792 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_19
timestamp 1679581782
transform 1 0 2400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_26
timestamp 1679581782
transform 1 0 3072 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_33
timestamp 1677580104
transform 1 0 3744 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_45
timestamp 1679581782
transform 1 0 4896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_52
timestamp 1679577901
transform 1 0 5568 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_765
timestamp 1679581782
transform 1 0 74016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_772
timestamp 1679581782
transform 1 0 74688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_779
timestamp 1679581782
transform 1 0 75360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_786
timestamp 1679581782
transform 1 0 76032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_793
timestamp 1679581782
transform 1 0 76704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_800
timestamp 1679581782
transform 1 0 77376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_807
timestamp 1679581782
transform 1 0 78048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_814
timestamp 1679581782
transform 1 0 78720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_821
timestamp 1679581782
transform 1 0 79392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_828
timestamp 1679581782
transform 1 0 80064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_835
timestamp 1679581782
transform 1 0 80736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_842
timestamp 1679577901
transform 1 0 81408 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_846
timestamp 1677580104
transform 1 0 81792 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_0
timestamp 1677580104
transform 1 0 576 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_765
timestamp 1679581782
transform 1 0 74016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_772
timestamp 1679581782
transform 1 0 74688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_779
timestamp 1679581782
transform 1 0 75360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_786
timestamp 1679581782
transform 1 0 76032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_793
timestamp 1679581782
transform 1 0 76704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_800
timestamp 1679581782
transform 1 0 77376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_807
timestamp 1679581782
transform 1 0 78048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_814
timestamp 1679581782
transform 1 0 78720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_13
timestamp 1679581782
transform 1 0 1824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_20
timestamp 1679581782
transform 1 0 2496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_27
timestamp 1679577901
transform 1 0 3168 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_31
timestamp 1677579658
transform 1 0 3552 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_42
timestamp 1679581782
transform 1 0 4608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_49
timestamp 1679581782
transform 1 0 5280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_765
timestamp 1679581782
transform 1 0 74016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_772
timestamp 1679581782
transform 1 0 74688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_779
timestamp 1679581782
transform 1 0 75360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_786
timestamp 1679581782
transform 1 0 76032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_793
timestamp 1679581782
transform 1 0 76704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_800
timestamp 1679581782
transform 1 0 77376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_807
timestamp 1679581782
transform 1 0 78048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_814
timestamp 1679581782
transform 1 0 78720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_821
timestamp 1679577901
transform 1 0 79392 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_835
timestamp 1679581782
transform 1 0 80736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_842
timestamp 1679577901
transform 1 0 81408 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_846
timestamp 1677580104
transform 1 0 81792 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_4
timestamp 1677580104
transform 1 0 960 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_6
timestamp 1677579658
transform 1 0 1152 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_17
timestamp 1679581782
transform 1 0 2208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_24
timestamp 1679577901
transform 1 0 2880 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_28
timestamp 1677579658
transform 1 0 3264 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_765
timestamp 1679581782
transform 1 0 74016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_772
timestamp 1679581782
transform 1 0 74688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_779
timestamp 1679581782
transform 1 0 75360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_786
timestamp 1679581782
transform 1 0 76032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_793
timestamp 1679581782
transform 1 0 76704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_800
timestamp 1679581782
transform 1 0 77376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_807
timestamp 1679581782
transform 1 0 78048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_814
timestamp 1679581782
transform 1 0 78720 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_0
timestamp 1677580104
transform 1 0 576 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_44
timestamp 1679581782
transform 1 0 4800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_51
timestamp 1679577901
transform 1 0 5472 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_55
timestamp 1677579658
transform 1 0 5856 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_765
timestamp 1679581782
transform 1 0 74016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_772
timestamp 1679581782
transform 1 0 74688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_779
timestamp 1679581782
transform 1 0 75360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_786
timestamp 1679581782
transform 1 0 76032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_793
timestamp 1679577901
transform 1 0 76704 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_797
timestamp 1677579658
transform 1 0 77088 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_802
timestamp 1679581782
transform 1 0 77568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_809
timestamp 1679581782
transform 1 0 78240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_836
timestamp 1679581782
transform 1 0 80832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_843
timestamp 1679577901
transform 1 0 81504 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_847
timestamp 1677579658
transform 1 0 81888 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_4
timestamp 1679577901
transform 1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_8
timestamp 1677579658
transform 1 0 1344 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_16
timestamp 1679581782
transform 1 0 2112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_23
timestamp 1679577901
transform 1 0 2784 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_27
timestamp 1677580104
transform 1 0 3168 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_765
timestamp 1679581782
transform 1 0 74016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_772
timestamp 1679581782
transform 1 0 74688 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_779
timestamp 1677579658
transform 1 0 75360 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_820
timestamp 1677579658
transform 1 0 79296 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_4
timestamp 1677580104
transform 1 0 960 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_6
timestamp 1677579658
transform 1 0 1152 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_17
timestamp 1679581782
transform 1 0 2208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_24
timestamp 1679581782
transform 1 0 2880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_41
timestamp 1679581782
transform 1 0 4512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_48
timestamp 1679581782
transform 1 0 5184 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_55
timestamp 1677579658
transform 1 0 5856 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_765
timestamp 1679581782
transform 1 0 74016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_772
timestamp 1679581782
transform 1 0 74688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_779
timestamp 1679581782
transform 1 0 75360 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_786
timestamp 1677579658
transform 1 0 76032 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_791
timestamp 1679581782
transform 1 0 76512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_798
timestamp 1679581782
transform 1 0 77184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_805
timestamp 1679581782
transform 1 0 77856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_812
timestamp 1679581782
transform 1 0 78528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_819
timestamp 1679581782
transform 1 0 79200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_826
timestamp 1679581782
transform 1 0 79872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_833
timestamp 1679581782
transform 1 0 80544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_840
timestamp 1679581782
transform 1 0 81216 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_847
timestamp 1677579658
transform 1 0 81888 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_0
timestamp 1677580104
transform 1 0 576 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_765
timestamp 1679581782
transform 1 0 74016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_772
timestamp 1679581782
transform 1 0 74688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_779
timestamp 1679581782
transform 1 0 75360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_786
timestamp 1679581782
transform 1 0 76032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_793
timestamp 1679581782
transform 1 0 76704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_800
timestamp 1679581782
transform 1 0 77376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_807
timestamp 1679581782
transform 1 0 78048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_814
timestamp 1679581782
transform 1 0 78720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_821
timestamp 1679581782
transform 1 0 79392 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_828
timestamp 1677580104
transform 1 0 80064 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_830
timestamp 1677579658
transform 1 0 80256 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_841
timestamp 1679581782
transform 1 0 81312 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_4
timestamp 1677580104
transform 1 0 960 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_6
timestamp 1677579658
transform 1 0 1152 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679581782
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_25
timestamp 1679581782
transform 1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_32
timestamp 1679577901
transform 1 0 3648 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_36
timestamp 1677579658
transform 1 0 4032 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_47
timestamp 1679581782
transform 1 0 5088 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_54
timestamp 1677580104
transform 1 0 5760 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_765
timestamp 1679581782
transform 1 0 74016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_772
timestamp 1679581782
transform 1 0 74688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_779
timestamp 1679581782
transform 1 0 75360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_786
timestamp 1679581782
transform 1 0 76032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_793
timestamp 1679581782
transform 1 0 76704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_800
timestamp 1679581782
transform 1 0 77376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_807
timestamp 1679581782
transform 1 0 78048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_814
timestamp 1679581782
transform 1 0 78720 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_4
timestamp 1677580104
transform 1 0 960 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_24
timestamp 1679577901
transform 1 0 2880 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_28
timestamp 1677579658
transform 1 0 3264 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_765
timestamp 1679581782
transform 1 0 74016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_772
timestamp 1679581782
transform 1 0 74688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_779
timestamp 1679581782
transform 1 0 75360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_786
timestamp 1679581782
transform 1 0 76032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_793
timestamp 1679581782
transform 1 0 76704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_800
timestamp 1679581782
transform 1 0 77376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_807
timestamp 1679581782
transform 1 0 78048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_814
timestamp 1679581782
transform 1 0 78720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_821
timestamp 1679581782
transform 1 0 79392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_828
timestamp 1679581782
transform 1 0 80064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_835
timestamp 1679581782
transform 1 0 80736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_842
timestamp 1679577901
transform 1 0 81408 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_846
timestamp 1677580104
transform 1 0 81792 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_8
timestamp 1679577901
transform 1 0 1344 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_12
timestamp 1677580104
transform 1 0 1728 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_41
timestamp 1679581782
transform 1 0 4512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_48
timestamp 1679581782
transform 1 0 5184 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_55
timestamp 1677579658
transform 1 0 5856 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_790
timestamp 1679581782
transform 1 0 76416 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_797
timestamp 1679581782
transform 1 0 77088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_804
timestamp 1679581782
transform 1 0 77760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_811
timestamp 1679581782
transform 1 0 78432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_818
timestamp 1679581782
transform 1 0 79104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_825
timestamp 1679581782
transform 1 0 79776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_832
timestamp 1679581782
transform 1 0 80448 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_839
timestamp 1679581782
transform 1 0 81120 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_846
timestamp 1677580104
transform 1 0 81792 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_4
timestamp 1677580104
transform 1 0 960 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_20
timestamp 1677579658
transform 1 0 2496 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_29
timestamp 1679577901
transform 1 0 3360 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_33
timestamp 1677579658
transform 1 0 3744 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_44
timestamp 1679581782
transform 1 0 4800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_51
timestamp 1679577901
transform 1 0 5472 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_55
timestamp 1677579658
transform 1 0 5856 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_765
timestamp 1679581782
transform 1 0 74016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_772
timestamp 1679581782
transform 1 0 74688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_779
timestamp 1679581782
transform 1 0 75360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_786
timestamp 1679581782
transform 1 0 76032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_793
timestamp 1679581782
transform 1 0 76704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_800
timestamp 1679581782
transform 1 0 77376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_807
timestamp 1679581782
transform 1 0 78048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_814
timestamp 1679581782
transform 1 0 78720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_821
timestamp 1679581782
transform 1 0 79392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_828
timestamp 1679581782
transform 1 0 80064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_835
timestamp 1679581782
transform 1 0 80736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_842
timestamp 1679577901
transform 1 0 81408 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_846
timestamp 1677580104
transform 1 0 81792 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_0
timestamp 1677580104
transform 1 0 576 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_765
timestamp 1679581782
transform 1 0 74016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_772
timestamp 1679581782
transform 1 0 74688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_779
timestamp 1679581782
transform 1 0 75360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_786
timestamp 1679581782
transform 1 0 76032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_793
timestamp 1679581782
transform 1 0 76704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_800
timestamp 1679581782
transform 1 0 77376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_807
timestamp 1679581782
transform 1 0 78048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_814
timestamp 1679581782
transform 1 0 78720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_821
timestamp 1679581782
transform 1 0 79392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_828
timestamp 1679581782
transform 1 0 80064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_835
timestamp 1679581782
transform 1 0 80736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_842
timestamp 1679577901
transform 1 0 81408 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_846
timestamp 1677580104
transform 1 0 81792 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_11
timestamp 1677580104
transform 1 0 1632 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_17
timestamp 1679581782
transform 1 0 2208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_24
timestamp 1679581782
transform 1 0 2880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_31
timestamp 1679581782
transform 1 0 3552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_48
timestamp 1679581782
transform 1 0 5184 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_55
timestamp 1677579658
transform 1 0 5856 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_765
timestamp 1679581782
transform 1 0 74016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_772
timestamp 1679581782
transform 1 0 74688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_779
timestamp 1679581782
transform 1 0 75360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_786
timestamp 1679581782
transform 1 0 76032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_793
timestamp 1679581782
transform 1 0 76704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_800
timestamp 1679581782
transform 1 0 77376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_807
timestamp 1679581782
transform 1 0 78048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_814
timestamp 1679581782
transform 1 0 78720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_821
timestamp 1679581782
transform 1 0 79392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_828
timestamp 1679581782
transform 1 0 80064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_835
timestamp 1679577901
transform 1 0 80736 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_839
timestamp 1677579658
transform 1 0 81120 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_844
timestamp 1679577901
transform 1 0 81600 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_18
timestamp 1677579658
transform 1 0 2304 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_765
timestamp 1679581782
transform 1 0 74016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_772
timestamp 1679581782
transform 1 0 74688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_779
timestamp 1679581782
transform 1 0 75360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_786
timestamp 1679581782
transform 1 0 76032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_793
timestamp 1679581782
transform 1 0 76704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_800
timestamp 1679581782
transform 1 0 77376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_807
timestamp 1679581782
transform 1 0 78048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_814
timestamp 1679581782
transform 1 0 78720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_821
timestamp 1679581782
transform 1 0 79392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_828
timestamp 1679581782
transform 1 0 80064 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_835
timestamp 1677579658
transform 1 0 80736 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_873
timestamp 1679581782
transform 1 0 84384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_880
timestamp 1679581782
transform 1 0 85056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_887
timestamp 1679581782
transform 1 0 85728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_894
timestamp 1679581782
transform 1 0 86400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_901
timestamp 1679581782
transform 1 0 87072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_908
timestamp 1679581782
transform 1 0 87744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_915
timestamp 1679581782
transform 1 0 88416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_922
timestamp 1679581782
transform 1 0 89088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_929
timestamp 1679581782
transform 1 0 89760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_936
timestamp 1679581782
transform 1 0 90432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_943
timestamp 1679581782
transform 1 0 91104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_950
timestamp 1679581782
transform 1 0 91776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_957
timestamp 1679581782
transform 1 0 92448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_964
timestamp 1679581782
transform 1 0 93120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_971
timestamp 1679581782
transform 1 0 93792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_978
timestamp 1679581782
transform 1 0 94464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_985
timestamp 1679581782
transform 1 0 95136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_992
timestamp 1679581782
transform 1 0 95808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_999
timestamp 1679581782
transform 1 0 96480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1006
timestamp 1679581782
transform 1 0 97152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1013
timestamp 1679581782
transform 1 0 97824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1020
timestamp 1679581782
transform 1 0 98496 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_1027
timestamp 1677580104
transform 1 0 99168 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_18
timestamp 1679577901
transform 1 0 2304 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_49
timestamp 1679581782
transform 1 0 5280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_765
timestamp 1679581782
transform 1 0 74016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_772
timestamp 1679581782
transform 1 0 74688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_779
timestamp 1679581782
transform 1 0 75360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_786
timestamp 1679581782
transform 1 0 76032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_793
timestamp 1679581782
transform 1 0 76704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_800
timestamp 1679581782
transform 1 0 77376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_807
timestamp 1679581782
transform 1 0 78048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_814
timestamp 1679581782
transform 1 0 78720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_821
timestamp 1679581782
transform 1 0 79392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_828
timestamp 1679581782
transform 1 0 80064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_835
timestamp 1679581782
transform 1 0 80736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_842
timestamp 1679581782
transform 1 0 81408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_849
timestamp 1679581782
transform 1 0 82080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_856
timestamp 1679581782
transform 1 0 82752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_863
timestamp 1679581782
transform 1 0 83424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_870
timestamp 1679581782
transform 1 0 84096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_877
timestamp 1679581782
transform 1 0 84768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_884
timestamp 1679581782
transform 1 0 85440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_891
timestamp 1679581782
transform 1 0 86112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_898
timestamp 1679581782
transform 1 0 86784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_905
timestamp 1679581782
transform 1 0 87456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_912
timestamp 1679581782
transform 1 0 88128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_919
timestamp 1679581782
transform 1 0 88800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_926
timestamp 1679581782
transform 1 0 89472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_933
timestamp 1679581782
transform 1 0 90144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_940
timestamp 1679581782
transform 1 0 90816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_947
timestamp 1679581782
transform 1 0 91488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_954
timestamp 1679581782
transform 1 0 92160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_961
timestamp 1679581782
transform 1 0 92832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_968
timestamp 1679581782
transform 1 0 93504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_975
timestamp 1679581782
transform 1 0 94176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_982
timestamp 1679581782
transform 1 0 94848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_989
timestamp 1679581782
transform 1 0 95520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_996
timestamp 1679581782
transform 1 0 96192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1003
timestamp 1679581782
transform 1 0 96864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1010
timestamp 1679581782
transform 1 0 97536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1017
timestamp 1679581782
transform 1 0 98208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_1024
timestamp 1679577901
transform 1 0 98880 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_1028
timestamp 1677579658
transform 1 0 99264 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679581782
transform 1 0 3264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_45
timestamp 1679581782
transform 1 0 4896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_52
timestamp 1679577901
transform 1 0 5568 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_765
timestamp 1679581782
transform 1 0 74016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_772
timestamp 1679581782
transform 1 0 74688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_779
timestamp 1679581782
transform 1 0 75360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_786
timestamp 1679581782
transform 1 0 76032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_793
timestamp 1679581782
transform 1 0 76704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_800
timestamp 1679581782
transform 1 0 77376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_807
timestamp 1679581782
transform 1 0 78048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_814
timestamp 1679581782
transform 1 0 78720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_821
timestamp 1679581782
transform 1 0 79392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_828
timestamp 1679581782
transform 1 0 80064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_835
timestamp 1679581782
transform 1 0 80736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_842
timestamp 1679581782
transform 1 0 81408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_849
timestamp 1679581782
transform 1 0 82080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_856
timestamp 1679581782
transform 1 0 82752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_863
timestamp 1679581782
transform 1 0 83424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_870
timestamp 1679581782
transform 1 0 84096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_877
timestamp 1679581782
transform 1 0 84768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_884
timestamp 1679581782
transform 1 0 85440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_891
timestamp 1679581782
transform 1 0 86112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_898
timestamp 1679581782
transform 1 0 86784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_905
timestamp 1679581782
transform 1 0 87456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_912
timestamp 1679581782
transform 1 0 88128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_919
timestamp 1679581782
transform 1 0 88800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_926
timestamp 1679581782
transform 1 0 89472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_933
timestamp 1679581782
transform 1 0 90144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_940
timestamp 1679581782
transform 1 0 90816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_947
timestamp 1679581782
transform 1 0 91488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_954
timestamp 1679581782
transform 1 0 92160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_961
timestamp 1679581782
transform 1 0 92832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_968
timestamp 1679581782
transform 1 0 93504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_975
timestamp 1679581782
transform 1 0 94176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_982
timestamp 1679581782
transform 1 0 94848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_989
timestamp 1679581782
transform 1 0 95520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_996
timestamp 1679581782
transform 1 0 96192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1003
timestamp 1679581782
transform 1 0 96864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1010
timestamp 1679581782
transform 1 0 97536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1017
timestamp 1679581782
transform 1 0 98208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_1024
timestamp 1679577901
transform 1 0 98880 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_1028
timestamp 1677579658
transform 1 0 99264 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_8
timestamp 1679581782
transform 1 0 1344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_15
timestamp 1679581782
transform 1 0 2016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_22
timestamp 1679581782
transform 1 0 2688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_765
timestamp 1679581782
transform 1 0 74016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_772
timestamp 1679581782
transform 1 0 74688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_779
timestamp 1679581782
transform 1 0 75360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_786
timestamp 1679581782
transform 1 0 76032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_793
timestamp 1679581782
transform 1 0 76704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_800
timestamp 1679581782
transform 1 0 77376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_807
timestamp 1679581782
transform 1 0 78048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_814
timestamp 1679581782
transform 1 0 78720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_821
timestamp 1679581782
transform 1 0 79392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_828
timestamp 1679581782
transform 1 0 80064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_835
timestamp 1679581782
transform 1 0 80736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_842
timestamp 1679581782
transform 1 0 81408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_849
timestamp 1679581782
transform 1 0 82080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_856
timestamp 1679577901
transform 1 0 82752 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_860
timestamp 1677580104
transform 1 0 83136 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_27
timestamp 1679581782
transform 1 0 3168 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_34
timestamp 1677580104
transform 1 0 3840 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_36
timestamp 1677579658
transform 1 0 4032 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_45
timestamp 1679581782
transform 1 0 4896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_52
timestamp 1679577901
transform 1 0 5568 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_765
timestamp 1679581782
transform 1 0 74016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_772
timestamp 1679581782
transform 1 0 74688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_779
timestamp 1679581782
transform 1 0 75360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_786
timestamp 1679581782
transform 1 0 76032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_793
timestamp 1679581782
transform 1 0 76704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_800
timestamp 1679581782
transform 1 0 77376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_807
timestamp 1679581782
transform 1 0 78048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_814
timestamp 1679581782
transform 1 0 78720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_821
timestamp 1679581782
transform 1 0 79392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_828
timestamp 1679581782
transform 1 0 80064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_835
timestamp 1679581782
transform 1 0 80736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_842
timestamp 1679581782
transform 1 0 81408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_849
timestamp 1679581782
transform 1 0 82080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_856
timestamp 1679577901
transform 1 0 82752 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_860
timestamp 1677580104
transform 1 0 83136 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_0
timestamp 1677580104
transform 1 0 576 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_19
timestamp 1679577901
transform 1 0 2400 0 1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_30_50
timestamp 1679577901
transform 1 0 5376 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_54
timestamp 1677580104
transform 1 0 5760 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_765
timestamp 1679581782
transform 1 0 74016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_772
timestamp 1679581782
transform 1 0 74688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_779
timestamp 1679581782
transform 1 0 75360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_786
timestamp 1679581782
transform 1 0 76032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_793
timestamp 1679581782
transform 1 0 76704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_800
timestamp 1679581782
transform 1 0 77376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_807
timestamp 1679581782
transform 1 0 78048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_814
timestamp 1679581782
transform 1 0 78720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_821
timestamp 1679581782
transform 1 0 79392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_828
timestamp 1679581782
transform 1 0 80064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_835
timestamp 1679581782
transform 1 0 80736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_842
timestamp 1679581782
transform 1 0 81408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_849
timestamp 1679581782
transform 1 0 82080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_856
timestamp 1679577901
transform 1 0 82752 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_860
timestamp 1677580104
transform 1 0 83136 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_8
timestamp 1679581782
transform 1 0 1344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_18
timestamp 1679581782
transform 1 0 2304 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_25
timestamp 1677579658
transform 1 0 2976 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_41
timestamp 1679581782
transform 1 0 4512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_48
timestamp 1679581782
transform 1 0 5184 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_55
timestamp 1677579658
transform 1 0 5856 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_765
timestamp 1679581782
transform 1 0 74016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_772
timestamp 1679581782
transform 1 0 74688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_779
timestamp 1679581782
transform 1 0 75360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_786
timestamp 1679581782
transform 1 0 76032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_793
timestamp 1679581782
transform 1 0 76704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_800
timestamp 1679581782
transform 1 0 77376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_807
timestamp 1679581782
transform 1 0 78048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_814
timestamp 1679581782
transform 1 0 78720 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_821
timestamp 1677580104
transform 1 0 79392 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_848
timestamp 1679581782
transform 1 0 81984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_855
timestamp 1679581782
transform 1 0 82656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_16
timestamp 1679581782
transform 1 0 2112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_23
timestamp 1679577901
transform 1 0 2784 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_27
timestamp 1677580104
transform 1 0 3168 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_765
timestamp 1679581782
transform 1 0 74016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_772
timestamp 1679581782
transform 1 0 74688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_779
timestamp 1679581782
transform 1 0 75360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_786
timestamp 1679581782
transform 1 0 76032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_793
timestamp 1679581782
transform 1 0 76704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_800
timestamp 1679581782
transform 1 0 77376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_807
timestamp 1679581782
transform 1 0 78048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_814
timestamp 1679581782
transform 1 0 78720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_821
timestamp 1679581782
transform 1 0 79392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_828
timestamp 1679581782
transform 1 0 80064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_835
timestamp 1679581782
transform 1 0 80736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_842
timestamp 1679581782
transform 1 0 81408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_849
timestamp 1679581782
transform 1 0 82080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_856
timestamp 1679577901
transform 1 0 82752 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_860
timestamp 1677580104
transform 1 0 83136 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_46
timestamp 1679581782
transform 1 0 4992 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_53
timestamp 1677580104
transform 1 0 5664 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_55
timestamp 1677579658
transform 1 0 5856 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_765
timestamp 1679581782
transform 1 0 74016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_772
timestamp 1679581782
transform 1 0 74688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_779
timestamp 1679581782
transform 1 0 75360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_786
timestamp 1679581782
transform 1 0 76032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_793
timestamp 1679581782
transform 1 0 76704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_800
timestamp 1679581782
transform 1 0 77376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_807
timestamp 1679581782
transform 1 0 78048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_814
timestamp 1679581782
transform 1 0 78720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_821
timestamp 1679581782
transform 1 0 79392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_828
timestamp 1679581782
transform 1 0 80064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_835
timestamp 1679581782
transform 1 0 80736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_842
timestamp 1679581782
transform 1 0 81408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_849
timestamp 1679581782
transform 1 0 82080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_856
timestamp 1679577901
transform 1 0 82752 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_860
timestamp 1677580104
transform 1 0 83136 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_0
timestamp 1679577901
transform 1 0 576 0 1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_34_13
timestamp 1679577901
transform 1 0 1824 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_17
timestamp 1677579658
transform 1 0 2208 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_23
timestamp 1679577901
transform 1 0 2784 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_44
timestamp 1679581782
transform 1 0 4800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_51
timestamp 1679577901
transform 1 0 5472 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_55
timestamp 1677579658
transform 1 0 5856 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_765
timestamp 1679581782
transform 1 0 74016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_772
timestamp 1679581782
transform 1 0 74688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_779
timestamp 1679581782
transform 1 0 75360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_786
timestamp 1679581782
transform 1 0 76032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_793
timestamp 1679581782
transform 1 0 76704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_800
timestamp 1679581782
transform 1 0 77376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_807
timestamp 1679581782
transform 1 0 78048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_814
timestamp 1679581782
transform 1 0 78720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_821
timestamp 1679581782
transform 1 0 79392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_828
timestamp 1679581782
transform 1 0 80064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_835
timestamp 1679577901
transform 1 0 80736 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_839
timestamp 1677580104
transform 1 0 81120 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_851
timestamp 1679581782
transform 1 0 82272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_858
timestamp 1679577901
transform 1 0 82944 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_7
timestamp 1679577901
transform 1 0 1248 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_11
timestamp 1677579658
transform 1 0 1632 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_19
timestamp 1677580104
transform 1 0 2400 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_21
timestamp 1677579658
transform 1 0 2592 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_27
timestamp 1677580104
transform 1 0 3168 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_765
timestamp 1679581782
transform 1 0 74016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_772
timestamp 1679581782
transform 1 0 74688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_779
timestamp 1679581782
transform 1 0 75360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_786
timestamp 1679581782
transform 1 0 76032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_793
timestamp 1679581782
transform 1 0 76704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_800
timestamp 1679581782
transform 1 0 77376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_807
timestamp 1679581782
transform 1 0 78048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_814
timestamp 1679581782
transform 1 0 78720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_821
timestamp 1679581782
transform 1 0 79392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_828
timestamp 1679581782
transform 1 0 80064 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_0
timestamp 1677579658
transform 1 0 576 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_765
timestamp 1679581782
transform 1 0 74016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_772
timestamp 1679581782
transform 1 0 74688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_779
timestamp 1679581782
transform 1 0 75360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_786
timestamp 1679581782
transform 1 0 76032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_793
timestamp 1679581782
transform 1 0 76704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_800
timestamp 1679581782
transform 1 0 77376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_807
timestamp 1679581782
transform 1 0 78048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_814
timestamp 1679581782
transform 1 0 78720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_821
timestamp 1679581782
transform 1 0 79392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_828
timestamp 1679581782
transform 1 0 80064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_835
timestamp 1679581782
transform 1 0 80736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_842
timestamp 1679581782
transform 1 0 81408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_849
timestamp 1679581782
transform 1 0 82080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_856
timestamp 1679577901
transform 1 0 82752 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_860
timestamp 1677580104
transform 1 0 83136 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_7
timestamp 1677580104
transform 1 0 1248 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_18
timestamp 1677580104
transform 1 0 2304 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_20
timestamp 1677579658
transform 1 0 2496 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_27
timestamp 1677579658
transform 1 0 3168 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_38
timestamp 1677580104
transform 1 0 4224 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_765
timestamp 1679581782
transform 1 0 74016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_772
timestamp 1679581782
transform 1 0 74688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_779
timestamp 1679581782
transform 1 0 75360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_786
timestamp 1679581782
transform 1 0 76032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_793
timestamp 1679581782
transform 1 0 76704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_800
timestamp 1679581782
transform 1 0 77376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_807
timestamp 1679581782
transform 1 0 78048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_814
timestamp 1679581782
transform 1 0 78720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_821
timestamp 1679581782
transform 1 0 79392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_828
timestamp 1679581782
transform 1 0 80064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_835
timestamp 1679581782
transform 1 0 80736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_842
timestamp 1679581782
transform 1 0 81408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_849
timestamp 1679581782
transform 1 0 82080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_856
timestamp 1679577901
transform 1 0 82752 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_860
timestamp 1677580104
transform 1 0 83136 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_38_0
timestamp 1679577901
transform 1 0 576 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_4
timestamp 1677579658
transform 1 0 960 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_23
timestamp 1679577901
transform 1 0 2784 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_27
timestamp 1677580104
transform 1 0 3168 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_765
timestamp 1679581782
transform 1 0 74016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_772
timestamp 1679581782
transform 1 0 74688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_779
timestamp 1679581782
transform 1 0 75360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_786
timestamp 1679581782
transform 1 0 76032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_793
timestamp 1679581782
transform 1 0 76704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_800
timestamp 1679581782
transform 1 0 77376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_807
timestamp 1679581782
transform 1 0 78048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_814
timestamp 1679581782
transform 1 0 78720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_821
timestamp 1679581782
transform 1 0 79392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_828
timestamp 1679581782
transform 1 0 80064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_835
timestamp 1679581782
transform 1 0 80736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_842
timestamp 1679581782
transform 1 0 81408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_849
timestamp 1679581782
transform 1 0 82080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_856
timestamp 1679577901
transform 1 0 82752 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_860
timestamp 1677580104
transform 1 0 83136 0 1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_39_0
timestamp 1679577901
transform 1 0 576 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_4
timestamp 1677580104
transform 1 0 960 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_33
timestamp 1679581782
transform 1 0 3744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_40
timestamp 1679581782
transform 1 0 4416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_47
timestamp 1679581782
transform 1 0 5088 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_54
timestamp 1677580104
transform 1 0 5760 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_765
timestamp 1679581782
transform 1 0 74016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_772
timestamp 1679581782
transform 1 0 74688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_779
timestamp 1679581782
transform 1 0 75360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_786
timestamp 1679581782
transform 1 0 76032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_793
timestamp 1679581782
transform 1 0 76704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_800
timestamp 1679581782
transform 1 0 77376 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_807
timestamp 1677579658
transform 1 0 78048 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_824
timestamp 1679581782
transform 1 0 79680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_831
timestamp 1679581782
transform 1 0 80352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_838
timestamp 1679581782
transform 1 0 81024 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_845
timestamp 1677579658
transform 1 0 81696 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_15
timestamp 1677580104
transform 1 0 2016 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_17
timestamp 1677579658
transform 1 0 2208 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_55
timestamp 1677579658
transform 1 0 5856 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_765
timestamp 1679581782
transform 1 0 74016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_772
timestamp 1679581782
transform 1 0 74688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_779
timestamp 1679581782
transform 1 0 75360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_786
timestamp 1679581782
transform 1 0 76032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_793
timestamp 1679581782
transform 1 0 76704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_800
timestamp 1679581782
transform 1 0 77376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_807
timestamp 1679581782
transform 1 0 78048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_814
timestamp 1679581782
transform 1 0 78720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_821
timestamp 1679581782
transform 1 0 79392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_828
timestamp 1679581782
transform 1 0 80064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_835
timestamp 1679577901
transform 1 0 80736 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_839
timestamp 1677580104
transform 1 0 81120 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_851
timestamp 1679581782
transform 1 0 82272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_858
timestamp 1679577901
transform 1 0 82944 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_7
timestamp 1679577901
transform 1 0 1248 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_11
timestamp 1677580104
transform 1 0 1632 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_17
timestamp 1679581782
transform 1 0 2208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_24
timestamp 1679581782
transform 1 0 2880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_31
timestamp 1679581782
transform 1 0 3552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_38
timestamp 1679581782
transform 1 0 4224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_45
timestamp 1679581782
transform 1 0 4896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_52
timestamp 1679577901
transform 1 0 5568 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_765
timestamp 1679581782
transform 1 0 74016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_772
timestamp 1679581782
transform 1 0 74688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_779
timestamp 1679581782
transform 1 0 75360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_786
timestamp 1679581782
transform 1 0 76032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_793
timestamp 1679581782
transform 1 0 76704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_800
timestamp 1679581782
transform 1 0 77376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_807
timestamp 1679581782
transform 1 0 78048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_814
timestamp 1679581782
transform 1 0 78720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_821
timestamp 1679581782
transform 1 0 79392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_828
timestamp 1679581782
transform 1 0 80064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_76
timestamp 1679581782
transform 1 0 7872 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_83
timestamp 1677580104
transform 1 0 8544 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_95
timestamp 1677579658
transform 1 0 9696 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_123
timestamp 1679581782
transform 1 0 12384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_130
timestamp 1679577901
transform 1 0 13056 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_134
timestamp 1677580104
transform 1 0 13440 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_146
timestamp 1679581782
transform 1 0 14592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_163
timestamp 1679581782
transform 1 0 16224 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_170
timestamp 1677580104
transform 1 0 16896 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_209
timestamp 1679577901
transform 1 0 20640 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_213
timestamp 1677580104
transform 1 0 21024 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_242
timestamp 1679581782
transform 1 0 23808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_249
timestamp 1679581782
transform 1 0 24480 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_256
timestamp 1677580104
transform 1 0 25152 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_261
timestamp 1679581782
transform 1 0 25632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_268
timestamp 1679581782
transform 1 0 26304 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_275
timestamp 1677579658
transform 1 0 26976 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_286
timestamp 1679581782
transform 1 0 28032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_293
timestamp 1679577901
transform 1 0 28704 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_297
timestamp 1677580104
transform 1 0 29088 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_326
timestamp 1679581782
transform 1 0 31872 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_333
timestamp 1679577901
transform 1 0 32544 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_337
timestamp 1677579658
transform 1 0 32928 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679581782
transform 1 0 39552 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_413
timestamp 1677580104
transform 1 0 40224 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_425
timestamp 1679581782
transform 1 0 41376 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_436
timestamp 1677579658
transform 1 0 42432 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_462
timestamp 1677580104
transform 1 0 44928 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_464
timestamp 1677579658
transform 1 0 45120 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_475
timestamp 1679581782
transform 1 0 46176 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_482
timestamp 1677580104
transform 1 0 46848 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_484
timestamp 1677579658
transform 1 0 47040 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_561
timestamp 1679581782
transform 1 0 54432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_568
timestamp 1679581782
transform 1 0 55104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_575
timestamp 1679581782
transform 1 0 55776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_582
timestamp 1679581782
transform 1 0 56448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_589
timestamp 1679581782
transform 1 0 57120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_596
timestamp 1679581782
transform 1 0 57792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_603
timestamp 1679581782
transform 1 0 58464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_610
timestamp 1679581782
transform 1 0 59136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_617
timestamp 1679581782
transform 1 0 59808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_624
timestamp 1679581782
transform 1 0 60480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_631
timestamp 1679581782
transform 1 0 61152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_638
timestamp 1679581782
transform 1 0 61824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_645
timestamp 1679581782
transform 1 0 62496 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_652
timestamp 1679581782
transform 1 0 63168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_659
timestamp 1679581782
transform 1 0 63840 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_666
timestamp 1679577901
transform 1 0 64512 0 1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_42_686
timestamp 1679581782
transform 1 0 66432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_693
timestamp 1679581782
transform 1 0 67104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_700
timestamp 1679581782
transform 1 0 67776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_707
timestamp 1679577901
transform 1 0 68448 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_711
timestamp 1677580104
transform 1 0 68832 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_726
timestamp 1679581782
transform 1 0 70272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_733
timestamp 1679581782
transform 1 0 70944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_740
timestamp 1679581782
transform 1 0 71616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_747
timestamp 1679581782
transform 1 0 72288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_754
timestamp 1679581782
transform 1 0 72960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_761
timestamp 1679581782
transform 1 0 73632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_768
timestamp 1679581782
transform 1 0 74304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_775
timestamp 1679581782
transform 1 0 74976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_782
timestamp 1679581782
transform 1 0 75648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_789
timestamp 1679581782
transform 1 0 76320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_796
timestamp 1679581782
transform 1 0 76992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_803
timestamp 1679581782
transform 1 0 77664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_810
timestamp 1679581782
transform 1 0 78336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_817
timestamp 1679581782
transform 1 0 79008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_824
timestamp 1679581782
transform 1 0 79680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_831
timestamp 1679581782
transform 1 0 80352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_838
timestamp 1679581782
transform 1 0 81024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_845
timestamp 1679581782
transform 1 0 81696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_852
timestamp 1679581782
transform 1 0 82368 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_859
timestamp 1677580104
transform 1 0 83040 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_861
timestamp 1677579658
transform 1 0 83232 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_133
timestamp 1679577901
transform 1 0 13344 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_137
timestamp 1677580104
transform 1 0 13728 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_166
timestamp 1677580104
transform 1 0 16512 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_168
timestamp 1677579658
transform 1 0 16704 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_179
timestamp 1679581782
transform 1 0 17760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_186
timestamp 1679581782
transform 1 0 18432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_193
timestamp 1679581782
transform 1 0 19104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_200
timestamp 1679581782
transform 1 0 19776 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_207
timestamp 1677579658
transform 1 0 20448 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_231
timestamp 1677579658
transform 1 0 22752 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_43_272
timestamp 1679577901
transform 1 0 26688 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_4  FILLER_43_303
timestamp 1679577901
transform 1 0 29664 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_354
timestamp 1679581782
transform 1 0 34560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_415
timestamp 1679581782
transform 1 0 40416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_422
timestamp 1679577901
transform 1 0 41088 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_426
timestamp 1677579658
transform 1 0 41472 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_454
timestamp 1679581782
transform 1 0 44160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_545
timestamp 1679581782
transform 1 0 52896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_552
timestamp 1679581782
transform 1 0 53568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_559
timestamp 1679581782
transform 1 0 54240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_566
timestamp 1679581782
transform 1 0 54912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_573
timestamp 1679581782
transform 1 0 55584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_580
timestamp 1679581782
transform 1 0 56256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_587
timestamp 1679581782
transform 1 0 56928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_594
timestamp 1679581782
transform 1 0 57600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_601
timestamp 1679581782
transform 1 0 58272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_608
timestamp 1679581782
transform 1 0 58944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_615
timestamp 1679581782
transform 1 0 59616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_622
timestamp 1679581782
transform 1 0 60288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_629
timestamp 1679581782
transform 1 0 60960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_636
timestamp 1679581782
transform 1 0 61632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_643
timestamp 1679581782
transform 1 0 62304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_650
timestamp 1679581782
transform 1 0 62976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_657
timestamp 1679581782
transform 1 0 63648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_664
timestamp 1679581782
transform 1 0 64320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_671
timestamp 1679581782
transform 1 0 64992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_678
timestamp 1679581782
transform 1 0 65664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_685
timestamp 1679581782
transform 1 0 66336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_692
timestamp 1679581782
transform 1 0 67008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_699
timestamp 1679581782
transform 1 0 67680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_706
timestamp 1679581782
transform 1 0 68352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_713
timestamp 1679581782
transform 1 0 69024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_720
timestamp 1679581782
transform 1 0 69696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_727
timestamp 1679581782
transform 1 0 70368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_734
timestamp 1679581782
transform 1 0 71040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_741
timestamp 1679581782
transform 1 0 71712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_748
timestamp 1679581782
transform 1 0 72384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_755
timestamp 1679581782
transform 1 0 73056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_762
timestamp 1679581782
transform 1 0 73728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_769
timestamp 1679581782
transform 1 0 74400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_776
timestamp 1679581782
transform 1 0 75072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_783
timestamp 1679581782
transform 1 0 75744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_790
timestamp 1679581782
transform 1 0 76416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_797
timestamp 1679581782
transform 1 0 77088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_804
timestamp 1679581782
transform 1 0 77760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_811
timestamp 1679581782
transform 1 0 78432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_818
timestamp 1679581782
transform 1 0 79104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_825
timestamp 1679581782
transform 1 0 79776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_832
timestamp 1679581782
transform 1 0 80448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_839
timestamp 1679577901
transform 1 0 81120 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_853
timestamp 1679581782
transform 1 0 82464 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_860
timestamp 1677580104
transform 1 0 83136 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679581782
transform 1 0 6624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679581782
transform 1 0 7296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679581782
transform 1 0 7968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679581782
transform 1 0 8640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679581782
transform 1 0 9312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679581782
transform 1 0 9984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679581782
transform 1 0 10656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679581782
transform 1 0 11328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679581782
transform 1 0 12000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679581782
transform 1 0 12672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679581782
transform 1 0 13344 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_140
timestamp 1677579658
transform 1 0 14016 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_208
timestamp 1677580104
transform 1 0 20544 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_236
timestamp 1679581782
transform 1 0 23232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_243
timestamp 1679581782
transform 1 0 23904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_250
timestamp 1679581782
transform 1 0 24576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_257
timestamp 1679581782
transform 1 0 25248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_264
timestamp 1679581782
transform 1 0 25920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_271
timestamp 1679581782
transform 1 0 26592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_278
timestamp 1679581782
transform 1 0 27264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_285
timestamp 1679581782
transform 1 0 27936 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_292
timestamp 1677580104
transform 1 0 28608 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_294
timestamp 1677579658
transform 1 0 28800 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_305
timestamp 1679581782
transform 1 0 29856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_312
timestamp 1679581782
transform 1 0 30528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_319
timestamp 1679581782
transform 1 0 31200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_326
timestamp 1679577901
transform 1 0 31872 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679581782
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679581782
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679581782
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_401
timestamp 1679581782
transform 1 0 39072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_408
timestamp 1679581782
transform 1 0 39744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_415
timestamp 1679581782
transform 1 0 40416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_422
timestamp 1679581782
transform 1 0 41088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_429
timestamp 1679581782
transform 1 0 41760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_436
timestamp 1679581782
transform 1 0 42432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_443
timestamp 1679581782
transform 1 0 43104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_450
timestamp 1679581782
transform 1 0 43776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_457
timestamp 1679581782
transform 1 0 44448 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_464
timestamp 1677580104
transform 1 0 45120 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_470
timestamp 1679581782
transform 1 0 45696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_477
timestamp 1679581782
transform 1 0 46368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_484
timestamp 1679581782
transform 1 0 47040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_491
timestamp 1679581782
transform 1 0 47712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_498
timestamp 1679581782
transform 1 0 48384 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_505
timestamp 1677579658
transform 1 0 49056 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_539
timestamp 1679581782
transform 1 0 52320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_546
timestamp 1679581782
transform 1 0 52992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_553
timestamp 1679581782
transform 1 0 53664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_560
timestamp 1679581782
transform 1 0 54336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_567
timestamp 1679581782
transform 1 0 55008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_574
timestamp 1679581782
transform 1 0 55680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_581
timestamp 1679581782
transform 1 0 56352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_588
timestamp 1679581782
transform 1 0 57024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_595
timestamp 1679581782
transform 1 0 57696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_602
timestamp 1679581782
transform 1 0 58368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_609
timestamp 1679581782
transform 1 0 59040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_616
timestamp 1679581782
transform 1 0 59712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_623
timestamp 1679581782
transform 1 0 60384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_630
timestamp 1679581782
transform 1 0 61056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_637
timestamp 1679581782
transform 1 0 61728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_644
timestamp 1679581782
transform 1 0 62400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_651
timestamp 1679581782
transform 1 0 63072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_658
timestamp 1679581782
transform 1 0 63744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_665
timestamp 1679581782
transform 1 0 64416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_672
timestamp 1679581782
transform 1 0 65088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_679
timestamp 1679581782
transform 1 0 65760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_686
timestamp 1679581782
transform 1 0 66432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_693
timestamp 1679581782
transform 1 0 67104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_700
timestamp 1679581782
transform 1 0 67776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_707
timestamp 1679581782
transform 1 0 68448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_714
timestamp 1679581782
transform 1 0 69120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_721
timestamp 1679581782
transform 1 0 69792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_728
timestamp 1679581782
transform 1 0 70464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_735
timestamp 1679581782
transform 1 0 71136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_742
timestamp 1679581782
transform 1 0 71808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_749
timestamp 1679581782
transform 1 0 72480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_756
timestamp 1679581782
transform 1 0 73152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_763
timestamp 1679581782
transform 1 0 73824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_770
timestamp 1679581782
transform 1 0 74496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_777
timestamp 1679581782
transform 1 0 75168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_784
timestamp 1679581782
transform 1 0 75840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_791
timestamp 1679581782
transform 1 0 76512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_798
timestamp 1679581782
transform 1 0 77184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_805
timestamp 1679581782
transform 1 0 77856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_812
timestamp 1679581782
transform 1 0 78528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_819
timestamp 1679581782
transform 1 0 79200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_826
timestamp 1679581782
transform 1 0 79872 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_833
timestamp 1677580104
transform 1 0 80544 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_147
timestamp 1677580104
transform 1 0 14688 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_149
timestamp 1677579658
transform 1 0 14880 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_329
timestamp 1677579658
transform 1 0 32160 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_45_340
timestamp 1679577901
transform 1 0 33216 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_354
timestamp 1679581782
transform 1 0 34560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_361
timestamp 1679581782
transform 1 0 35232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_368
timestamp 1679581782
transform 1 0 35904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_375
timestamp 1679581782
transform 1 0 36576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_382
timestamp 1679581782
transform 1 0 37248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_389
timestamp 1679581782
transform 1 0 37920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_396
timestamp 1679581782
transform 1 0 38592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_403
timestamp 1679581782
transform 1 0 39264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_410
timestamp 1679581782
transform 1 0 39936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_417
timestamp 1679581782
transform 1 0 40608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_424
timestamp 1679581782
transform 1 0 41280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_431
timestamp 1679581782
transform 1 0 41952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_438
timestamp 1679581782
transform 1 0 42624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_445
timestamp 1679581782
transform 1 0 43296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_452
timestamp 1679581782
transform 1 0 43968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_459
timestamp 1679581782
transform 1 0 44640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_466
timestamp 1679581782
transform 1 0 45312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_473
timestamp 1679581782
transform 1 0 45984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_480
timestamp 1679581782
transform 1 0 46656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_487
timestamp 1679581782
transform 1 0 47328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_494
timestamp 1679581782
transform 1 0 48000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_501
timestamp 1679581782
transform 1 0 48672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_508
timestamp 1679581782
transform 1 0 49344 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_515
timestamp 1677579658
transform 1 0 50016 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_519
timestamp 1679581782
transform 1 0 50400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_526
timestamp 1679581782
transform 1 0 51072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_533
timestamp 1679581782
transform 1 0 51744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_540
timestamp 1679581782
transform 1 0 52416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_547
timestamp 1679581782
transform 1 0 53088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_554
timestamp 1679581782
transform 1 0 53760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_561
timestamp 1679581782
transform 1 0 54432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_568
timestamp 1679581782
transform 1 0 55104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_575
timestamp 1679581782
transform 1 0 55776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_582
timestamp 1679581782
transform 1 0 56448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_589
timestamp 1679581782
transform 1 0 57120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_596
timestamp 1679581782
transform 1 0 57792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_603
timestamp 1679581782
transform 1 0 58464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_610
timestamp 1679581782
transform 1 0 59136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_617
timestamp 1679581782
transform 1 0 59808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_624
timestamp 1679581782
transform 1 0 60480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_631
timestamp 1679581782
transform 1 0 61152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_638
timestamp 1679581782
transform 1 0 61824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_645
timestamp 1679581782
transform 1 0 62496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_652
timestamp 1679581782
transform 1 0 63168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_659
timestamp 1679581782
transform 1 0 63840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_666
timestamp 1679581782
transform 1 0 64512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_673
timestamp 1679581782
transform 1 0 65184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_680
timestamp 1679581782
transform 1 0 65856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_687
timestamp 1679581782
transform 1 0 66528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_694
timestamp 1679581782
transform 1 0 67200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_701
timestamp 1679581782
transform 1 0 67872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_708
timestamp 1679581782
transform 1 0 68544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_715
timestamp 1679581782
transform 1 0 69216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_722
timestamp 1679581782
transform 1 0 69888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_729
timestamp 1679581782
transform 1 0 70560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_736
timestamp 1679581782
transform 1 0 71232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_743
timestamp 1679581782
transform 1 0 71904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_750
timestamp 1679581782
transform 1 0 72576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_757
timestamp 1679581782
transform 1 0 73248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_764
timestamp 1679581782
transform 1 0 73920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_771
timestamp 1679581782
transform 1 0 74592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_778
timestamp 1679581782
transform 1 0 75264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_785
timestamp 1679581782
transform 1 0 75936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_792
timestamp 1679581782
transform 1 0 76608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_799
timestamp 1679581782
transform 1 0 77280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_806
timestamp 1679581782
transform 1 0 77952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_813
timestamp 1679581782
transform 1 0 78624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_820
timestamp 1679581782
transform 1 0 79296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_827
timestamp 1679581782
transform 1 0 79968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_834
timestamp 1679581782
transform 1 0 80640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_841
timestamp 1679581782
transform 1 0 81312 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_848
timestamp 1677580104
transform 1 0 81984 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_854
timestamp 1679581782
transform 1 0 82560 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_861
timestamp 1677579658
transform 1 0 83232 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_119
timestamp 1677579658
transform 1 0 12000 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_136
timestamp 1679581782
transform 1 0 13632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_143
timestamp 1679581782
transform 1 0 14304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_150
timestamp 1679581782
transform 1 0 14976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_157
timestamp 1679581782
transform 1 0 15648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_164
timestamp 1679581782
transform 1 0 16320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_171
timestamp 1679581782
transform 1 0 16992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_178
timestamp 1679581782
transform 1 0 17664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_185
timestamp 1679581782
transform 1 0 18336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_192
timestamp 1679581782
transform 1 0 19008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_199
timestamp 1679581782
transform 1 0 19680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_206
timestamp 1679581782
transform 1 0 20352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_213
timestamp 1679581782
transform 1 0 21024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_220
timestamp 1679581782
transform 1 0 21696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_227
timestamp 1679581782
transform 1 0 22368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_234
timestamp 1679581782
transform 1 0 23040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_241
timestamp 1679581782
transform 1 0 23712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_248
timestamp 1679581782
transform 1 0 24384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_255
timestamp 1679581782
transform 1 0 25056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_262
timestamp 1679581782
transform 1 0 25728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_269
timestamp 1679581782
transform 1 0 26400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_276
timestamp 1679581782
transform 1 0 27072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_283
timestamp 1679581782
transform 1 0 27744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_290
timestamp 1679581782
transform 1 0 28416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_297
timestamp 1679581782
transform 1 0 29088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_304
timestamp 1679581782
transform 1 0 29760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_311
timestamp 1679581782
transform 1 0 30432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_318
timestamp 1679581782
transform 1 0 31104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_325
timestamp 1679581782
transform 1 0 31776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_332
timestamp 1679581782
transform 1 0 32448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_339
timestamp 1679581782
transform 1 0 33120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_346
timestamp 1679581782
transform 1 0 33792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_353
timestamp 1679581782
transform 1 0 34464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_360
timestamp 1679581782
transform 1 0 35136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_367
timestamp 1679581782
transform 1 0 35808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_374
timestamp 1679581782
transform 1 0 36480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_381
timestamp 1679581782
transform 1 0 37152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_388
timestamp 1679581782
transform 1 0 37824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_395
timestamp 1679581782
transform 1 0 38496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_402
timestamp 1679581782
transform 1 0 39168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_409
timestamp 1679581782
transform 1 0 39840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_416
timestamp 1679581782
transform 1 0 40512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_423
timestamp 1679581782
transform 1 0 41184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_430
timestamp 1679581782
transform 1 0 41856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_437
timestamp 1679581782
transform 1 0 42528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_444
timestamp 1679581782
transform 1 0 43200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_451
timestamp 1679581782
transform 1 0 43872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_458
timestamp 1679581782
transform 1 0 44544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_465
timestamp 1679581782
transform 1 0 45216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_472
timestamp 1679581782
transform 1 0 45888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_479
timestamp 1679581782
transform 1 0 46560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_486
timestamp 1679581782
transform 1 0 47232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_493
timestamp 1679581782
transform 1 0 47904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_500
timestamp 1679581782
transform 1 0 48576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_507
timestamp 1679581782
transform 1 0 49248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_514
timestamp 1679581782
transform 1 0 49920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_521
timestamp 1679581782
transform 1 0 50592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_528
timestamp 1679581782
transform 1 0 51264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_535
timestamp 1679581782
transform 1 0 51936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_542
timestamp 1679581782
transform 1 0 52608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_549
timestamp 1679581782
transform 1 0 53280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_556
timestamp 1679581782
transform 1 0 53952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_563
timestamp 1679581782
transform 1 0 54624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_570
timestamp 1679581782
transform 1 0 55296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_577
timestamp 1679581782
transform 1 0 55968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_584
timestamp 1679581782
transform 1 0 56640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_591
timestamp 1679581782
transform 1 0 57312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_598
timestamp 1679581782
transform 1 0 57984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_605
timestamp 1679581782
transform 1 0 58656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_612
timestamp 1679581782
transform 1 0 59328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_619
timestamp 1679581782
transform 1 0 60000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_626
timestamp 1679581782
transform 1 0 60672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_633
timestamp 1679581782
transform 1 0 61344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_640
timestamp 1679581782
transform 1 0 62016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_647
timestamp 1679581782
transform 1 0 62688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_654
timestamp 1679581782
transform 1 0 63360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_661
timestamp 1679581782
transform 1 0 64032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_668
timestamp 1679581782
transform 1 0 64704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_675
timestamp 1679581782
transform 1 0 65376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_682
timestamp 1679581782
transform 1 0 66048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_689
timestamp 1679581782
transform 1 0 66720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_696
timestamp 1679581782
transform 1 0 67392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_703
timestamp 1679581782
transform 1 0 68064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_710
timestamp 1679581782
transform 1 0 68736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_717
timestamp 1679581782
transform 1 0 69408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_724
timestamp 1679581782
transform 1 0 70080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_731
timestamp 1679581782
transform 1 0 70752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_738
timestamp 1679581782
transform 1 0 71424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_745
timestamp 1679581782
transform 1 0 72096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_752
timestamp 1679581782
transform 1 0 72768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_759
timestamp 1679581782
transform 1 0 73440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_766
timestamp 1679581782
transform 1 0 74112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_773
timestamp 1679581782
transform 1 0 74784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_780
timestamp 1679581782
transform 1 0 75456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_787
timestamp 1679581782
transform 1 0 76128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_794
timestamp 1679581782
transform 1 0 76800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_801
timestamp 1679581782
transform 1 0 77472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_808
timestamp 1679581782
transform 1 0 78144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_815
timestamp 1679581782
transform 1 0 78816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_822
timestamp 1679581782
transform 1 0 79488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_829
timestamp 1679581782
transform 1 0 80160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_836
timestamp 1679581782
transform 1 0 80832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_843
timestamp 1679581782
transform 1 0 81504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_850
timestamp 1679581782
transform 1 0 82176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_857
timestamp 1679577901
transform 1 0 82848 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_861
timestamp 1677579658
transform 1 0 83232 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679581782
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679581782
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679581782
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_861
timestamp 1677579658
transform 1 0 83232 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679581782
transform 1 0 56352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679581782
transform 1 0 57024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679581782
transform 1 0 57696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679581782
transform 1 0 58368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679581782
transform 1 0 59040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679581782
transform 1 0 59712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679581782
transform 1 0 60384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679581782
transform 1 0 61056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679581782
transform 1 0 61728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679581782
transform 1 0 62400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679581782
transform 1 0 63744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679581782
transform 1 0 64416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679581782
transform 1 0 65088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679581782
transform 1 0 65760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679581782
transform 1 0 66432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679581782
transform 1 0 67104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679581782
transform 1 0 67776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679581782
transform 1 0 68448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679581782
transform 1 0 69120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679581782
transform 1 0 69792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679581782
transform 1 0 70464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679581782
transform 1 0 71136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679581782
transform 1 0 71808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679581782
transform 1 0 72480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679581782
transform 1 0 73152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679581782
transform 1 0 73824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679581782
transform 1 0 74496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679581782
transform 1 0 75168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679581782
transform 1 0 75840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679581782
transform 1 0 76512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679581782
transform 1 0 77184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679581782
transform 1 0 77856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679581782
transform 1 0 78528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679581782
transform 1 0 79200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679581782
transform 1 0 79872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679581782
transform 1 0 80544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_840
timestamp 1679581782
transform 1 0 81216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_847
timestamp 1679581782
transform 1 0 81888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_854
timestamp 1679581782
transform 1 0 82560 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_861
timestamp 1677579658
transform 1 0 83232 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679581782
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679581782
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679581782
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679581782
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679581782
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679581782
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679581782
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679581782
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679581782
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679581782
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679581782
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679581782
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679581782
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_214
timestamp 1679581782
transform 1 0 21120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_221
timestamp 1679581782
transform 1 0 21792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_228
timestamp 1679581782
transform 1 0 22464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_235
timestamp 1679581782
transform 1 0 23136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_242
timestamp 1679581782
transform 1 0 23808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_249
timestamp 1679581782
transform 1 0 24480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_256
timestamp 1679581782
transform 1 0 25152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_263
timestamp 1679581782
transform 1 0 25824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_270
timestamp 1679581782
transform 1 0 26496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_277
timestamp 1679581782
transform 1 0 27168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_284
timestamp 1679581782
transform 1 0 27840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_291
timestamp 1679581782
transform 1 0 28512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_298
timestamp 1679581782
transform 1 0 29184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_305
timestamp 1679581782
transform 1 0 29856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_312
timestamp 1679581782
transform 1 0 30528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_319
timestamp 1679581782
transform 1 0 31200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_326
timestamp 1679581782
transform 1 0 31872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_333
timestamp 1679581782
transform 1 0 32544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_340
timestamp 1679581782
transform 1 0 33216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_347
timestamp 1679581782
transform 1 0 33888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_354
timestamp 1679581782
transform 1 0 34560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_361
timestamp 1679581782
transform 1 0 35232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_368
timestamp 1679581782
transform 1 0 35904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_375
timestamp 1679581782
transform 1 0 36576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_382
timestamp 1679581782
transform 1 0 37248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_389
timestamp 1679581782
transform 1 0 37920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_396
timestamp 1679581782
transform 1 0 38592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679581782
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679581782
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_417
timestamp 1679581782
transform 1 0 40608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_424
timestamp 1679581782
transform 1 0 41280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_431
timestamp 1679581782
transform 1 0 41952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_438
timestamp 1679581782
transform 1 0 42624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_445
timestamp 1679581782
transform 1 0 43296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_452
timestamp 1679581782
transform 1 0 43968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_459
timestamp 1679581782
transform 1 0 44640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_466
timestamp 1679581782
transform 1 0 45312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_473
timestamp 1679581782
transform 1 0 45984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_480
timestamp 1679581782
transform 1 0 46656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_487
timestamp 1679581782
transform 1 0 47328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_494
timestamp 1679581782
transform 1 0 48000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_501
timestamp 1679581782
transform 1 0 48672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_508
timestamp 1679581782
transform 1 0 49344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_515
timestamp 1679581782
transform 1 0 50016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_522
timestamp 1679581782
transform 1 0 50688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_529
timestamp 1679581782
transform 1 0 51360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_536
timestamp 1679581782
transform 1 0 52032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_543
timestamp 1679581782
transform 1 0 52704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_550
timestamp 1679581782
transform 1 0 53376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_557
timestamp 1679581782
transform 1 0 54048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_564
timestamp 1679581782
transform 1 0 54720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_571
timestamp 1679581782
transform 1 0 55392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_578
timestamp 1679581782
transform 1 0 56064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_585
timestamp 1679581782
transform 1 0 56736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_592
timestamp 1679581782
transform 1 0 57408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_599
timestamp 1679581782
transform 1 0 58080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_606
timestamp 1679581782
transform 1 0 58752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_613
timestamp 1679581782
transform 1 0 59424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_620
timestamp 1679581782
transform 1 0 60096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_627
timestamp 1679581782
transform 1 0 60768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_634
timestamp 1679581782
transform 1 0 61440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_641
timestamp 1679581782
transform 1 0 62112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_648
timestamp 1679581782
transform 1 0 62784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_655
timestamp 1679581782
transform 1 0 63456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_662
timestamp 1679581782
transform 1 0 64128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_669
timestamp 1679581782
transform 1 0 64800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_676
timestamp 1679581782
transform 1 0 65472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_683
timestamp 1679581782
transform 1 0 66144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_690
timestamp 1679581782
transform 1 0 66816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_697
timestamp 1679581782
transform 1 0 67488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_704
timestamp 1679581782
transform 1 0 68160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_711
timestamp 1679581782
transform 1 0 68832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_718
timestamp 1679581782
transform 1 0 69504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_725
timestamp 1679581782
transform 1 0 70176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_732
timestamp 1679581782
transform 1 0 70848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_739
timestamp 1679581782
transform 1 0 71520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_746
timestamp 1679581782
transform 1 0 72192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_753
timestamp 1679581782
transform 1 0 72864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_760
timestamp 1679581782
transform 1 0 73536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_767
timestamp 1679581782
transform 1 0 74208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_774
timestamp 1679581782
transform 1 0 74880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_781
timestamp 1679581782
transform 1 0 75552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_788
timestamp 1679581782
transform 1 0 76224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_795
timestamp 1679581782
transform 1 0 76896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_802
timestamp 1679581782
transform 1 0 77568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_809
timestamp 1679581782
transform 1 0 78240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_816
timestamp 1679581782
transform 1 0 78912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_823
timestamp 1679581782
transform 1 0 79584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_830
timestamp 1679581782
transform 1 0 80256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_837
timestamp 1679581782
transform 1 0 80928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_844
timestamp 1679581782
transform 1 0 81600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_851
timestamp 1679581782
transform 1 0 82272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_858
timestamp 1679577901
transform 1 0 82944 0 -1 38556
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_43
timestamp 1680000637
transform -1 0 1344 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_44
timestamp 1680000637
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_45
timestamp 1680000637
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_46
timestamp 1680000637
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_47
timestamp 1680000637
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_48
timestamp 1680000637
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_49
timestamp 1680000637
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tielo  heichips25_template
timestamp 1680000637
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_50
timestamp 1680000637
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_51
timestamp 1680000637
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_52
timestamp 1680000637
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_53
timestamp 1680000637
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_54
timestamp 1680000637
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_55
timestamp 1680000637
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_56
timestamp 1680000637
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_57
timestamp 1680000637
transform -1 0 1344 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 960 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 1344 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform -1 0 960 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use adc  u_adc
timestamp 0
transform 1 0 84000 0 1 1000
box 0 0 1 1
use delay_line  u_delay_line
timestamp 0
transform 1 0 85400 0 1 24200
box 0 0 1 1
use multimode_dll  u_multimode_dll
timestamp 0
transform 1 0 8000 0 1 6000
box 0 0 1 1
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 712 95476 38600 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via5 65100 22800 65100 22800 0 VGND
rlabel via5 63860 27560 63860 27560 0 VPWR
rlabel metal3 1152 26208 1152 26208 0 _000_
rlabel metal2 768 28602 768 28602 0 _001_
rlabel metal3 2112 29946 2112 29946 0 _002_
rlabel metal2 3504 29316 3504 29316 0 _003_
rlabel metal3 5280 27048 5280 27048 0 _004_
rlabel metal3 3792 24444 3792 24444 0 _005_
rlabel metal2 2880 24003 2880 24003 0 _006_
rlabel metal2 2400 30660 2400 30660 0 _007_
rlabel metal2 27168 33390 27168 33390 0 _008_
rlabel metal2 29280 32844 29280 32844 0 _009_
rlabel metal2 31104 33600 31104 33600 0 _010_
rlabel metal3 34896 33684 34896 33684 0 _011_
rlabel metal2 41664 33390 41664 33390 0 _012_
rlabel metal3 50160 33768 50160 33768 0 _013_
rlabel metal2 52224 33822 52224 33822 0 _014_
rlabel metal2 47520 33402 47520 33402 0 _015_
rlabel metal2 44928 33402 44928 33402 0 _016_
rlabel metal2 37920 33978 37920 33978 0 _017_
rlabel metal2 32352 34650 32352 34650 0 _018_
rlabel metal2 34368 33894 34368 33894 0 _019_
rlabel metal2 32832 2898 32832 2898 0 _020_
rlabel metal2 35808 2688 35808 2688 0 _021_
rlabel metal2 46752 2898 46752 2898 0 _022_
rlabel metal2 49632 2898 49632 2898 0 _023_
rlabel metal2 52800 2898 52800 2898 0 _024_
rlabel metal2 55344 2604 55344 2604 0 _025_
rlabel metal2 55104 1890 55104 1890 0 _026_
rlabel metal2 52512 1890 52512 1890 0 _027_
rlabel metal2 49920 1638 49920 1638 0 _028_
rlabel metal2 47328 1638 47328 1638 0 _029_
rlabel metal2 38976 2898 38976 2898 0 _030_
rlabel metal2 37680 1932 37680 1932 0 _031_
rlabel metal2 37248 1890 37248 1890 0 _032_
rlabel metal2 32160 1848 32160 1848 0 _033_
rlabel metal2 30336 1176 30336 1176 0 _034_
rlabel metal2 28800 2898 28800 2898 0 _035_
rlabel metal2 27744 1848 27744 1848 0 _036_
rlabel metal2 21024 1638 21024 1638 0 _037_
rlabel metal2 20112 2604 20112 2604 0 _038_
rlabel metal2 22656 3360 22656 3360 0 _039_
rlabel metal2 22656 1386 22656 1386 0 _040_
rlabel metal2 24096 1848 24096 1848 0 _041_
rlabel metal2 26016 2688 26016 2688 0 _042_
rlabel metal2 40512 1176 40512 1176 0 _043_
rlabel metal2 44544 1848 44544 1848 0 _044_
rlabel metal2 45696 2688 45696 2688 0 _045_
rlabel metal2 4224 15582 4224 15582 0 _046_
rlabel metal2 3504 18564 3504 18564 0 _047_
rlabel metal2 3456 20034 3456 20034 0 _048_
rlabel metal2 9888 32928 9888 32928 0 _049_
rlabel metal2 14016 33390 14016 33390 0 _050_
rlabel metal2 17712 33516 17712 33516 0 _051_
rlabel metal2 15408 34272 15408 34272 0 _052_
rlabel metal2 3888 21420 3888 21420 0 _053_
rlabel metal2 3552 7686 3552 7686 0 _054_
rlabel metal2 2880 8736 2880 8736 0 _055_
rlabel metal2 1536 9702 1536 9702 0 _056_
rlabel metal2 1344 12222 1344 12222 0 _057_
rlabel metal2 1200 13860 1200 13860 0 _058_
rlabel metal2 2016 16758 2016 16758 0 _059_
rlabel metal3 1248 18564 1248 18564 0 _060_
rlabel metal2 2496 20286 2496 20286 0 _061_
rlabel metal2 5280 32760 5280 32760 0 _062_
rlabel metal2 18144 32928 18144 32928 0 _063_
rlabel metal2 21360 32844 21360 32844 0 _064_
rlabel metal2 25344 34146 25344 34146 0 _065_
rlabel metal2 16896 3150 16896 3150 0 _066_
rlabel metal2 13824 3360 13824 3360 0 _067_
rlabel metal2 4224 4872 4224 4872 0 _068_
rlabel metal2 4032 9408 4032 9408 0 _069_
rlabel metal3 3600 10836 3600 10836 0 _070_
rlabel metal3 3696 12348 3696 12348 0 _071_
rlabel metal2 3648 14238 3648 14238 0 _072_
rlabel metal2 76800 13272 76800 13272 0 _073_
rlabel metal2 79488 11970 79488 11970 0 _074_
rlabel metal2 79968 12516 79968 12516 0 _075_
rlabel metal2 79488 10458 79488 10458 0 _076_
rlabel metal2 79488 4410 79488 4410 0 _077_
rlabel metal2 79488 1848 79488 1848 0 _078_
rlabel metal2 79536 2520 79536 2520 0 _079_
rlabel metal3 79824 6468 79824 6468 0 _080_
rlabel metal2 79488 15246 79488 15246 0 _081_
rlabel metal2 81888 19992 81888 19992 0 _082_
rlabel metal3 81120 27636 81120 27636 0 _083_
rlabel metal3 81120 32172 81120 32172 0 _084_
rlabel metal3 81216 33516 81216 33516 0 _085_
rlabel metal3 1008 23100 1008 23100 0 _086_
rlabel metal2 4464 28140 4464 28140 0 _087_
rlabel metal2 4272 24780 4272 24780 0 _088_
rlabel metal3 3312 5124 3312 5124 0 _089_
rlabel metal3 2064 11844 2064 11844 0 _090_
rlabel metal2 1440 5376 1440 5376 0 _091_
rlabel metal2 1728 5418 1728 5418 0 _092_
rlabel metal2 2016 5208 2016 5208 0 _093_
rlabel metal3 4320 13020 4320 13020 0 _094_
rlabel metal3 1920 15540 1920 15540 0 _095_
rlabel metal3 4320 14448 4320 14448 0 _096_
rlabel metal2 1920 24906 1920 24906 0 _097_
rlabel metal3 5520 23016 5520 23016 0 _098_
rlabel metal3 4896 25914 4896 25914 0 _099_
rlabel metal2 2592 26376 2592 26376 0 _100_
rlabel metal2 3744 28602 3744 28602 0 _101_
rlabel metal2 2016 25620 2016 25620 0 _102_
rlabel metal2 1824 23980 1824 23980 0 _103_
rlabel metal2 1728 26166 1728 26166 0 _104_
rlabel metal2 3648 27132 3648 27132 0 _105_
rlabel metal2 1776 29148 1776 29148 0 _106_
rlabel metal2 1584 29148 1584 29148 0 _107_
rlabel metal2 2688 29274 2688 29274 0 _108_
rlabel metal2 2304 29820 2304 29820 0 _109_
rlabel metal3 3792 28476 3792 28476 0 _110_
rlabel metal2 3840 26250 3840 26250 0 _111_
rlabel metal2 4512 26712 4512 26712 0 _112_
rlabel metal2 4656 26796 4656 26796 0 _113_
rlabel metal2 3936 25284 3936 25284 0 _114_
rlabel metal2 4128 25242 4128 25242 0 _115_
rlabel metal4 1728 7056 1728 7056 0 adc_data\[0\]
rlabel metal3 1776 11172 1776 11172 0 adc_data\[1\]
rlabel metal2 1296 8400 1296 8400 0 adc_data\[2\]
rlabel metal4 99960 6160 99960 6160 0 adc_data\[3\]
rlabel metal2 30816 2058 30816 2058 0 adc_data\[4\]
rlabel metal2 89280 920 89280 920 0 adc_data\[5\]
rlabel metal4 73056 6972 73056 6972 0 adc_data\[6\]
rlabel metal4 99960 11326 99960 11326 0 adc_data\[7\]
rlabel metal3 2910 36708 2910 36708 0 clk
rlabel metal2 40717 5866 40717 5866 0 clk0_out
rlabel metal2 37453 5866 37453 5866 0 clk1_out
rlabel metal2 37680 5814 37680 5814 0 clk2_out
rlabel metal3 3984 21504 3984 21504 0 clk_delayed
rlabel metal2 65952 33012 65952 33012 0 clk_regs
rlabel metal2 79776 23688 79776 23688 0 clknet_0_clk
rlabel metal2 21792 33852 21792 33852 0 clknet_0_clk_regs
rlabel metal4 26880 5964 26880 5964 0 clknet_1_0__leaf_clk
rlabel metal3 89664 24528 89664 24528 0 clknet_1_1__leaf_clk
rlabel metal2 4704 18648 4704 18648 0 clknet_4_0_0_clk_regs
rlabel metal2 44448 2310 44448 2310 0 clknet_4_10_0_clk_regs
rlabel metal3 41040 33684 41040 33684 0 clknet_4_11_0_clk_regs
rlabel metal2 80736 4956 80736 4956 0 clknet_4_12_0_clk_regs
rlabel metal2 46080 2310 46080 2310 0 clknet_4_13_0_clk_regs
rlabel metal3 79392 13188 79392 13188 0 clknet_4_14_0_clk_regs
rlabel metal3 81936 20076 81936 20076 0 clknet_4_15_0_clk_regs
rlabel metal2 4128 20748 4128 20748 0 clknet_4_1_0_clk_regs
rlabel metal2 4752 5628 4752 5628 0 clknet_4_2_0_clk_regs
rlabel metal3 4752 13188 4752 13188 0 clknet_4_3_0_clk_regs
rlabel metal2 2064 26124 2064 26124 0 clknet_4_4_0_clk_regs
rlabel metal2 2496 30786 2496 30786 0 clknet_4_5_0_clk_regs
rlabel metal2 24096 33726 24096 33726 0 clknet_4_6_0_clk_regs
rlabel metal2 26592 33558 26592 33558 0 clknet_4_7_0_clk_regs
rlabel metal3 25584 2604 25584 2604 0 clknet_4_8_0_clk_regs
rlabel metal3 24624 1092 24624 1092 0 clknet_4_9_0_clk_regs
rlabel metal2 1536 30282 1536 30282 0 data\[0\]
rlabel metal2 38496 34062 38496 34062 0 data\[10\]
rlabel metal2 32640 35112 32640 35112 0 data\[11\]
rlabel metal2 34224 35196 34224 35196 0 data\[12\]
rlabel metal2 34944 3528 34944 3528 0 data\[13\]
rlabel metal2 46368 3234 46368 3234 0 data\[14\]
rlabel metal3 46464 3570 46464 3570 0 data\[15\]
rlabel metal2 47328 4704 47328 4704 0 data\[16\]
rlabel metal2 46944 4578 46944 4578 0 data\[17\]
rlabel metal2 47136 4662 47136 4662 0 data\[18\]
rlabel metal2 47424 3444 47424 3444 0 data\[19\]
rlabel metal2 29616 33432 29616 33432 0 data\[1\]
rlabel metal2 47232 1260 47232 1260 0 data\[20\]
rlabel metal2 44736 1050 44736 1050 0 data\[21\]
rlabel metal2 44928 2856 44928 2856 0 data\[22\]
rlabel metal3 38640 2856 38640 2856 0 data\[23\]
rlabel metal2 40032 2100 40032 2100 0 data\[24\]
rlabel metal2 34848 2058 34848 2058 0 data\[25\]
rlabel metal2 34512 2100 34512 2100 0 data\[26\]
rlabel metal3 34032 1344 34032 1344 0 data\[27\]
rlabel metal2 27168 2394 27168 2394 0 data\[28\]
rlabel metal2 27264 1890 27264 1890 0 data\[29\]
rlabel metal2 31776 31500 31776 31500 0 data\[2\]
rlabel metal2 20448 4578 20448 4578 0 data\[30\]
rlabel metal2 22080 3612 22080 3612 0 data\[31\]
rlabel metal2 22176 3738 22176 3738 0 data\[32\]
rlabel metal2 23424 2184 23424 2184 0 data\[33\]
rlabel metal2 23520 3864 23520 3864 0 data\[34\]
rlabel metal2 39888 1092 39888 1092 0 data\[35\]
rlabel metal2 40032 1470 40032 1470 0 data\[36\]
rlabel metal2 41664 2100 41664 2100 0 data\[37\]
rlabel metal2 42816 2646 42816 2646 0 data\[38\]
rlabel metal3 5376 17304 5376 17304 0 data\[39\]
rlabel metal3 31104 33684 31104 33684 0 data\[3\]
rlabel metal2 5856 17934 5856 17934 0 data\[40\]
rlabel metal3 5952 19992 5952 19992 0 data\[41\]
rlabel metal2 14112 32760 14112 32760 0 data\[42\]
rlabel metal4 17472 32886 17472 32886 0 data\[43\]
rlabel metal2 20448 33852 20448 33852 0 data\[44\]
rlabel metal3 4704 21588 4704 21588 0 data\[45\]
rlabel metal2 5904 22092 5904 22092 0 data\[46\]
rlabel metal3 4896 7140 4896 7140 0 data\[47\]
rlabel metal2 5280 9996 5280 9996 0 data\[48\]
rlabel metal2 3264 10206 3264 10206 0 data\[49\]
rlabel metal3 39312 33432 39312 33432 0 data\[4\]
rlabel metal2 3744 12222 3744 12222 0 data\[50\]
rlabel metal2 3408 14952 3408 14952 0 data\[51\]
rlabel metal2 2016 17502 2016 17502 0 data\[52\]
rlabel metal3 3648 18312 3648 18312 0 data\[53\]
rlabel metal2 5232 21000 5232 21000 0 data\[54\]
rlabel metal2 17568 32676 17568 32676 0 data\[55\]
rlabel metal3 20784 33096 20784 33096 0 data\[56\]
rlabel metal2 23712 31500 23712 31500 0 data\[57\]
rlabel metal2 18253 30026 18253 30026 0 data\[58\]
rlabel metal2 19296 3696 19296 3696 0 data\[59\]
rlabel metal2 49296 33516 49296 33516 0 data\[5\]
rlabel metal2 4608 4536 4608 4536 0 data\[60\]
rlabel metal3 5424 5712 5424 5712 0 data\[61\]
rlabel metal2 5856 10668 5856 10668 0 data\[62\]
rlabel metal2 5856 11550 5856 11550 0 data\[63\]
rlabel metal2 5904 13440 5904 13440 0 data\[64\]
rlabel metal2 5856 14322 5856 14322 0 data\[65\]
rlabel metal2 79392 12432 79392 12432 0 data\[66\]
rlabel metal2 81888 11634 81888 11634 0 data\[67\]
rlabel metal2 81936 13440 81936 13440 0 data\[68\]
rlabel metal2 80400 6048 80400 6048 0 data\[69\]
rlabel metal3 51840 34314 51840 34314 0 data\[6\]
rlabel metal2 81984 3948 81984 3948 0 data\[70\]
rlabel metal2 81888 1218 81888 1218 0 data\[71\]
rlabel metal2 81936 2436 81936 2436 0 data\[72\]
rlabel metal2 81888 6048 81888 6048 0 data\[73\]
rlabel metal2 81360 19488 81360 19488 0 data\[74\]
rlabel metal2 81408 22428 81408 22428 0 data\[75\]
rlabel metal2 81696 27078 81696 27078 0 data\[76\]
rlabel metal3 84316 32004 84316 32004 0 data\[77\]
rlabel metal2 83232 35364 83232 35364 0 data\[78\]
rlabel metal2 54336 32550 54336 32550 0 data\[7\]
rlabel metal2 49632 33432 49632 33432 0 data\[8\]
rlabel metal2 38592 33768 38592 33768 0 data\[9\]
rlabel metal2 38784 31656 38784 31656 0 delaynet_0_clk
rlabel metal2 25728 5628 25728 5628 0 ena
rlabel metal3 366 15708 366 15708 0 net
rlabel metal3 1392 32088 1392 32088 0 net1
rlabel metal3 1296 7140 1296 7140 0 net10
rlabel metal3 1248 7056 1248 7056 0 net11
rlabel metal2 1920 13524 1920 13524 0 net12
rlabel metal3 1488 15456 1488 15456 0 net13
rlabel metal2 2304 16128 2304 16128 0 net14
rlabel metal2 4224 7098 4224 7098 0 net15
rlabel metal2 1440 17724 1440 17724 0 net16
rlabel metal3 3984 20076 3984 20076 0 net17
rlabel metal2 20688 33600 20688 33600 0 net18
rlabel metal2 26880 2310 26880 2310 0 net19
rlabel metal2 864 23730 864 23730 0 net2
rlabel metal2 38304 1134 38304 1134 0 net20
rlabel metal2 22080 34272 22080 34272 0 net21
rlabel metal2 21312 3192 21312 3192 0 net22
rlabel metal3 4512 22848 4512 22848 0 net23
rlabel metal2 42384 2604 42384 2604 0 net24
rlabel metal4 63360 4116 63360 4116 0 net25
rlabel metal2 80256 1344 80256 1344 0 net26
rlabel metal2 81024 20874 81024 20874 0 net27
rlabel metal2 3840 10248 3840 10248 0 net28
rlabel metal2 3792 5628 3792 5628 0 net29
rlabel metal2 912 24780 912 24780 0 net3
rlabel metal2 3264 17766 3264 17766 0 net30
rlabel metal3 1152 26124 1152 26124 0 net31
rlabel metal2 1104 26880 1104 26880 0 net32
rlabel metal2 1728 32298 1728 32298 0 net33
rlabel metal2 26400 4116 26400 4116 0 net34
rlabel metal2 39360 2562 39360 2562 0 net35
rlabel metal2 24960 33768 24960 33768 0 net36
rlabel metal2 23424 2898 23424 2898 0 net37
rlabel metal2 45312 2562 45312 2562 0 net38
rlabel metal2 45216 2730 45216 2730 0 net39
rlabel metal2 1392 20832 1392 20832 0 net4
rlabel metal2 79920 4116 79920 4116 0 net40
rlabel metal2 82272 20118 82272 20118 0 net41
rlabel metal2 2736 26964 2736 26964 0 net42
rlabel metal3 558 16548 558 16548 0 net43
rlabel metal3 366 17388 366 17388 0 net44
rlabel metal3 366 18228 366 18228 0 net45
rlabel metal3 366 19068 366 19068 0 net46
rlabel metal3 366 19908 366 19908 0 net47
rlabel metal3 366 20748 366 20748 0 net48
rlabel metal3 366 21588 366 21588 0 net49
rlabel metal2 624 24696 624 24696 0 net5
rlabel metal3 366 2268 366 2268 0 net50
rlabel metal3 366 3108 366 3108 0 net51
rlabel metal3 366 3948 366 3948 0 net52
rlabel metal3 366 4788 366 4788 0 net53
rlabel metal3 366 5628 366 5628 0 net54
rlabel metal3 366 6468 366 6468 0 net55
rlabel metal3 366 7308 366 7308 0 net56
rlabel metal3 558 8148 558 8148 0 net57
rlabel metal2 864 8778 864 8778 0 net6
rlabel metal2 912 9408 912 9408 0 net7
rlabel metal2 1104 9660 1104 9660 0 net8
rlabel metal2 1392 8316 1392 8316 0 net9
rlabel metal2 31728 5856 31728 5856 0 osc_out
rlabel metal3 366 37548 366 37548 0 rst_n
rlabel metal2 34765 5866 34765 5866 0 stable
rlabel metal2 1536 26040 1536 26040 0 u_shift_reg.bit_count\[0\]
rlabel metal2 2016 28938 2016 28938 0 u_shift_reg.bit_count\[1\]
rlabel metal2 2688 29778 2688 29778 0 u_shift_reg.bit_count\[2\]
rlabel metal3 4896 29148 4896 29148 0 u_shift_reg.bit_count\[3\]
rlabel metal2 4320 26754 4320 26754 0 u_shift_reg.bit_count\[4\]
rlabel metal2 4512 25620 4512 25620 0 u_shift_reg.bit_count\[5\]
rlabel metal2 3744 24570 3744 24570 0 u_shift_reg.bit_count\[6\]
rlabel metal2 2016 23520 2016 23520 0 u_shift_reg.locked
rlabel metal3 558 22428 558 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 558 24108 558 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal2 672 8946 672 8946 0 uio_out[0]
rlabel metal2 672 9744 672 9744 0 uio_out[1]
rlabel metal3 558 10668 558 10668 0 uio_out[2]
rlabel metal2 624 11172 624 11172 0 uio_out[3]
rlabel metal2 672 12138 672 12138 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 366 14028 366 14028 0 uio_out[6]
rlabel metal3 366 14868 366 14868 0 uio_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
