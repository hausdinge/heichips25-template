module heichips25_template (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net1;
 wire net2;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;

 sg13g2_inv_1 _31_ (.VDD(VPWR),
    .Y(_08_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _32_ (.VDD(VPWR),
    .Y(_09_),
    .A(net1),
    .VSS(VGND));
 sg13g2_and3_1 _33_ (.X(_10_),
    .A(net2),
    .B(net34),
    .C(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _34_ (.X(_11_),
    .A(net44),
    .B(net41),
    .C(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _35_ (.A(_10_),
    .B(_11_),
    .X(_12_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _36_ (.B1(net1),
    .VDD(VPWR),
    .Y(_13_),
    .VSS(VGND),
    .A1(net46),
    .A2(_12_));
 sg13g2_a21oi_1 _37_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net46),
    .A2(_12_),
    .Y(_00_),
    .B1(_13_));
 sg13g2_a21oi_1 _38_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net8),
    .A2(_12_),
    .Y(_14_),
    .B1(net38));
 sg13g2_and4_1 _39_ (.A(net38),
    .B(net8),
    .C(_10_),
    .D(_11_),
    .X(_15_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _40_ (.A(_09_),
    .B(net39),
    .C(_15_),
    .Y(_01_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _41_ (.B1(net1),
    .VDD(VPWR),
    .Y(_16_),
    .VSS(VGND),
    .A1(net36),
    .A2(_15_));
 sg13g2_a21oi_1 _42_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net36),
    .A2(_15_),
    .Y(_02_),
    .B1(_16_));
 sg13g2_o21ai_1 _43_ (.B1(net1),
    .VDD(VPWR),
    .Y(_17_),
    .VSS(VGND),
    .A1(net2),
    .A2(net47));
 sg13g2_a21oi_1 _44_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2),
    .A2(net47),
    .Y(_03_),
    .B1(_17_));
 sg13g2_a21oi_1 _45_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2),
    .A2(net3),
    .Y(_18_),
    .B1(net34));
 sg13g2_nor3_1 _46_ (.A(_09_),
    .B(_10_),
    .C(net35),
    .Y(_04_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _47_ (.B1(net1),
    .VDD(VPWR),
    .Y(_19_),
    .VSS(VGND),
    .A1(net48),
    .A2(_10_));
 sg13g2_a21oi_1 _48_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net48),
    .A2(_10_),
    .Y(_05_),
    .B1(_19_));
 sg13g2_a21oi_1 _49_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net5),
    .A2(_10_),
    .Y(_20_),
    .B1(net41));
 sg13g2_nand3_1 _50_ (.B(net5),
    .C(_10_),
    .A(net41),
    .Y(_21_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _51_ (.Y(_22_),
    .A(net1),
    .B(_21_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _52_ (.A(net42),
    .B(_22_),
    .Y(_06_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _53_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_08_),
    .C1(_09_),
    .B1(_21_),
    .A1(_10_),
    .Y(_07_),
    .A2(_11_));
 sg13g2_dfrbpq_1 _54_ (.RESET_B(net25),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00_),
    .Q(net8),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _55_ (.RESET_B(net24),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net40),
    .Q(net9),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _56_ (.RESET_B(net22),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net37),
    .Q(net10),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _57_ (.RESET_B(net20),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_03_),
    .Q(net3),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _58_ (.RESET_B(net),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_04_),
    .Q(net4),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_1 _59_ (.RESET_B(net23),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_05_),
    .Q(net5),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _60_ (.RESET_B(net19),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net43),
    .Q(net6),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_1 _61_ (.RESET_B(net21),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net45),
    .Q(net7),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_tiehi _60__20 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net19));
 sg13g2_tiehi _57__21 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net20));
 sg13g2_tiehi _61__22 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net21));
 sg13g2_tiehi _56__23 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net22));
 sg13g2_tiehi _59__24 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net23));
 sg13g2_tiehi _55__25 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net24));
 sg13g2_tiehi _54__26 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net25));
 sg13g2_tiehi heichips25_template (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net26));
 sg13g2_tiehi heichips25_template_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net27));
 sg13g2_tiehi heichips25_template_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net28));
 sg13g2_tiehi heichips25_template_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net29));
 sg13g2_tiehi heichips25_template_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net30));
 sg13g2_tiehi heichips25_template_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net31));
 sg13g2_tiehi heichips25_template_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net32));
 sg13g2_tiehi heichips25_template_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _78_ (.A(net3),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _79_ (.A(net4),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _80_ (.A(net5),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _81_ (.A(net6),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _82_ (.A(net7),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _83_ (.A(net8),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _84_ (.A(net9),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _85_ (.A(net10),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _58__19 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net));
 sg13g2_buf_16 clkbuf_1_0__f_clk (.X(clknet_1_0__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_1_1__f_clk (.X(clknet_1_1__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold34 (.A(net4),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold35 (.A(_18_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold36 (.A(net10),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold37 (.A(_02_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold38 (.A(net9),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold39 (.A(_14_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold40 (.A(_01_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold41 (.A(net6),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold42 (.A(_20_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold43 (.A(_06_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold44 (.A(net7),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold45 (.A(_07_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold46 (.A(net8),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold47 (.A(net3),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold48 (.A(net5),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net26;
 assign uio_oe[1] = net27;
 assign uio_oe[2] = net28;
 assign uio_oe[3] = net29;
 assign uio_oe[4] = net30;
 assign uio_oe[5] = net31;
 assign uio_oe[6] = net32;
 assign uio_oe[7] = net33;
endmodule
