magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771805714
<< metal1 >>
rect 576 38576 83328 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 83328 38576
rect 576 38512 83328 38536
rect 22051 38408 22109 38409
rect 22051 38368 22060 38408
rect 22100 38368 22109 38408
rect 22051 38367 22109 38368
rect 26571 38408 26613 38417
rect 26571 38368 26572 38408
rect 26612 38368 26613 38408
rect 26571 38359 26613 38368
rect 27523 38408 27581 38409
rect 27523 38368 27532 38408
rect 27572 38368 27581 38408
rect 27523 38367 27581 38368
rect 27619 38324 27677 38325
rect 27619 38284 27628 38324
rect 27668 38284 27677 38324
rect 27619 38283 27677 38284
rect 29443 38324 29501 38325
rect 29443 38284 29452 38324
rect 29492 38284 29501 38324
rect 29443 38283 29501 38284
rect 33675 38324 33717 38333
rect 33675 38284 33676 38324
rect 33716 38284 33717 38324
rect 33675 38275 33717 38284
rect 21955 38240 22013 38241
rect 21955 38200 21964 38240
rect 22004 38200 22013 38240
rect 21955 38199 22013 38200
rect 25987 38240 26045 38241
rect 25987 38200 25996 38240
rect 26036 38200 26045 38240
rect 25987 38199 26045 38200
rect 26475 38240 26517 38249
rect 26475 38200 26476 38240
rect 26516 38200 26517 38240
rect 26475 38191 26517 38200
rect 26667 38240 26709 38249
rect 26667 38200 26668 38240
rect 26708 38200 26709 38240
rect 26667 38191 26709 38200
rect 27723 38240 27765 38249
rect 27723 38200 27724 38240
rect 27764 38200 27765 38240
rect 27723 38191 27765 38200
rect 27819 38240 27861 38249
rect 27819 38200 27820 38240
rect 27860 38200 27861 38240
rect 27819 38191 27861 38200
rect 28963 38240 29021 38241
rect 28963 38200 28972 38240
rect 29012 38200 29021 38240
rect 28963 38199 29021 38200
rect 29251 38240 29309 38241
rect 29251 38200 29260 38240
rect 29300 38200 29309 38240
rect 29251 38199 29309 38200
rect 29739 38240 29781 38249
rect 29739 38200 29740 38240
rect 29780 38200 29781 38240
rect 29739 38191 29781 38200
rect 29923 38240 29981 38241
rect 29923 38200 29932 38240
rect 29972 38200 29981 38240
rect 29923 38199 29981 38200
rect 33283 38240 33341 38241
rect 33283 38200 33292 38240
rect 33332 38200 33341 38240
rect 33283 38199 33341 38200
rect 33579 38240 33621 38249
rect 33579 38200 33580 38240
rect 33620 38200 33621 38240
rect 33579 38191 33621 38200
rect 37515 38240 37557 38249
rect 37515 38200 37516 38240
rect 37556 38200 37557 38240
rect 37411 38198 37469 38199
rect 37411 38158 37420 38198
rect 37460 38158 37469 38198
rect 37515 38191 37557 38200
rect 37795 38240 37853 38241
rect 37795 38200 37804 38240
rect 37844 38200 37853 38240
rect 37795 38199 37853 38200
rect 37411 38157 37469 38158
rect 643 38156 701 38157
rect 643 38116 652 38156
rect 692 38116 701 38156
rect 643 38115 701 38116
rect 22723 38156 22781 38157
rect 22723 38116 22732 38156
rect 22772 38116 22781 38156
rect 22723 38115 22781 38116
rect 23683 38156 23741 38157
rect 23683 38116 23692 38156
rect 23732 38116 23741 38156
rect 23683 38115 23741 38116
rect 24259 38156 24317 38157
rect 24259 38116 24268 38156
rect 24308 38116 24317 38156
rect 24259 38115 24317 38116
rect 24643 38156 24701 38157
rect 24643 38116 24652 38156
rect 24692 38116 24701 38156
rect 24643 38115 24701 38116
rect 24459 38072 24501 38081
rect 24459 38032 24460 38072
rect 24500 38032 24501 38072
rect 24459 38023 24501 38032
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 21763 37988 21821 37989
rect 21763 37948 21772 37988
rect 21812 37948 21821 37988
rect 21763 37947 21821 37948
rect 22539 37988 22581 37997
rect 22539 37948 22540 37988
rect 22580 37948 22581 37988
rect 22539 37939 22581 37948
rect 23883 37988 23925 37997
rect 23883 37948 23884 37988
rect 23924 37948 23925 37988
rect 23883 37939 23925 37948
rect 24075 37988 24117 37997
rect 24075 37948 24076 37988
rect 24116 37948 24117 37988
rect 24075 37939 24117 37948
rect 26091 37988 26133 37997
rect 26091 37948 26092 37988
rect 26132 37948 26133 37988
rect 26091 37939 26133 37948
rect 27531 37988 27573 37997
rect 27531 37948 27532 37988
rect 27572 37948 27573 37988
rect 27531 37939 27573 37948
rect 29835 37988 29877 37997
rect 29835 37948 29836 37988
rect 29876 37948 29877 37988
rect 29835 37939 29877 37948
rect 33955 37988 34013 37989
rect 33955 37948 33964 37988
rect 34004 37948 34013 37988
rect 33955 37947 34013 37948
rect 37123 37988 37181 37989
rect 37123 37948 37132 37988
rect 37172 37948 37181 37988
rect 37123 37947 37181 37948
rect 576 37820 83328 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 83328 37820
rect 576 37756 83328 37780
rect 26667 37652 26709 37661
rect 26667 37612 26668 37652
rect 26708 37612 26709 37652
rect 26667 37603 26709 37612
rect 19747 37484 19805 37485
rect 19747 37444 19756 37484
rect 19796 37444 19805 37484
rect 19747 37443 19805 37444
rect 32899 37484 32957 37485
rect 32899 37444 32908 37484
rect 32948 37444 32957 37484
rect 32899 37443 32957 37444
rect 20619 37400 20661 37409
rect 20619 37360 20620 37400
rect 20660 37360 20661 37400
rect 20619 37351 20661 37360
rect 20715 37400 20757 37409
rect 20715 37360 20716 37400
rect 20756 37360 20757 37400
rect 20715 37351 20757 37360
rect 21003 37400 21045 37409
rect 21003 37360 21004 37400
rect 21044 37360 21045 37400
rect 21003 37351 21045 37360
rect 21379 37400 21437 37401
rect 21379 37360 21388 37400
rect 21428 37360 21437 37400
rect 21379 37359 21437 37360
rect 22243 37400 22301 37401
rect 22243 37360 22252 37400
rect 22292 37360 22301 37400
rect 22243 37359 22301 37360
rect 23971 37400 24029 37401
rect 23971 37360 23980 37400
rect 24020 37360 24029 37400
rect 23971 37359 24029 37360
rect 24835 37400 24893 37401
rect 24835 37360 24844 37400
rect 24884 37360 24893 37400
rect 24835 37359 24893 37360
rect 26371 37400 26429 37401
rect 26371 37360 26380 37400
rect 26420 37360 26429 37400
rect 26371 37359 26429 37360
rect 26475 37400 26517 37409
rect 26475 37360 26476 37400
rect 26516 37360 26517 37400
rect 26475 37351 26517 37360
rect 26667 37400 26709 37409
rect 26667 37360 26668 37400
rect 26708 37360 26709 37400
rect 26667 37351 26709 37360
rect 26859 37400 26901 37409
rect 26859 37360 26860 37400
rect 26900 37360 26901 37400
rect 26859 37351 26901 37360
rect 27235 37400 27293 37401
rect 27235 37360 27244 37400
rect 27284 37360 27293 37400
rect 27235 37359 27293 37360
rect 28099 37400 28157 37401
rect 28099 37360 28108 37400
rect 28148 37360 28157 37400
rect 28099 37359 28157 37360
rect 29731 37400 29789 37401
rect 29731 37360 29740 37400
rect 29780 37360 29789 37400
rect 29731 37359 29789 37360
rect 29827 37400 29885 37401
rect 29827 37360 29836 37400
rect 29876 37360 29885 37400
rect 29827 37359 29885 37360
rect 30595 37400 30653 37401
rect 30595 37360 30604 37400
rect 30644 37360 30653 37400
rect 30595 37359 30653 37360
rect 31459 37400 31517 37401
rect 31459 37360 31468 37400
rect 31508 37360 31517 37400
rect 31459 37359 31517 37360
rect 34435 37400 34493 37401
rect 34435 37360 34444 37400
rect 34484 37360 34493 37400
rect 34435 37359 34493 37360
rect 35299 37400 35357 37401
rect 35299 37360 35308 37400
rect 35348 37360 35357 37400
rect 35299 37359 35357 37360
rect 35691 37400 35733 37409
rect 35691 37360 35692 37400
rect 35732 37360 35733 37400
rect 35691 37351 35733 37360
rect 36651 37400 36693 37409
rect 36651 37360 36652 37400
rect 36692 37360 36693 37400
rect 36651 37351 36693 37360
rect 36931 37400 36989 37401
rect 36931 37360 36940 37400
rect 36980 37360 36989 37400
rect 36931 37359 36989 37360
rect 37323 37400 37365 37409
rect 37323 37360 37324 37400
rect 37364 37360 37365 37400
rect 37323 37351 37365 37360
rect 37699 37400 37757 37401
rect 37699 37360 37708 37400
rect 37748 37360 37757 37400
rect 37699 37359 37757 37360
rect 38563 37400 38621 37401
rect 38563 37360 38572 37400
rect 38612 37360 38621 37400
rect 38563 37359 38621 37360
rect 41059 37400 41117 37401
rect 41059 37360 41068 37400
rect 41108 37360 41117 37400
rect 41059 37359 41117 37360
rect 41923 37400 41981 37401
rect 41923 37360 41932 37400
rect 41972 37360 41981 37400
rect 41923 37359 41981 37360
rect 23595 37316 23637 37325
rect 23595 37276 23596 37316
rect 23636 37276 23637 37316
rect 23595 37267 23637 37276
rect 30219 37316 30261 37325
rect 30219 37276 30220 37316
rect 30260 37276 30261 37316
rect 30219 37267 30261 37276
rect 36555 37316 36597 37325
rect 36555 37276 36556 37316
rect 36596 37276 36597 37316
rect 36555 37267 36597 37276
rect 42315 37316 42357 37325
rect 42315 37276 42316 37316
rect 42356 37276 42357 37316
rect 42315 37267 42357 37276
rect 19563 37232 19605 37241
rect 19563 37192 19564 37232
rect 19604 37192 19605 37232
rect 19563 37183 19605 37192
rect 20419 37232 20477 37233
rect 20419 37192 20428 37232
rect 20468 37192 20477 37232
rect 20419 37191 20477 37192
rect 23395 37232 23453 37233
rect 23395 37192 23404 37232
rect 23444 37192 23453 37232
rect 23395 37191 23453 37192
rect 25987 37232 26045 37233
rect 25987 37192 25996 37232
rect 26036 37192 26045 37232
rect 25987 37191 26045 37192
rect 29251 37232 29309 37233
rect 29251 37192 29260 37232
rect 29300 37192 29309 37232
rect 29251 37191 29309 37192
rect 30027 37232 30069 37241
rect 30027 37192 30028 37232
rect 30068 37192 30069 37232
rect 30027 37183 30069 37192
rect 32611 37232 32669 37233
rect 32611 37192 32620 37232
rect 32660 37192 32669 37232
rect 32611 37191 32669 37192
rect 33099 37232 33141 37241
rect 33099 37192 33100 37232
rect 33140 37192 33141 37232
rect 33099 37183 33141 37192
rect 33283 37232 33341 37233
rect 33283 37192 33292 37232
rect 33332 37192 33341 37232
rect 39715 37232 39773 37233
rect 33283 37191 33341 37192
rect 36267 37190 36309 37199
rect 39715 37192 39724 37232
rect 39764 37192 39773 37232
rect 39715 37191 39773 37192
rect 39907 37232 39965 37233
rect 39907 37192 39916 37232
rect 39956 37192 39965 37232
rect 39907 37191 39965 37192
rect 36267 37150 36268 37190
rect 36308 37150 36309 37190
rect 36267 37141 36309 37150
rect 576 37064 83328 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 83328 37064
rect 576 37000 83328 37024
rect 22539 36954 22581 36963
rect 22539 36914 22540 36954
rect 22580 36914 22581 36954
rect 22539 36905 22581 36914
rect 21091 36896 21149 36897
rect 21091 36856 21100 36896
rect 21140 36856 21149 36896
rect 21091 36855 21149 36856
rect 23403 36896 23445 36905
rect 23403 36856 23404 36896
rect 23444 36856 23445 36896
rect 23403 36847 23445 36856
rect 24835 36896 24893 36897
rect 24835 36856 24844 36896
rect 24884 36856 24893 36896
rect 24835 36855 24893 36856
rect 25123 36896 25181 36897
rect 25123 36856 25132 36896
rect 25172 36856 25181 36896
rect 25123 36855 25181 36856
rect 25603 36896 25661 36897
rect 25603 36856 25612 36896
rect 25652 36856 25661 36896
rect 25603 36855 25661 36856
rect 28099 36896 28157 36897
rect 28099 36856 28108 36896
rect 28148 36856 28157 36896
rect 28099 36855 28157 36856
rect 32035 36896 32093 36897
rect 32035 36856 32044 36896
rect 32084 36856 32093 36896
rect 32035 36855 32093 36856
rect 38467 36896 38525 36897
rect 38467 36856 38476 36896
rect 38516 36856 38525 36896
rect 38467 36855 38525 36856
rect 25315 36812 25373 36813
rect 25315 36772 25324 36812
rect 25364 36772 25373 36812
rect 25315 36771 25373 36772
rect 26275 36812 26333 36813
rect 26275 36772 26284 36812
rect 26324 36772 26333 36812
rect 26275 36771 26333 36772
rect 29643 36812 29685 36821
rect 29643 36772 29644 36812
rect 29684 36772 29685 36812
rect 29643 36763 29685 36772
rect 32715 36812 32757 36821
rect 32715 36772 32716 36812
rect 32756 36772 32757 36812
rect 32715 36763 32757 36772
rect 36075 36812 36117 36821
rect 36075 36772 36076 36812
rect 36116 36772 36117 36812
rect 36075 36763 36117 36772
rect 40011 36812 40053 36821
rect 40011 36772 40012 36812
rect 40052 36772 40053 36812
rect 40011 36763 40053 36772
rect 33091 36741 33149 36742
rect 18699 36728 18741 36737
rect 18699 36688 18700 36728
rect 18740 36688 18741 36728
rect 18699 36679 18741 36688
rect 19075 36728 19133 36729
rect 19075 36688 19084 36728
rect 19124 36688 19133 36728
rect 19075 36687 19133 36688
rect 19939 36728 19997 36729
rect 19939 36688 19948 36728
rect 19988 36688 19997 36728
rect 19939 36687 19997 36688
rect 21379 36728 21437 36729
rect 21379 36688 21388 36728
rect 21428 36688 21437 36728
rect 21379 36687 21437 36688
rect 22347 36728 22389 36737
rect 22347 36688 22348 36728
rect 22388 36688 22389 36728
rect 22347 36679 22389 36688
rect 22435 36728 22493 36729
rect 22435 36688 22444 36728
rect 22484 36688 22493 36728
rect 22435 36687 22493 36688
rect 23019 36728 23061 36737
rect 23019 36688 23020 36728
rect 23060 36688 23061 36728
rect 23019 36679 23061 36688
rect 23107 36728 23165 36729
rect 23107 36688 23116 36728
rect 23156 36688 23165 36728
rect 23107 36687 23165 36688
rect 23875 36728 23933 36729
rect 23875 36688 23884 36728
rect 23924 36688 23933 36728
rect 23875 36687 23933 36688
rect 23979 36728 24021 36737
rect 23979 36688 23980 36728
rect 24020 36688 24021 36728
rect 23979 36679 24021 36688
rect 24163 36728 24221 36729
rect 24163 36688 24172 36728
rect 24212 36688 24221 36728
rect 24163 36687 24221 36688
rect 24355 36728 24413 36729
rect 24355 36688 24364 36728
rect 24404 36688 24413 36728
rect 24355 36687 24413 36688
rect 24459 36728 24501 36737
rect 24459 36688 24460 36728
rect 24500 36688 24501 36728
rect 24459 36679 24501 36688
rect 24651 36728 24693 36737
rect 24651 36688 24652 36728
rect 24692 36688 24693 36728
rect 24651 36679 24693 36688
rect 24931 36728 24989 36729
rect 24931 36688 24940 36728
rect 24980 36688 24989 36728
rect 24931 36687 24989 36688
rect 25515 36728 25557 36737
rect 25515 36688 25516 36728
rect 25556 36688 25557 36728
rect 25515 36679 25557 36688
rect 25611 36728 25653 36737
rect 25611 36688 25612 36728
rect 25652 36688 25653 36728
rect 25611 36679 25653 36688
rect 26371 36728 26429 36729
rect 26371 36688 26380 36728
rect 26420 36688 26429 36728
rect 26371 36687 26429 36688
rect 26755 36728 26813 36729
rect 26755 36688 26764 36728
rect 26804 36688 26813 36728
rect 26755 36687 26813 36688
rect 27147 36728 27189 36737
rect 27147 36688 27148 36728
rect 27188 36688 27189 36728
rect 27147 36679 27189 36688
rect 27243 36728 27285 36737
rect 27243 36688 27244 36728
rect 27284 36688 27285 36728
rect 27243 36679 27285 36688
rect 27339 36728 27381 36737
rect 27339 36688 27340 36728
rect 27380 36688 27381 36728
rect 27339 36679 27381 36688
rect 27435 36728 27477 36737
rect 27435 36688 27436 36728
rect 27476 36688 27477 36728
rect 27435 36679 27477 36688
rect 28003 36728 28061 36729
rect 28003 36688 28012 36728
rect 28052 36688 28061 36728
rect 28003 36687 28061 36688
rect 30019 36728 30077 36729
rect 30019 36688 30028 36728
rect 30068 36688 30077 36728
rect 30019 36687 30077 36688
rect 30883 36728 30941 36729
rect 30883 36688 30892 36728
rect 30932 36688 30941 36728
rect 33091 36701 33100 36741
rect 33140 36701 33149 36741
rect 33091 36700 33149 36701
rect 33955 36728 34013 36729
rect 30883 36687 30941 36688
rect 33955 36688 33964 36728
rect 34004 36688 34013 36728
rect 33955 36687 34013 36688
rect 35307 36728 35349 36737
rect 35307 36688 35308 36728
rect 35348 36688 35349 36728
rect 35307 36679 35349 36688
rect 35499 36728 35541 36737
rect 35499 36688 35500 36728
rect 35540 36688 35541 36728
rect 35499 36679 35541 36688
rect 35691 36728 35733 36737
rect 35691 36688 35692 36728
rect 35732 36688 35733 36728
rect 35691 36679 35733 36688
rect 35883 36728 35925 36737
rect 35883 36688 35884 36728
rect 35924 36688 35925 36728
rect 35883 36679 35925 36688
rect 36451 36728 36509 36729
rect 36451 36688 36460 36728
rect 36500 36688 36509 36728
rect 36451 36687 36509 36688
rect 37315 36728 37373 36729
rect 37315 36688 37324 36728
rect 37364 36688 37373 36728
rect 37315 36687 37373 36688
rect 39619 36728 39677 36729
rect 39619 36688 39628 36728
rect 39668 36688 39677 36728
rect 39619 36687 39677 36688
rect 39915 36728 39957 36737
rect 39915 36688 39916 36728
rect 39956 36688 39957 36728
rect 39915 36679 39957 36688
rect 41547 36728 41589 36737
rect 41547 36688 41548 36728
rect 41588 36688 41589 36728
rect 41547 36679 41589 36688
rect 41923 36728 41981 36729
rect 41923 36688 41932 36728
rect 41972 36688 41981 36728
rect 41923 36687 41981 36688
rect 42787 36728 42845 36729
rect 42787 36688 42796 36728
rect 42836 36688 42845 36728
rect 42787 36687 42845 36688
rect 32515 36644 32573 36645
rect 32515 36604 32524 36644
rect 32564 36604 32573 36644
rect 32515 36603 32573 36604
rect 35787 36644 35829 36653
rect 35787 36604 35788 36644
rect 35828 36604 35829 36644
rect 35787 36595 35829 36604
rect 22059 36560 22101 36569
rect 22059 36520 22060 36560
rect 22100 36520 22101 36560
rect 22059 36511 22101 36520
rect 24171 36560 24213 36569
rect 24171 36520 24172 36560
rect 24212 36520 24213 36560
rect 24171 36511 24213 36520
rect 27619 36560 27677 36561
rect 27619 36520 27628 36560
rect 27668 36520 27677 36560
rect 27619 36519 27677 36520
rect 27811 36560 27869 36561
rect 27811 36520 27820 36560
rect 27860 36520 27869 36560
rect 27811 36519 27869 36520
rect 40291 36560 40349 36561
rect 40291 36520 40300 36560
rect 40340 36520 40349 36560
rect 40291 36519 40349 36520
rect 21291 36476 21333 36485
rect 21291 36436 21292 36476
rect 21332 36436 21333 36476
rect 21291 36427 21333 36436
rect 24651 36476 24693 36485
rect 24651 36436 24652 36476
rect 24692 36436 24693 36476
rect 24651 36427 24693 36436
rect 32331 36476 32373 36485
rect 32331 36436 32332 36476
rect 32372 36436 32373 36476
rect 32331 36427 32373 36436
rect 35107 36476 35165 36477
rect 35107 36436 35116 36476
rect 35156 36436 35165 36476
rect 35107 36435 35165 36436
rect 35307 36476 35349 36485
rect 35307 36436 35308 36476
rect 35348 36436 35349 36476
rect 35307 36427 35349 36436
rect 43939 36476 43997 36477
rect 43939 36436 43948 36476
rect 43988 36436 43997 36476
rect 43939 36435 43997 36436
rect 576 36308 83328 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 83328 36308
rect 576 36244 83328 36268
rect 20523 36140 20565 36149
rect 20523 36100 20524 36140
rect 20564 36100 20565 36140
rect 20523 36091 20565 36100
rect 21963 36140 22005 36149
rect 21963 36100 21964 36140
rect 22004 36100 22005 36140
rect 21963 36091 22005 36100
rect 25699 36140 25757 36141
rect 25699 36100 25708 36140
rect 25748 36100 25757 36140
rect 25699 36099 25757 36100
rect 32227 36140 32285 36141
rect 32227 36100 32236 36140
rect 32276 36100 32285 36140
rect 32227 36099 32285 36100
rect 41635 36140 41693 36141
rect 41635 36100 41644 36140
rect 41684 36100 41693 36140
rect 41635 36099 41693 36100
rect 16867 36056 16925 36057
rect 16867 36016 16876 36056
rect 16916 36016 16925 36056
rect 16867 36015 16925 36016
rect 19171 36056 19229 36057
rect 19171 36016 19180 36056
rect 19220 36016 19229 36056
rect 19171 36015 19229 36016
rect 20323 36056 20381 36057
rect 20323 36016 20332 36056
rect 20372 36016 20381 36056
rect 20323 36015 20381 36016
rect 22915 36056 22973 36057
rect 22915 36016 22924 36056
rect 22964 36016 22973 36056
rect 22915 36015 22973 36016
rect 27811 36056 27869 36057
rect 27811 36016 27820 36056
rect 27860 36016 27869 36056
rect 27811 36015 27869 36016
rect 35115 36056 35157 36065
rect 35115 36016 35116 36056
rect 35156 36016 35157 36056
rect 35115 36007 35157 36016
rect 36451 36056 36509 36057
rect 36451 36016 36460 36056
rect 36500 36016 36509 36056
rect 36451 36015 36509 36016
rect 40579 36056 40637 36057
rect 40579 36016 40588 36056
rect 40628 36016 40637 36056
rect 40579 36015 40637 36016
rect 43747 36056 43805 36057
rect 43747 36016 43756 36056
rect 43796 36016 43805 36056
rect 43747 36015 43805 36016
rect 46243 36056 46301 36057
rect 46243 36016 46252 36056
rect 46292 36016 46301 36056
rect 46243 36015 46301 36016
rect 49603 36056 49661 36057
rect 49603 36016 49612 36056
rect 49652 36016 49661 36056
rect 49603 36015 49661 36016
rect 51331 36056 51389 36057
rect 51331 36016 51340 36056
rect 51380 36016 51389 36056
rect 51331 36015 51389 36016
rect 52291 36056 52349 36057
rect 52291 36016 52300 36056
rect 52340 36016 52349 36056
rect 52291 36015 52349 36016
rect 13891 35972 13949 35973
rect 13891 35932 13900 35972
rect 13940 35932 13949 35972
rect 13891 35931 13949 35932
rect 35307 35972 35349 35981
rect 35307 35932 35308 35972
rect 35348 35932 35349 35972
rect 35307 35923 35349 35932
rect 43939 35972 43997 35973
rect 43939 35932 43948 35972
rect 43988 35932 43997 35972
rect 43939 35931 43997 35932
rect 44515 35972 44573 35973
rect 44515 35932 44524 35972
rect 44564 35932 44573 35972
rect 44515 35931 44573 35932
rect 35115 35899 35157 35908
rect 16195 35888 16253 35889
rect 16195 35848 16204 35888
rect 16244 35848 16253 35888
rect 16195 35847 16253 35848
rect 16491 35888 16533 35897
rect 16491 35848 16492 35888
rect 16532 35848 16533 35888
rect 16491 35839 16533 35848
rect 18499 35888 18557 35889
rect 18499 35848 18508 35888
rect 18548 35848 18557 35888
rect 18499 35847 18557 35848
rect 18795 35888 18837 35897
rect 18795 35848 18796 35888
rect 18836 35848 18837 35888
rect 18795 35839 18837 35848
rect 19651 35888 19709 35889
rect 19651 35848 19660 35888
rect 19700 35848 19709 35888
rect 19651 35847 19709 35848
rect 19947 35888 19989 35897
rect 19947 35848 19948 35888
rect 19988 35848 19989 35888
rect 19947 35839 19989 35848
rect 20811 35888 20853 35897
rect 20811 35848 20812 35888
rect 20852 35848 20853 35888
rect 20811 35839 20853 35848
rect 20899 35888 20957 35889
rect 20899 35848 20908 35888
rect 20948 35848 20957 35888
rect 20899 35847 20957 35848
rect 21195 35888 21237 35897
rect 21195 35848 21196 35888
rect 21236 35848 21237 35888
rect 21195 35839 21237 35848
rect 21483 35888 21525 35897
rect 21483 35848 21484 35888
rect 21524 35848 21525 35888
rect 21483 35839 21525 35848
rect 21667 35888 21725 35889
rect 21667 35848 21676 35888
rect 21716 35848 21725 35888
rect 21667 35847 21725 35848
rect 21771 35888 21813 35897
rect 21771 35848 21772 35888
rect 21812 35848 21813 35888
rect 21771 35839 21813 35848
rect 21955 35888 22013 35889
rect 21955 35848 21964 35888
rect 22004 35848 22013 35888
rect 21955 35847 22013 35848
rect 22243 35888 22301 35889
rect 22243 35848 22252 35888
rect 22292 35848 22301 35888
rect 22243 35847 22301 35848
rect 22539 35888 22581 35897
rect 22539 35848 22540 35888
rect 22580 35848 22581 35888
rect 22539 35839 22581 35848
rect 23307 35888 23349 35897
rect 23307 35848 23308 35888
rect 23348 35848 23349 35888
rect 23307 35839 23349 35848
rect 23683 35888 23741 35889
rect 23683 35848 23692 35888
rect 23732 35848 23741 35888
rect 23683 35847 23741 35848
rect 24547 35888 24605 35889
rect 24547 35848 24556 35888
rect 24596 35848 24605 35888
rect 24547 35847 24605 35848
rect 27091 35888 27149 35889
rect 27091 35848 27100 35888
rect 27140 35848 27149 35888
rect 27091 35847 27149 35848
rect 27531 35888 27573 35897
rect 27531 35848 27532 35888
rect 27572 35848 27573 35888
rect 27531 35839 27573 35848
rect 27723 35888 27765 35897
rect 27723 35848 27724 35888
rect 27764 35848 27765 35888
rect 27723 35839 27765 35848
rect 27819 35888 27861 35897
rect 27819 35848 27820 35888
rect 27860 35848 27861 35888
rect 27819 35839 27861 35848
rect 31555 35888 31613 35889
rect 31555 35848 31564 35888
rect 31604 35848 31613 35888
rect 31555 35847 31613 35848
rect 31851 35888 31893 35897
rect 31851 35848 31852 35888
rect 31892 35848 31893 35888
rect 31851 35839 31893 35848
rect 31947 35888 31989 35897
rect 31947 35848 31948 35888
rect 31988 35848 31989 35888
rect 31947 35839 31989 35848
rect 32515 35888 32573 35889
rect 32515 35848 32524 35888
rect 32564 35848 32573 35888
rect 32515 35847 32573 35848
rect 34819 35888 34877 35889
rect 34819 35848 34828 35888
rect 34868 35848 34877 35888
rect 34819 35847 34877 35848
rect 34923 35888 34965 35897
rect 34923 35848 34924 35888
rect 34964 35848 34965 35888
rect 35115 35859 35116 35899
rect 35156 35859 35157 35899
rect 35115 35850 35157 35859
rect 35395 35888 35453 35889
rect 34923 35839 34965 35848
rect 35395 35848 35404 35888
rect 35444 35848 35453 35888
rect 35395 35847 35453 35848
rect 35595 35888 35637 35897
rect 35595 35848 35596 35888
rect 35636 35848 35637 35888
rect 35595 35839 35637 35848
rect 35787 35888 35829 35897
rect 35787 35848 35788 35888
rect 35828 35848 35829 35888
rect 35787 35839 35829 35848
rect 35979 35888 36021 35897
rect 35979 35848 35980 35888
rect 36020 35848 36021 35888
rect 35979 35839 36021 35848
rect 36171 35888 36213 35897
rect 36171 35848 36172 35888
rect 36212 35848 36213 35888
rect 36171 35839 36213 35848
rect 36259 35888 36317 35889
rect 36259 35848 36268 35888
rect 36308 35848 36317 35888
rect 36259 35847 36317 35848
rect 36747 35888 36789 35897
rect 36747 35848 36748 35888
rect 36788 35848 36789 35888
rect 36747 35839 36789 35848
rect 36843 35888 36885 35897
rect 36843 35848 36844 35888
rect 36884 35848 36885 35888
rect 36843 35839 36885 35848
rect 37123 35888 37181 35889
rect 37123 35848 37132 35888
rect 37172 35848 37181 35888
rect 37123 35847 37181 35848
rect 39907 35888 39965 35889
rect 39907 35848 39916 35888
rect 39956 35848 39965 35888
rect 39907 35847 39965 35848
rect 40203 35888 40245 35897
rect 40203 35848 40204 35888
rect 40244 35848 40245 35888
rect 40203 35839 40245 35848
rect 40299 35888 40341 35897
rect 40299 35848 40300 35888
rect 40340 35848 40341 35888
rect 40299 35839 40341 35848
rect 40963 35888 41021 35889
rect 40963 35848 40972 35888
rect 41012 35848 41021 35888
rect 40963 35847 41021 35848
rect 41259 35888 41301 35897
rect 41259 35848 41260 35888
rect 41300 35848 41301 35888
rect 41259 35839 41301 35848
rect 41355 35888 41397 35897
rect 41355 35848 41356 35888
rect 41396 35848 41397 35888
rect 41355 35839 41397 35848
rect 43075 35888 43133 35889
rect 43075 35848 43084 35888
rect 43124 35848 43133 35888
rect 43075 35847 43133 35848
rect 43371 35888 43413 35897
rect 43371 35848 43372 35888
rect 43412 35848 43413 35888
rect 43371 35839 43413 35848
rect 45571 35888 45629 35889
rect 45571 35848 45580 35888
rect 45620 35848 45629 35888
rect 45571 35847 45629 35848
rect 45867 35888 45909 35897
rect 45867 35848 45868 35888
rect 45908 35848 45909 35888
rect 45867 35839 45909 35848
rect 48931 35888 48989 35889
rect 48931 35848 48940 35888
rect 48980 35848 48989 35888
rect 48931 35847 48989 35848
rect 49227 35888 49269 35897
rect 49227 35848 49228 35888
rect 49268 35848 49269 35888
rect 49227 35839 49269 35848
rect 50659 35888 50717 35889
rect 50659 35848 50668 35888
rect 50708 35848 50717 35888
rect 50659 35847 50717 35848
rect 50955 35888 50997 35897
rect 50955 35848 50956 35888
rect 50996 35848 50997 35888
rect 50955 35839 50997 35848
rect 51619 35888 51677 35889
rect 51619 35848 51628 35888
rect 51668 35848 51677 35888
rect 51619 35847 51677 35848
rect 51915 35888 51957 35897
rect 51915 35848 51916 35888
rect 51956 35848 51957 35888
rect 51915 35839 51957 35848
rect 16587 35804 16629 35813
rect 16587 35764 16588 35804
rect 16628 35764 16629 35804
rect 16587 35755 16629 35764
rect 18891 35804 18933 35813
rect 18891 35764 18892 35804
rect 18932 35764 18933 35804
rect 18891 35755 18933 35764
rect 20043 35804 20085 35813
rect 20043 35764 20044 35804
rect 20084 35764 20085 35804
rect 20043 35755 20085 35764
rect 22635 35804 22677 35813
rect 22635 35764 22636 35804
rect 22676 35764 22677 35804
rect 22635 35755 22677 35764
rect 26179 35804 26237 35805
rect 26179 35764 26188 35804
rect 26228 35764 26237 35804
rect 26179 35763 26237 35764
rect 43467 35804 43509 35813
rect 43467 35764 43468 35804
rect 43508 35764 43509 35804
rect 43467 35755 43509 35764
rect 45963 35804 46005 35813
rect 45963 35764 45964 35804
rect 46004 35764 46005 35804
rect 45963 35755 46005 35764
rect 49323 35804 49365 35813
rect 49323 35764 49324 35804
rect 49364 35764 49365 35804
rect 49323 35755 49365 35764
rect 51051 35804 51093 35813
rect 51051 35764 51052 35804
rect 51092 35764 51093 35804
rect 51051 35755 51093 35764
rect 52011 35804 52053 35813
rect 52011 35764 52012 35804
rect 52052 35764 52053 35804
rect 52011 35755 52053 35764
rect 14091 35720 14133 35729
rect 14091 35680 14092 35720
rect 14132 35680 14133 35720
rect 14091 35671 14133 35680
rect 21003 35716 21045 35725
rect 21003 35676 21004 35716
rect 21044 35676 21045 35716
rect 21003 35667 21045 35676
rect 21387 35720 21429 35729
rect 21387 35680 21388 35720
rect 21428 35680 21429 35720
rect 21387 35671 21429 35680
rect 34347 35720 34389 35729
rect 34347 35680 34348 35720
rect 34388 35680 34389 35720
rect 34347 35671 34389 35680
rect 35691 35720 35733 35729
rect 35691 35680 35692 35720
rect 35732 35680 35733 35720
rect 35691 35671 35733 35680
rect 36067 35720 36125 35721
rect 36067 35680 36076 35720
rect 36116 35680 36125 35720
rect 36067 35679 36125 35680
rect 44139 35720 44181 35729
rect 44139 35680 44140 35720
rect 44180 35680 44181 35720
rect 44139 35671 44181 35680
rect 44715 35720 44757 35729
rect 44715 35680 44716 35720
rect 44756 35680 44757 35720
rect 44715 35671 44757 35680
rect 576 35552 83328 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 83328 35552
rect 576 35488 83328 35512
rect 17539 35384 17597 35385
rect 17539 35344 17548 35384
rect 17588 35344 17597 35384
rect 17539 35343 17597 35344
rect 28483 35384 28541 35385
rect 28483 35344 28492 35384
rect 28532 35344 28541 35384
rect 28483 35343 28541 35344
rect 33379 35384 33437 35385
rect 33379 35344 33388 35384
rect 33428 35344 33437 35384
rect 33379 35343 33437 35344
rect 38371 35384 38429 35385
rect 38371 35344 38380 35384
rect 38420 35344 38429 35384
rect 38371 35343 38429 35344
rect 43267 35384 43325 35385
rect 43267 35344 43276 35384
rect 43316 35344 43325 35384
rect 43267 35343 43325 35344
rect 44323 35384 44381 35385
rect 44323 35344 44332 35384
rect 44372 35344 44381 35384
rect 44323 35343 44381 35344
rect 51907 35384 51965 35385
rect 51907 35344 51916 35384
rect 51956 35344 51965 35384
rect 51907 35343 51965 35344
rect 19947 35300 19989 35309
rect 19947 35260 19948 35300
rect 19988 35260 19989 35300
rect 19947 35251 19989 35260
rect 20715 35300 20757 35309
rect 20715 35260 20716 35300
rect 20756 35260 20757 35300
rect 20715 35251 20757 35260
rect 26091 35300 26133 35309
rect 26091 35260 26092 35300
rect 26132 35260 26133 35300
rect 26091 35251 26133 35260
rect 35787 35300 35829 35309
rect 35787 35260 35788 35300
rect 35828 35260 35829 35300
rect 35787 35251 35829 35260
rect 35979 35300 36021 35309
rect 35979 35260 35980 35300
rect 36020 35260 36021 35300
rect 35979 35251 36021 35260
rect 46731 35300 46773 35309
rect 46731 35260 46732 35300
rect 46772 35260 46773 35300
rect 46731 35251 46773 35260
rect 49515 35300 49557 35309
rect 49515 35260 49516 35300
rect 49556 35260 49557 35300
rect 49515 35251 49557 35260
rect 52107 35300 52149 35309
rect 52107 35260 52108 35300
rect 52148 35260 52149 35300
rect 52107 35251 52149 35260
rect 13227 35216 13269 35225
rect 13227 35176 13228 35216
rect 13268 35176 13269 35216
rect 13227 35167 13269 35176
rect 13323 35216 13365 35225
rect 13323 35176 13324 35216
rect 13364 35176 13365 35216
rect 13323 35167 13365 35176
rect 13603 35216 13661 35217
rect 13603 35176 13612 35216
rect 13652 35176 13661 35216
rect 13603 35175 13661 35176
rect 14083 35216 14141 35217
rect 14083 35176 14092 35216
rect 14132 35176 14141 35216
rect 14083 35175 14141 35176
rect 14379 35216 14421 35225
rect 14379 35176 14380 35216
rect 14420 35176 14421 35216
rect 14379 35167 14421 35176
rect 14475 35216 14517 35225
rect 14475 35176 14476 35216
rect 14516 35176 14517 35216
rect 14475 35167 14517 35176
rect 14955 35216 14997 35225
rect 14955 35176 14956 35216
rect 14996 35176 14997 35216
rect 14955 35167 14997 35176
rect 15331 35216 15389 35217
rect 15331 35176 15340 35216
rect 15380 35176 15389 35216
rect 15331 35175 15389 35176
rect 16195 35216 16253 35217
rect 16195 35176 16204 35216
rect 16244 35176 16253 35216
rect 16195 35175 16253 35176
rect 18691 35216 18749 35217
rect 18691 35176 18700 35216
rect 18740 35176 18749 35216
rect 18691 35175 18749 35176
rect 19555 35216 19613 35217
rect 19555 35176 19564 35216
rect 19604 35176 19613 35216
rect 19555 35175 19613 35176
rect 21091 35216 21149 35217
rect 21091 35176 21100 35216
rect 21140 35176 21149 35216
rect 21091 35175 21149 35176
rect 21955 35216 22013 35217
rect 21955 35176 21964 35216
rect 22004 35176 22013 35216
rect 21955 35175 22013 35176
rect 25035 35216 25077 35225
rect 25035 35176 25036 35216
rect 25076 35176 25077 35216
rect 25035 35167 25077 35176
rect 26467 35216 26525 35217
rect 26467 35176 26476 35216
rect 26516 35176 26525 35216
rect 26467 35175 26525 35176
rect 27331 35216 27389 35217
rect 27331 35176 27340 35216
rect 27380 35176 27389 35216
rect 27331 35175 27389 35176
rect 30027 35216 30069 35225
rect 30027 35176 30028 35216
rect 30068 35176 30069 35216
rect 30027 35167 30069 35176
rect 30403 35216 30461 35217
rect 30403 35176 30412 35216
rect 30452 35176 30461 35216
rect 30403 35175 30461 35176
rect 31267 35216 31325 35217
rect 31267 35176 31276 35216
rect 31316 35176 31325 35216
rect 31267 35175 31325 35176
rect 34531 35216 34589 35217
rect 34531 35176 34540 35216
rect 34580 35176 34589 35216
rect 34531 35175 34589 35176
rect 35395 35216 35453 35217
rect 35395 35176 35404 35216
rect 35444 35176 35453 35216
rect 35395 35175 35453 35176
rect 36355 35216 36413 35217
rect 36355 35176 36364 35216
rect 36404 35176 36413 35216
rect 36355 35175 36413 35176
rect 37219 35216 37277 35217
rect 37219 35176 37228 35216
rect 37268 35176 37277 35216
rect 37219 35175 37277 35176
rect 40003 35216 40061 35217
rect 40003 35176 40012 35216
rect 40052 35176 40061 35216
rect 40003 35175 40061 35176
rect 40299 35216 40341 35225
rect 40299 35176 40300 35216
rect 40340 35176 40341 35216
rect 40299 35167 40341 35176
rect 40395 35216 40437 35225
rect 40395 35176 40396 35216
rect 40436 35176 40437 35216
rect 40395 35167 40437 35176
rect 40875 35216 40917 35225
rect 40875 35176 40876 35216
rect 40916 35176 40917 35216
rect 40875 35167 40917 35176
rect 41251 35216 41309 35217
rect 41251 35176 41260 35216
rect 41300 35176 41309 35216
rect 41251 35175 41309 35176
rect 42115 35216 42173 35217
rect 42115 35176 42124 35216
rect 42164 35176 42173 35216
rect 42115 35175 42173 35176
rect 45475 35216 45533 35217
rect 45475 35176 45484 35216
rect 45524 35176 45533 35216
rect 45475 35175 45533 35176
rect 46339 35216 46397 35217
rect 46339 35176 46348 35216
rect 46388 35176 46397 35216
rect 46339 35175 46397 35176
rect 46923 35216 46965 35225
rect 46923 35176 46924 35216
rect 46964 35176 46965 35216
rect 46923 35167 46965 35176
rect 47299 35216 47357 35217
rect 47299 35176 47308 35216
rect 47348 35176 47357 35216
rect 47299 35175 47357 35176
rect 48163 35216 48221 35217
rect 48163 35176 48172 35216
rect 48212 35176 48221 35216
rect 48163 35175 48221 35176
rect 49891 35216 49949 35217
rect 49891 35176 49900 35216
rect 49940 35176 49949 35216
rect 49891 35175 49949 35176
rect 50755 35216 50813 35217
rect 50755 35176 50764 35216
rect 50804 35176 50813 35216
rect 50755 35175 50813 35176
rect 52483 35216 52541 35217
rect 52483 35176 52492 35216
rect 52532 35176 52541 35216
rect 52483 35175 52541 35176
rect 53347 35216 53405 35217
rect 53347 35176 53356 35216
rect 53396 35176 53405 35216
rect 53347 35175 53405 35176
rect 64587 35216 64629 35225
rect 64587 35176 64588 35216
rect 64628 35176 64629 35216
rect 64587 35167 64629 35176
rect 70147 35216 70205 35217
rect 70147 35176 70156 35216
rect 70196 35176 70205 35216
rect 70147 35175 70205 35176
rect 10627 35132 10685 35133
rect 10627 35092 10636 35132
rect 10676 35092 10685 35132
rect 10627 35091 10685 35092
rect 20323 35132 20381 35133
rect 20323 35092 20332 35132
rect 20372 35092 20381 35132
rect 20323 35091 20381 35092
rect 43651 35132 43709 35133
rect 43651 35092 43660 35132
rect 43700 35092 43709 35132
rect 43651 35091 43709 35092
rect 43939 35132 43997 35133
rect 43939 35092 43948 35132
rect 43988 35092 43997 35132
rect 43939 35091 43997 35092
rect 14755 35048 14813 35049
rect 14755 35008 14764 35048
rect 14804 35008 14813 35048
rect 14755 35007 14813 35008
rect 20139 35048 20181 35057
rect 20139 35008 20140 35048
rect 20180 35008 20181 35048
rect 20139 34999 20181 35008
rect 40675 35048 40733 35049
rect 40675 35008 40684 35048
rect 40724 35008 40733 35048
rect 40675 35007 40733 35008
rect 64395 35048 64437 35057
rect 64395 35008 64396 35048
rect 64436 35008 64437 35048
rect 64395 34999 64437 35008
rect 10443 34964 10485 34973
rect 10443 34924 10444 34964
rect 10484 34924 10485 34964
rect 10443 34915 10485 34924
rect 12931 34964 12989 34965
rect 12931 34924 12940 34964
rect 12980 34924 12989 34964
rect 12931 34923 12989 34924
rect 17347 34964 17405 34965
rect 17347 34924 17356 34964
rect 17396 34924 17405 34964
rect 17347 34923 17405 34924
rect 17539 34964 17597 34965
rect 17539 34924 17548 34964
rect 17588 34924 17597 34964
rect 17539 34923 17597 34924
rect 23107 34964 23165 34965
rect 23107 34924 23116 34964
rect 23156 34924 23165 34964
rect 23107 34923 23165 34924
rect 25227 34964 25269 34973
rect 25227 34924 25228 34964
rect 25268 34924 25269 34964
rect 25227 34915 25269 34924
rect 32419 34964 32477 34965
rect 32419 34924 32428 34964
rect 32468 34924 32477 34964
rect 32419 34923 32477 34924
rect 43467 34964 43509 34973
rect 43467 34924 43468 34964
rect 43508 34924 43509 34964
rect 43467 34915 43509 34924
rect 44139 34964 44181 34973
rect 44139 34924 44140 34964
rect 44180 34924 44181 34964
rect 44139 34915 44181 34924
rect 49315 34964 49373 34965
rect 49315 34924 49324 34964
rect 49364 34924 49373 34964
rect 49315 34923 49373 34924
rect 51907 34964 51965 34965
rect 51907 34924 51916 34964
rect 51956 34924 51965 34964
rect 51907 34923 51965 34924
rect 54499 34964 54557 34965
rect 54499 34924 54508 34964
rect 54548 34924 54557 34964
rect 54499 34923 54557 34924
rect 576 34796 83328 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 83328 34796
rect 576 34732 83328 34756
rect 19267 34628 19325 34629
rect 19267 34588 19276 34628
rect 19316 34588 19325 34628
rect 19267 34587 19325 34588
rect 30211 34628 30269 34629
rect 30211 34588 30220 34628
rect 30260 34588 30269 34628
rect 30211 34587 30269 34588
rect 46531 34628 46589 34629
rect 46531 34588 46540 34628
rect 46580 34588 46589 34628
rect 46531 34587 46589 34588
rect 47979 34628 48021 34637
rect 47979 34588 47980 34628
rect 48020 34588 48021 34628
rect 47979 34579 48021 34588
rect 7563 34544 7605 34553
rect 7563 34504 7564 34544
rect 7604 34504 7605 34544
rect 7563 34495 7605 34504
rect 10627 34544 10685 34545
rect 10627 34504 10636 34544
rect 10676 34504 10685 34544
rect 10627 34503 10685 34504
rect 26475 34544 26517 34553
rect 26475 34504 26476 34544
rect 26516 34504 26517 34544
rect 26475 34495 26517 34504
rect 27427 34544 27485 34545
rect 27427 34504 27436 34544
rect 27476 34504 27485 34544
rect 27427 34503 27485 34504
rect 31939 34544 31997 34545
rect 31939 34504 31948 34544
rect 31988 34504 31997 34544
rect 31939 34503 31997 34504
rect 36931 34544 36989 34545
rect 36931 34504 36940 34544
rect 36980 34504 36989 34544
rect 36931 34503 36989 34504
rect 70923 34544 70965 34553
rect 70923 34504 70924 34544
rect 70964 34504 70965 34544
rect 70923 34495 70965 34504
rect 25515 34460 25557 34469
rect 25515 34420 25516 34460
rect 25556 34420 25557 34460
rect 25515 34411 25557 34420
rect 26275 34460 26333 34461
rect 26275 34420 26284 34460
rect 26324 34420 26333 34460
rect 26275 34419 26333 34420
rect 7843 34376 7901 34377
rect 7843 34336 7852 34376
rect 7892 34336 7901 34376
rect 7843 34335 7901 34336
rect 9955 34376 10013 34377
rect 9955 34336 9964 34376
rect 10004 34336 10013 34376
rect 9955 34335 10013 34336
rect 10251 34376 10293 34385
rect 10251 34336 10252 34376
rect 10292 34336 10293 34376
rect 10251 34327 10293 34336
rect 10827 34376 10869 34385
rect 10827 34336 10828 34376
rect 10868 34336 10869 34376
rect 10827 34327 10869 34336
rect 11203 34376 11261 34377
rect 11203 34336 11212 34376
rect 11252 34336 11261 34376
rect 11203 34335 11261 34336
rect 12067 34376 12125 34377
rect 12067 34336 12076 34376
rect 12116 34336 12125 34376
rect 12067 34335 12125 34336
rect 13419 34376 13461 34385
rect 13419 34336 13420 34376
rect 13460 34336 13461 34376
rect 13419 34327 13461 34336
rect 13795 34376 13853 34377
rect 13795 34336 13804 34376
rect 13844 34336 13853 34376
rect 13795 34335 13853 34336
rect 14659 34376 14717 34377
rect 14659 34336 14668 34376
rect 14708 34336 14717 34376
rect 14659 34335 14717 34336
rect 16875 34376 16917 34385
rect 16875 34336 16876 34376
rect 16916 34336 16917 34376
rect 16875 34327 16917 34336
rect 17307 34376 17349 34385
rect 17307 34336 17308 34376
rect 17348 34336 17349 34376
rect 17307 34327 17349 34336
rect 18115 34376 18173 34377
rect 18115 34336 18124 34376
rect 18164 34336 18173 34376
rect 18115 34335 18173 34336
rect 19555 34376 19613 34377
rect 19555 34336 19564 34376
rect 19604 34336 19613 34376
rect 19555 34335 19613 34336
rect 20515 34376 20573 34377
rect 20515 34336 20524 34376
rect 20564 34336 20573 34376
rect 20515 34335 20573 34336
rect 20995 34376 21053 34377
rect 20995 34336 21004 34376
rect 21044 34336 21053 34376
rect 20995 34335 21053 34336
rect 21283 34376 21341 34377
rect 21283 34336 21292 34376
rect 21332 34336 21341 34376
rect 21283 34335 21341 34336
rect 22243 34376 22301 34377
rect 22243 34336 22252 34376
rect 22292 34336 22301 34376
rect 22243 34335 22301 34336
rect 23115 34376 23157 34385
rect 23115 34336 23116 34376
rect 23156 34336 23157 34376
rect 23115 34327 23157 34336
rect 23491 34376 23549 34377
rect 23491 34336 23500 34376
rect 23540 34336 23549 34376
rect 23491 34335 23549 34336
rect 24355 34376 24413 34377
rect 24355 34336 24364 34376
rect 24404 34336 24413 34376
rect 24355 34335 24413 34336
rect 26755 34376 26813 34377
rect 26755 34336 26764 34376
rect 26804 34336 26813 34376
rect 26755 34335 26813 34336
rect 27051 34376 27093 34385
rect 27051 34336 27052 34376
rect 27092 34336 27093 34376
rect 27051 34327 27093 34336
rect 27627 34376 27669 34385
rect 27627 34336 27628 34376
rect 27668 34336 27669 34376
rect 27627 34327 27669 34336
rect 28003 34376 28061 34377
rect 28003 34336 28012 34376
rect 28052 34336 28061 34376
rect 28003 34335 28061 34336
rect 28867 34376 28925 34377
rect 28867 34336 28876 34376
rect 28916 34336 28925 34376
rect 28867 34335 28925 34336
rect 30507 34376 30549 34385
rect 30507 34336 30508 34376
rect 30548 34336 30549 34376
rect 30507 34327 30549 34336
rect 30603 34376 30645 34385
rect 30603 34336 30604 34376
rect 30644 34336 30645 34376
rect 30603 34327 30645 34336
rect 30883 34376 30941 34377
rect 30883 34336 30892 34376
rect 30932 34336 30941 34376
rect 30883 34335 30941 34336
rect 31267 34376 31325 34377
rect 31267 34336 31276 34376
rect 31316 34336 31325 34376
rect 31267 34335 31325 34336
rect 31563 34376 31605 34385
rect 31563 34336 31564 34376
rect 31604 34336 31605 34376
rect 31563 34327 31605 34336
rect 32139 34376 32181 34385
rect 32139 34336 32140 34376
rect 32180 34336 32181 34376
rect 32139 34327 32181 34336
rect 32515 34376 32573 34377
rect 32515 34336 32524 34376
rect 32564 34336 32573 34376
rect 32515 34335 32573 34336
rect 33379 34376 33437 34377
rect 33379 34336 33388 34376
rect 33428 34336 33437 34376
rect 33379 34335 33437 34336
rect 35683 34376 35741 34377
rect 35683 34336 35692 34376
rect 35732 34336 35741 34376
rect 35683 34335 35741 34336
rect 36259 34376 36317 34377
rect 36259 34336 36268 34376
rect 36308 34336 36317 34376
rect 36259 34335 36317 34336
rect 36555 34376 36597 34385
rect 36555 34336 36556 34376
rect 36596 34336 36597 34376
rect 36555 34327 36597 34336
rect 38083 34376 38141 34377
rect 38083 34336 38092 34376
rect 38132 34336 38141 34376
rect 38083 34335 38141 34336
rect 39139 34376 39197 34377
rect 39139 34336 39148 34376
rect 39188 34336 39197 34376
rect 39139 34335 39197 34336
rect 40003 34376 40061 34377
rect 40003 34336 40012 34376
rect 40052 34336 40061 34376
rect 40003 34335 40061 34336
rect 42219 34376 42261 34385
rect 42219 34336 42220 34376
rect 42260 34336 42261 34376
rect 42219 34327 42261 34336
rect 43651 34376 43709 34377
rect 43651 34336 43660 34376
rect 43700 34336 43709 34376
rect 43651 34335 43709 34336
rect 43947 34376 43989 34385
rect 43947 34336 43948 34376
rect 43988 34336 43989 34376
rect 43947 34327 43989 34336
rect 44323 34376 44381 34377
rect 44323 34336 44332 34376
rect 44372 34336 44381 34376
rect 44323 34335 44381 34336
rect 45187 34376 45245 34377
rect 45187 34336 45196 34376
rect 45236 34336 45245 34376
rect 45187 34335 45245 34336
rect 46827 34376 46869 34385
rect 46827 34336 46828 34376
rect 46868 34336 46869 34376
rect 46827 34327 46869 34336
rect 46923 34376 46965 34385
rect 46923 34336 46924 34376
rect 46964 34336 46965 34376
rect 46923 34327 46965 34336
rect 47203 34376 47261 34377
rect 47203 34336 47212 34376
rect 47252 34336 47261 34376
rect 47203 34335 47261 34336
rect 49603 34376 49661 34377
rect 49603 34336 49612 34376
rect 49652 34336 49661 34376
rect 49603 34335 49661 34336
rect 50851 34376 50909 34377
rect 50851 34336 50860 34376
rect 50900 34336 50909 34376
rect 50851 34335 50909 34336
rect 52483 34376 52541 34377
rect 52483 34336 52492 34376
rect 52532 34336 52541 34376
rect 52483 34335 52541 34336
rect 53155 34376 53213 34377
rect 53155 34336 53164 34376
rect 53204 34336 53213 34376
rect 53155 34335 53213 34336
rect 54019 34376 54077 34377
rect 54019 34336 54028 34376
rect 54068 34336 54077 34376
rect 54019 34335 54077 34336
rect 61507 34376 61565 34377
rect 61507 34336 61516 34376
rect 61556 34336 61565 34376
rect 61507 34335 61565 34336
rect 62467 34376 62525 34377
rect 62467 34336 62476 34376
rect 62516 34336 62525 34376
rect 62467 34335 62525 34336
rect 62755 34376 62813 34377
rect 62755 34336 62764 34376
rect 62804 34336 62813 34376
rect 62755 34335 62813 34336
rect 64203 34376 64245 34385
rect 64203 34336 64204 34376
rect 64244 34336 64245 34376
rect 64203 34327 64245 34336
rect 65443 34376 65501 34377
rect 65443 34336 65452 34376
rect 65492 34336 65501 34376
rect 65443 34335 65501 34336
rect 66315 34376 66357 34385
rect 66315 34336 66316 34376
rect 66356 34336 66357 34376
rect 66315 34327 66357 34336
rect 68035 34376 68093 34377
rect 68035 34336 68044 34376
rect 68084 34336 68093 34376
rect 68035 34335 68093 34336
rect 68907 34376 68949 34385
rect 68907 34336 68908 34376
rect 68948 34336 68949 34376
rect 68907 34327 68949 34336
rect 69283 34376 69341 34377
rect 69283 34336 69292 34376
rect 69332 34336 69341 34376
rect 69283 34335 69341 34336
rect 70155 34376 70197 34385
rect 70155 34336 70156 34376
rect 70196 34336 70197 34376
rect 70155 34327 70197 34336
rect 70627 34376 70685 34377
rect 70627 34336 70636 34376
rect 70676 34336 70685 34376
rect 70627 34335 70685 34336
rect 10347 34292 10389 34301
rect 10347 34252 10348 34292
rect 10388 34252 10389 34292
rect 10347 34243 10389 34252
rect 27147 34292 27189 34301
rect 27147 34252 27148 34292
rect 27188 34252 27189 34292
rect 27147 34243 27189 34252
rect 31659 34292 31701 34301
rect 31659 34252 31660 34292
rect 31700 34252 31701 34292
rect 31659 34243 31701 34252
rect 36651 34292 36693 34301
rect 36651 34252 36652 34292
rect 36692 34252 36693 34292
rect 36651 34243 36693 34252
rect 38763 34292 38805 34301
rect 38763 34252 38764 34292
rect 38804 34252 38805 34292
rect 38763 34243 38805 34252
rect 52779 34292 52821 34301
rect 52779 34252 52780 34292
rect 52820 34252 52821 34292
rect 52779 34243 52821 34252
rect 7371 34208 7413 34217
rect 7371 34168 7372 34208
rect 7412 34168 7413 34208
rect 7371 34159 7413 34168
rect 13219 34208 13277 34209
rect 13219 34168 13228 34208
rect 13268 34168 13277 34208
rect 13219 34167 13277 34168
rect 15811 34208 15869 34209
rect 15811 34168 15820 34208
rect 15860 34168 15869 34208
rect 15811 34167 15869 34168
rect 19267 34208 19325 34209
rect 19267 34168 19276 34208
rect 19316 34168 19325 34208
rect 19267 34167 19325 34168
rect 30019 34208 30077 34209
rect 30019 34168 30028 34208
rect 30068 34168 30077 34208
rect 30019 34167 30077 34168
rect 34531 34208 34589 34209
rect 34531 34168 34540 34208
rect 34580 34168 34589 34208
rect 34531 34167 34589 34168
rect 35211 34208 35253 34217
rect 35211 34168 35212 34208
rect 35252 34168 35253 34208
rect 35211 34159 35253 34168
rect 37611 34208 37653 34217
rect 37611 34168 37612 34208
rect 37652 34168 37653 34208
rect 37611 34159 37653 34168
rect 41155 34208 41213 34209
rect 41155 34168 41164 34208
rect 41204 34168 41213 34208
rect 41155 34167 41213 34168
rect 46339 34208 46397 34209
rect 46339 34168 46348 34208
rect 46388 34168 46397 34208
rect 46339 34167 46397 34168
rect 50379 34208 50421 34217
rect 50379 34168 50380 34208
rect 50420 34168 50421 34208
rect 50379 34159 50421 34168
rect 52011 34208 52053 34217
rect 52011 34168 52012 34208
rect 52052 34168 52053 34208
rect 52011 34159 52053 34168
rect 55171 34208 55229 34209
rect 55171 34168 55180 34208
rect 55220 34168 55229 34208
rect 55171 34167 55229 34168
rect 64587 34208 64629 34217
rect 64587 34168 64588 34208
rect 64628 34168 64629 34208
rect 64587 34159 64629 34168
rect 68523 34208 68565 34217
rect 68523 34168 68524 34208
rect 68564 34168 68565 34208
rect 68523 34159 68565 34168
rect 576 34040 83328 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 83328 34040
rect 576 33976 83328 34000
rect 80811 33704 80853 33713
rect 80811 33664 80812 33704
rect 80852 33664 80853 33704
rect 80811 33655 80853 33664
rect 81187 33704 81245 33705
rect 81187 33664 81196 33704
rect 81236 33664 81245 33704
rect 81187 33663 81245 33664
rect 82051 33704 82109 33705
rect 82051 33664 82060 33704
rect 82100 33664 82109 33704
rect 82051 33663 82109 33664
rect 83203 33452 83261 33453
rect 83203 33412 83212 33452
rect 83252 33412 83261 33452
rect 83203 33411 83261 33412
rect 576 33284 5952 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 5952 33284
rect 576 33220 5952 33244
rect 74016 33284 83328 33308
rect 74016 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 83328 33284
rect 74016 33220 83328 33244
rect 80515 33116 80573 33117
rect 80515 33076 80524 33116
rect 80564 33076 80573 33116
rect 80515 33075 80573 33076
rect 5539 32948 5597 32949
rect 5539 32908 5548 32948
rect 5588 32908 5597 32948
rect 5539 32907 5597 32908
rect 80131 32948 80189 32949
rect 80131 32908 80140 32948
rect 80180 32908 80189 32948
rect 80131 32907 80189 32908
rect 82051 32948 82109 32949
rect 82051 32908 82060 32948
rect 82100 32908 82109 32948
rect 82051 32907 82109 32908
rect 80811 32864 80853 32873
rect 80811 32824 80812 32864
rect 80852 32824 80853 32864
rect 80811 32815 80853 32824
rect 80907 32864 80949 32873
rect 80907 32824 80908 32864
rect 80948 32824 80949 32864
rect 80907 32815 80949 32824
rect 81187 32864 81245 32865
rect 81187 32824 81196 32864
rect 81236 32824 81245 32864
rect 81187 32823 81245 32824
rect 5355 32696 5397 32705
rect 5355 32656 5356 32696
rect 5396 32656 5397 32696
rect 5355 32647 5397 32656
rect 80331 32696 80373 32705
rect 80331 32656 80332 32696
rect 80372 32656 80373 32696
rect 80331 32647 80373 32656
rect 81867 32696 81909 32705
rect 81867 32656 81868 32696
rect 81908 32656 81909 32696
rect 81867 32647 81909 32656
rect 576 32528 5952 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 5952 32528
rect 576 32464 5952 32488
rect 74016 32528 83328 32552
rect 74016 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 83328 32528
rect 74016 32464 83328 32488
rect 4587 32360 4629 32369
rect 4587 32320 4588 32360
rect 4628 32320 4629 32360
rect 4587 32311 4629 32320
rect 5731 32192 5789 32193
rect 5731 32152 5740 32192
rect 5780 32152 5789 32192
rect 5731 32151 5789 32152
rect 80811 32192 80853 32201
rect 80811 32152 80812 32192
rect 80852 32152 80853 32192
rect 80811 32143 80853 32152
rect 81187 32192 81245 32193
rect 81187 32152 81196 32192
rect 81236 32152 81245 32192
rect 81187 32151 81245 32152
rect 82051 32192 82109 32193
rect 82051 32152 82060 32192
rect 82100 32152 82109 32192
rect 82051 32151 82109 32152
rect 4387 32108 4445 32109
rect 4387 32068 4396 32108
rect 4436 32068 4445 32108
rect 4387 32067 4445 32068
rect 4587 31940 4629 31949
rect 4587 31900 4588 31940
rect 4628 31900 4629 31940
rect 4587 31891 4629 31900
rect 5067 31940 5109 31949
rect 5067 31900 5068 31940
rect 5108 31900 5109 31940
rect 5067 31891 5109 31900
rect 83203 31940 83261 31941
rect 83203 31900 83212 31940
rect 83252 31900 83261 31940
rect 83203 31899 83261 31900
rect 576 31772 5952 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 5952 31772
rect 576 31708 5952 31732
rect 74016 31772 83328 31796
rect 74016 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 83328 31772
rect 74016 31708 83328 31732
rect 5827 31604 5885 31605
rect 5827 31564 5836 31604
rect 5876 31564 5885 31604
rect 5827 31563 5885 31564
rect 80707 31604 80765 31605
rect 80707 31564 80716 31604
rect 80756 31564 80765 31604
rect 80707 31563 80765 31564
rect 80323 31436 80381 31437
rect 80323 31396 80332 31436
rect 80372 31396 80381 31436
rect 80323 31395 80381 31396
rect 3811 31352 3869 31353
rect 3811 31312 3820 31352
rect 3860 31312 3869 31352
rect 3811 31311 3869 31312
rect 4675 31352 4733 31353
rect 4675 31312 4684 31352
rect 4724 31312 4733 31352
rect 4675 31311 4733 31312
rect 81099 31352 81141 31361
rect 81099 31312 81100 31352
rect 81140 31312 81141 31352
rect 81099 31303 81141 31312
rect 81379 31352 81437 31353
rect 81379 31312 81388 31352
rect 81428 31312 81437 31352
rect 81379 31311 81437 31312
rect 3435 31268 3477 31277
rect 3435 31228 3436 31268
rect 3476 31228 3477 31268
rect 3435 31219 3477 31228
rect 81003 31268 81045 31277
rect 81003 31228 81004 31268
rect 81044 31228 81045 31268
rect 81003 31219 81045 31228
rect 5827 31184 5885 31185
rect 5827 31144 5836 31184
rect 5876 31144 5885 31184
rect 5827 31143 5885 31144
rect 80139 31184 80181 31193
rect 80139 31144 80140 31184
rect 80180 31144 80181 31184
rect 80139 31135 80181 31144
rect 576 31016 5952 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 5952 31016
rect 576 30952 5952 30976
rect 74016 31016 83328 31040
rect 74016 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 83328 31016
rect 74016 30952 83328 30976
rect 82915 30848 82973 30849
rect 82915 30808 82924 30848
rect 82964 30808 82973 30848
rect 82915 30807 82973 30808
rect 4491 30764 4533 30773
rect 4491 30724 4492 30764
rect 4532 30724 4533 30764
rect 4491 30715 4533 30724
rect 80043 30764 80085 30773
rect 80043 30724 80044 30764
rect 80084 30724 80085 30764
rect 80043 30715 80085 30724
rect 4587 30680 4629 30689
rect 4587 30640 4588 30680
rect 4628 30640 4629 30680
rect 4587 30631 4629 30640
rect 4867 30680 4925 30681
rect 4867 30640 4876 30680
rect 4916 30640 4925 30680
rect 4867 30639 4925 30640
rect 79651 30680 79709 30681
rect 79651 30640 79660 30680
rect 79700 30640 79709 30680
rect 79651 30639 79709 30640
rect 79947 30680 79989 30689
rect 79947 30640 79948 30680
rect 79988 30640 79989 30680
rect 79947 30631 79989 30640
rect 80523 30680 80565 30689
rect 80523 30640 80524 30680
rect 80564 30640 80565 30680
rect 80523 30631 80565 30640
rect 80899 30680 80957 30681
rect 80899 30640 80908 30680
rect 80948 30640 80957 30680
rect 80899 30639 80957 30640
rect 81763 30680 81821 30681
rect 81763 30640 81772 30680
rect 81812 30640 81821 30680
rect 81763 30639 81821 30640
rect 79171 30596 79229 30597
rect 79171 30556 79180 30596
rect 79220 30556 79229 30596
rect 79171 30555 79229 30556
rect 4195 30512 4253 30513
rect 4195 30472 4204 30512
rect 4244 30472 4253 30512
rect 4195 30471 4253 30472
rect 80323 30512 80381 30513
rect 80323 30472 80332 30512
rect 80372 30472 80381 30512
rect 80323 30471 80381 30472
rect 79371 30428 79413 30437
rect 79371 30388 79372 30428
rect 79412 30388 79413 30428
rect 79371 30379 79413 30388
rect 576 30260 5952 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 5952 30260
rect 576 30196 5952 30220
rect 74016 30260 83328 30284
rect 74016 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 83328 30260
rect 74016 30196 83328 30220
rect 81379 30008 81437 30009
rect 81379 29968 81388 30008
rect 81428 29968 81437 30008
rect 81379 29967 81437 29968
rect 79171 29840 79229 29841
rect 79171 29800 79180 29840
rect 79220 29800 79229 29840
rect 79171 29799 79229 29800
rect 80035 29840 80093 29841
rect 80035 29800 80044 29840
rect 80084 29800 80093 29840
rect 80035 29799 80093 29800
rect 81675 29840 81717 29849
rect 81675 29800 81676 29840
rect 81716 29800 81717 29840
rect 81675 29791 81717 29800
rect 81771 29840 81813 29849
rect 81771 29800 81772 29840
rect 81812 29800 81813 29840
rect 81771 29791 81813 29800
rect 82051 29840 82109 29841
rect 82051 29800 82060 29840
rect 82100 29800 82109 29840
rect 82051 29799 82109 29800
rect 78795 29756 78837 29765
rect 78795 29716 78796 29756
rect 78836 29716 78837 29756
rect 78795 29707 78837 29716
rect 81187 29672 81245 29673
rect 81187 29632 81196 29672
rect 81236 29632 81245 29672
rect 81187 29631 81245 29632
rect 576 29504 5952 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 5952 29504
rect 576 29440 5952 29464
rect 74016 29504 83328 29528
rect 74016 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 83328 29504
rect 74016 29440 83328 29464
rect 83203 29336 83261 29337
rect 83203 29296 83212 29336
rect 83252 29296 83261 29336
rect 83203 29295 83261 29296
rect 79659 29252 79701 29261
rect 79659 29212 79660 29252
rect 79700 29212 79701 29252
rect 79659 29203 79701 29212
rect 80811 29252 80853 29261
rect 80811 29212 80812 29252
rect 80852 29212 80853 29252
rect 80811 29203 80853 29212
rect 4579 29168 4637 29169
rect 4579 29128 4588 29168
rect 4628 29128 4637 29168
rect 4579 29127 4637 29128
rect 5443 29168 5501 29169
rect 5443 29128 5452 29168
rect 5492 29128 5501 29168
rect 5443 29127 5501 29128
rect 5835 29168 5877 29177
rect 5835 29128 5836 29168
rect 5876 29128 5877 29168
rect 5835 29119 5877 29128
rect 79755 29168 79797 29177
rect 79755 29128 79756 29168
rect 79796 29128 79797 29168
rect 79755 29119 79797 29128
rect 80035 29168 80093 29169
rect 80035 29128 80044 29168
rect 80084 29128 80093 29168
rect 80035 29127 80093 29128
rect 81187 29168 81245 29169
rect 81187 29128 81196 29168
rect 81236 29128 81245 29168
rect 81187 29127 81245 29128
rect 82051 29168 82109 29169
rect 82051 29128 82060 29168
rect 82100 29128 82109 29168
rect 82051 29127 82109 29128
rect 79363 29000 79421 29001
rect 79363 28960 79372 29000
rect 79412 28960 79421 29000
rect 79363 28959 79421 28960
rect 3427 28916 3485 28917
rect 3427 28876 3436 28916
rect 3476 28876 3485 28916
rect 3427 28875 3485 28876
rect 576 28748 5952 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 5952 28748
rect 576 28684 5952 28708
rect 74016 28748 83328 28772
rect 74016 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 83328 28748
rect 74016 28684 83328 28708
rect 5155 28580 5213 28581
rect 5155 28540 5164 28580
rect 5204 28540 5213 28580
rect 5155 28539 5213 28540
rect 83203 28580 83261 28581
rect 83203 28540 83212 28580
rect 83252 28540 83261 28580
rect 83203 28539 83261 28540
rect 80611 28496 80669 28497
rect 80611 28456 80620 28496
rect 80660 28456 80669 28496
rect 80611 28455 80669 28456
rect 4483 28328 4541 28329
rect 4483 28288 4492 28328
rect 4532 28288 4541 28328
rect 4483 28287 4541 28288
rect 4779 28328 4821 28337
rect 4779 28288 4780 28328
rect 4820 28288 4821 28328
rect 4779 28279 4821 28288
rect 74179 28328 74237 28329
rect 74179 28288 74188 28328
rect 74228 28288 74237 28328
rect 74179 28287 74237 28288
rect 79939 28328 79997 28329
rect 79939 28288 79948 28328
rect 79988 28288 79997 28328
rect 79939 28287 79997 28288
rect 80235 28328 80277 28337
rect 80235 28288 80236 28328
rect 80276 28288 80277 28328
rect 80235 28279 80277 28288
rect 80331 28328 80373 28337
rect 80331 28288 80332 28328
rect 80372 28288 80373 28328
rect 80331 28279 80373 28288
rect 80811 28328 80853 28337
rect 80811 28288 80812 28328
rect 80852 28288 80853 28328
rect 80811 28279 80853 28288
rect 81187 28328 81245 28329
rect 81187 28288 81196 28328
rect 81236 28288 81245 28328
rect 81187 28287 81245 28288
rect 82051 28328 82109 28329
rect 82051 28288 82060 28328
rect 82100 28288 82109 28328
rect 82051 28287 82109 28288
rect 4875 28244 4917 28253
rect 4875 28204 4876 28244
rect 4916 28204 4917 28244
rect 4875 28195 4917 28204
rect 75819 28160 75861 28169
rect 75819 28120 75820 28160
rect 75860 28120 75861 28160
rect 75819 28111 75861 28120
rect 576 27992 5952 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 5952 27992
rect 576 27928 5952 27952
rect 74016 27992 83328 28016
rect 74016 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 83328 27992
rect 74016 27928 83328 27952
rect 80523 27740 80565 27749
rect 80523 27700 80524 27740
rect 80564 27700 80565 27740
rect 80523 27691 80565 27700
rect 80131 27656 80189 27657
rect 80131 27616 80140 27656
rect 80180 27616 80189 27656
rect 80131 27615 80189 27616
rect 80427 27656 80469 27665
rect 80427 27616 80428 27656
rect 80468 27616 80469 27656
rect 80427 27607 80469 27616
rect 80803 27404 80861 27405
rect 80803 27364 80812 27404
rect 80852 27364 80861 27404
rect 80803 27363 80861 27364
rect 576 27236 5952 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 5952 27236
rect 576 27172 5952 27196
rect 74016 27236 83328 27260
rect 74016 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 83328 27236
rect 74016 27172 83328 27196
rect 83203 27068 83261 27069
rect 83203 27028 83212 27068
rect 83252 27028 83261 27068
rect 83203 27027 83261 27028
rect 79843 26984 79901 26985
rect 79843 26944 79852 26984
rect 79892 26944 79901 26984
rect 79843 26943 79901 26944
rect 80235 26816 80277 26825
rect 80235 26776 80236 26816
rect 80276 26776 80277 26816
rect 80235 26767 80277 26776
rect 80515 26816 80573 26817
rect 80515 26776 80524 26816
rect 80564 26776 80573 26816
rect 80515 26775 80573 26776
rect 80811 26816 80853 26825
rect 80811 26776 80812 26816
rect 80852 26776 80853 26816
rect 80811 26767 80853 26776
rect 81187 26816 81245 26817
rect 81187 26776 81196 26816
rect 81236 26776 81245 26816
rect 81187 26775 81245 26776
rect 82051 26816 82109 26817
rect 82051 26776 82060 26816
rect 82100 26776 82109 26816
rect 82051 26775 82109 26776
rect 80139 26732 80181 26741
rect 80139 26692 80140 26732
rect 80180 26692 80181 26732
rect 80139 26683 80181 26692
rect 576 26480 5952 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 5952 26480
rect 576 26416 5952 26440
rect 74016 26480 83328 26504
rect 74016 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 83328 26480
rect 74016 26416 83328 26440
rect 5827 26312 5885 26313
rect 5827 26272 5836 26312
rect 5876 26272 5885 26312
rect 5827 26271 5885 26272
rect 80235 26228 80277 26237
rect 80235 26188 80236 26228
rect 80276 26188 80277 26228
rect 80235 26179 80277 26188
rect 3435 26144 3477 26153
rect 3435 26104 3436 26144
rect 3476 26104 3477 26144
rect 3435 26095 3477 26104
rect 3811 26144 3869 26145
rect 3811 26104 3820 26144
rect 3860 26104 3869 26144
rect 3811 26103 3869 26104
rect 4675 26144 4733 26145
rect 4675 26104 4684 26144
rect 4724 26104 4733 26144
rect 4675 26103 4733 26104
rect 80611 26144 80669 26145
rect 80611 26104 80620 26144
rect 80660 26104 80669 26144
rect 80611 26103 80669 26104
rect 81475 26144 81533 26145
rect 81475 26104 81484 26144
rect 81524 26104 81533 26144
rect 81475 26103 81533 26104
rect 82627 25976 82685 25977
rect 82627 25936 82636 25976
rect 82676 25936 82685 25976
rect 82627 25935 82685 25936
rect 5827 25892 5885 25893
rect 5827 25852 5836 25892
rect 5876 25852 5885 25892
rect 5827 25851 5885 25852
rect 576 25724 5952 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 5952 25724
rect 576 25660 5952 25684
rect 74016 25724 83328 25748
rect 74016 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 83328 25724
rect 74016 25660 83328 25684
rect 4195 25556 4253 25557
rect 4195 25516 4204 25556
rect 4244 25516 4253 25556
rect 4195 25515 4253 25516
rect 80227 25472 80285 25473
rect 80227 25432 80236 25472
rect 80276 25432 80285 25472
rect 80227 25431 80285 25432
rect 81187 25472 81245 25473
rect 81187 25432 81196 25472
rect 81236 25432 81245 25472
rect 81187 25431 81245 25432
rect 643 25388 701 25389
rect 643 25348 652 25388
rect 692 25348 701 25388
rect 643 25347 701 25348
rect 4491 25304 4533 25313
rect 4491 25264 4492 25304
rect 4532 25264 4533 25304
rect 4491 25255 4533 25264
rect 4587 25304 4629 25313
rect 4587 25264 4588 25304
rect 4628 25264 4629 25304
rect 4587 25255 4629 25264
rect 4867 25304 4925 25305
rect 4867 25264 4876 25304
rect 4916 25264 4925 25304
rect 4867 25263 4925 25264
rect 80619 25304 80661 25313
rect 80619 25264 80620 25304
rect 80660 25264 80661 25304
rect 80619 25255 80661 25264
rect 80899 25304 80957 25305
rect 80899 25264 80908 25304
rect 80948 25264 80957 25304
rect 80899 25263 80957 25264
rect 81483 25304 81525 25313
rect 81483 25264 81484 25304
rect 81524 25264 81525 25304
rect 81483 25255 81525 25264
rect 81579 25304 81621 25313
rect 81579 25264 81580 25304
rect 81620 25264 81621 25304
rect 81579 25255 81621 25264
rect 81859 25304 81917 25305
rect 81859 25264 81868 25304
rect 81908 25264 81917 25304
rect 81859 25263 81917 25264
rect 80523 25220 80565 25229
rect 80523 25180 80524 25220
rect 80564 25180 80565 25220
rect 80523 25171 80565 25180
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 576 24968 5952 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 5952 24968
rect 576 24904 5952 24928
rect 74016 24968 83328 24992
rect 74016 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 83328 24968
rect 74016 24904 83328 24928
rect 843 24800 885 24809
rect 843 24760 844 24800
rect 884 24760 885 24800
rect 843 24751 885 24760
rect 80235 24716 80277 24725
rect 80235 24676 80236 24716
rect 80276 24676 80277 24716
rect 80235 24667 80277 24676
rect 80611 24632 80669 24633
rect 80611 24592 80620 24632
rect 80660 24592 80669 24632
rect 80611 24591 80669 24592
rect 81475 24632 81533 24633
rect 81475 24592 81484 24632
rect 81524 24592 81533 24632
rect 81475 24591 81533 24592
rect 643 24548 701 24549
rect 643 24508 652 24548
rect 692 24508 701 24548
rect 643 24507 701 24508
rect 82635 24548 82677 24557
rect 82635 24508 82636 24548
rect 82676 24508 82677 24548
rect 82635 24499 82677 24508
rect 576 24212 5952 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 5952 24212
rect 576 24148 5952 24172
rect 74016 24212 83328 24236
rect 74016 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 83328 24212
rect 74016 24148 83328 24172
rect 843 24044 885 24053
rect 843 24004 844 24044
rect 884 24004 885 24044
rect 843 23995 885 24004
rect 5827 24044 5885 24045
rect 5827 24004 5836 24044
rect 5876 24004 5885 24044
rect 5827 24003 5885 24004
rect 83203 24044 83261 24045
rect 83203 24004 83212 24044
rect 83252 24004 83261 24044
rect 83203 24003 83261 24004
rect 643 23876 701 23877
rect 643 23836 652 23876
rect 692 23836 701 23876
rect 643 23835 701 23836
rect 3811 23792 3869 23793
rect 3811 23752 3820 23792
rect 3860 23752 3869 23792
rect 3811 23751 3869 23752
rect 4675 23792 4733 23793
rect 4675 23752 4684 23792
rect 4724 23752 4733 23792
rect 4675 23751 4733 23752
rect 80811 23792 80853 23801
rect 80811 23752 80812 23792
rect 80852 23752 80853 23792
rect 80811 23743 80853 23752
rect 81187 23792 81245 23793
rect 81187 23752 81196 23792
rect 81236 23752 81245 23792
rect 81187 23751 81245 23752
rect 82051 23792 82109 23793
rect 82051 23752 82060 23792
rect 82100 23752 82109 23792
rect 82051 23751 82109 23752
rect 3435 23708 3477 23717
rect 3435 23668 3436 23708
rect 3476 23668 3477 23708
rect 3435 23659 3477 23668
rect 576 23456 5952 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 5952 23456
rect 576 23392 5952 23416
rect 74016 23456 83328 23480
rect 74016 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 83328 23456
rect 74016 23392 83328 23416
rect 4203 23330 4245 23339
rect 843 23288 885 23297
rect 843 23248 844 23288
rect 884 23248 885 23288
rect 4203 23290 4204 23330
rect 4244 23290 4245 23330
rect 4203 23281 4245 23290
rect 843 23239 885 23248
rect 4491 23204 4533 23213
rect 4491 23164 4492 23204
rect 4532 23164 4533 23204
rect 4491 23155 4533 23164
rect 3531 23120 3573 23129
rect 3531 23080 3532 23120
rect 3572 23080 3573 23120
rect 3531 23071 3573 23080
rect 3627 23120 3669 23129
rect 3627 23080 3628 23120
rect 3668 23080 3669 23120
rect 3627 23071 3669 23080
rect 3907 23120 3965 23121
rect 3907 23080 3916 23120
rect 3956 23080 3965 23120
rect 3907 23079 3965 23080
rect 4587 23120 4629 23129
rect 4587 23080 4588 23120
rect 4628 23080 4629 23120
rect 4587 23071 4629 23080
rect 4867 23120 4925 23121
rect 4867 23080 4876 23120
rect 4916 23080 4925 23120
rect 4867 23079 4925 23080
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 3235 22868 3293 22869
rect 3235 22828 3244 22868
rect 3284 22828 3293 22868
rect 3235 22827 3293 22828
rect 576 22700 5952 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 5952 22700
rect 576 22636 5952 22660
rect 74016 22700 83328 22724
rect 74016 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 83328 22700
rect 74016 22636 83328 22660
rect 5827 22532 5885 22533
rect 5827 22492 5836 22532
rect 5876 22492 5885 22532
rect 5827 22491 5885 22492
rect 3435 22280 3477 22289
rect 3435 22240 3436 22280
rect 3476 22240 3477 22280
rect 3435 22231 3477 22240
rect 3811 22280 3869 22281
rect 3811 22240 3820 22280
rect 3860 22240 3869 22280
rect 3811 22239 3869 22240
rect 4675 22280 4733 22281
rect 4675 22240 4684 22280
rect 4724 22240 4733 22280
rect 4675 22239 4733 22240
rect 643 22112 701 22113
rect 643 22072 652 22112
rect 692 22072 701 22112
rect 643 22071 701 22072
rect 5827 22112 5885 22113
rect 5827 22072 5836 22112
rect 5876 22072 5885 22112
rect 5827 22071 5885 22072
rect 576 21944 5952 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 5952 21944
rect 576 21880 5952 21904
rect 74016 21944 99360 21968
rect 74016 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 74016 21880 99360 21904
rect 3339 21692 3381 21701
rect 3339 21652 3340 21692
rect 3380 21652 3381 21692
rect 3339 21643 3381 21652
rect 3435 21608 3477 21617
rect 3435 21568 3436 21608
rect 3476 21568 3477 21608
rect 3435 21559 3477 21568
rect 3715 21608 3773 21609
rect 3715 21568 3724 21608
rect 3764 21568 3773 21608
rect 3715 21567 3773 21568
rect 3043 21356 3101 21357
rect 3043 21316 3052 21356
rect 3092 21316 3101 21356
rect 3043 21315 3101 21316
rect 576 21188 5952 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 5952 21188
rect 576 21124 5952 21148
rect 74016 21188 99360 21212
rect 74016 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 74016 21124 99360 21148
rect 5347 21020 5405 21021
rect 5347 20980 5356 21020
rect 5396 20980 5405 21020
rect 5347 20979 5405 20980
rect 84451 21020 84509 21021
rect 84451 20980 84460 21020
rect 84500 20980 84509 21020
rect 84451 20979 84509 20980
rect 81763 20936 81821 20937
rect 81763 20896 81772 20936
rect 81812 20896 81821 20936
rect 81763 20895 81821 20896
rect 2955 20768 2997 20777
rect 2955 20728 2956 20768
rect 2996 20728 2997 20768
rect 2955 20719 2997 20728
rect 3331 20768 3389 20769
rect 3331 20728 3340 20768
rect 3380 20728 3389 20768
rect 3331 20727 3389 20728
rect 4195 20768 4253 20769
rect 4195 20728 4204 20768
rect 4244 20728 4253 20768
rect 4195 20727 4253 20728
rect 81091 20768 81149 20769
rect 81091 20728 81100 20768
rect 81140 20728 81149 20768
rect 81091 20727 81149 20728
rect 81387 20768 81429 20777
rect 81387 20728 81388 20768
rect 81428 20728 81429 20768
rect 81387 20719 81429 20728
rect 81483 20768 81525 20777
rect 81483 20728 81484 20768
rect 81524 20728 81525 20768
rect 81483 20719 81525 20728
rect 82435 20768 82493 20769
rect 82435 20728 82444 20768
rect 82484 20728 82493 20768
rect 82435 20727 82493 20728
rect 83299 20768 83357 20769
rect 83299 20728 83308 20768
rect 83348 20728 83357 20768
rect 83299 20727 83357 20728
rect 82059 20684 82101 20693
rect 82059 20644 82060 20684
rect 82100 20644 82101 20684
rect 82059 20635 82101 20644
rect 643 20600 701 20601
rect 643 20560 652 20600
rect 692 20560 701 20600
rect 643 20559 701 20560
rect 576 20432 5952 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 5952 20432
rect 576 20368 5952 20392
rect 74016 20432 99360 20456
rect 74016 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 74016 20368 99360 20392
rect 643 20264 701 20265
rect 643 20224 652 20264
rect 692 20224 701 20264
rect 643 20223 701 20224
rect 3435 20096 3477 20105
rect 3435 20056 3436 20096
rect 3476 20056 3477 20096
rect 3435 20047 3477 20056
rect 3811 20096 3869 20097
rect 3811 20056 3820 20096
rect 3860 20056 3869 20096
rect 3811 20055 3869 20056
rect 4675 20096 4733 20097
rect 4675 20056 4684 20096
rect 4724 20056 4733 20096
rect 4675 20055 4733 20056
rect 96739 20096 96797 20097
rect 96739 20056 96748 20096
rect 96788 20056 96797 20096
rect 96739 20055 96797 20056
rect 5835 20012 5877 20021
rect 5835 19972 5836 20012
rect 5876 19972 5877 20012
rect 5835 19963 5877 19972
rect 98571 19928 98613 19937
rect 98571 19888 98572 19928
rect 98612 19888 98613 19928
rect 98571 19879 98613 19888
rect 576 19676 5952 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 5952 19676
rect 576 19612 5952 19636
rect 74016 19676 99360 19700
rect 74016 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 74016 19612 99360 19636
rect 3619 19508 3677 19509
rect 3619 19468 3628 19508
rect 3668 19468 3677 19508
rect 3619 19467 3677 19468
rect 2851 19340 2909 19341
rect 2851 19300 2860 19340
rect 2900 19300 2909 19340
rect 2851 19299 2909 19300
rect 3427 19340 3485 19341
rect 3427 19300 3436 19340
rect 3476 19300 3485 19340
rect 3427 19299 3485 19300
rect 3915 19256 3957 19265
rect 3915 19216 3916 19256
rect 3956 19216 3957 19256
rect 3915 19207 3957 19216
rect 4011 19256 4053 19265
rect 4011 19216 4012 19256
rect 4052 19216 4053 19256
rect 4011 19207 4053 19216
rect 4291 19256 4349 19257
rect 4291 19216 4300 19256
rect 4340 19216 4349 19256
rect 4291 19215 4349 19216
rect 643 19088 701 19089
rect 643 19048 652 19088
rect 692 19048 701 19088
rect 643 19047 701 19048
rect 3051 19088 3093 19097
rect 3051 19048 3052 19088
rect 3092 19048 3093 19088
rect 3051 19039 3093 19048
rect 3243 19088 3285 19097
rect 3243 19048 3244 19088
rect 3284 19048 3285 19088
rect 3243 19039 3285 19048
rect 576 18920 5952 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 5952 18920
rect 576 18856 5952 18880
rect 74016 18920 80736 18944
rect 74016 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80736 18920
rect 74016 18856 80736 18880
rect 643 18752 701 18753
rect 643 18712 652 18752
rect 692 18712 701 18752
rect 643 18711 701 18712
rect 2955 18668 2997 18677
rect 2955 18628 2956 18668
rect 2996 18628 2997 18668
rect 2955 18619 2997 18628
rect 2563 18584 2621 18585
rect 2563 18544 2572 18584
rect 2612 18544 2621 18584
rect 2563 18543 2621 18544
rect 2859 18584 2901 18593
rect 2859 18544 2860 18584
rect 2900 18544 2901 18584
rect 2859 18535 2901 18544
rect 3435 18584 3477 18593
rect 3435 18544 3436 18584
rect 3476 18544 3477 18584
rect 3435 18535 3477 18544
rect 3811 18584 3869 18585
rect 3811 18544 3820 18584
rect 3860 18544 3869 18584
rect 3811 18543 3869 18544
rect 4675 18584 4733 18585
rect 4675 18544 4684 18584
rect 4724 18544 4733 18584
rect 4675 18543 4733 18544
rect 2275 18500 2333 18501
rect 2275 18460 2284 18500
rect 2324 18460 2333 18500
rect 2275 18459 2333 18460
rect 5835 18500 5877 18509
rect 5835 18460 5836 18500
rect 5876 18460 5877 18500
rect 5835 18451 5877 18460
rect 3235 18416 3293 18417
rect 3235 18376 3244 18416
rect 3284 18376 3293 18416
rect 3235 18375 3293 18376
rect 2091 18332 2133 18341
rect 2091 18292 2092 18332
rect 2132 18292 2133 18332
rect 2091 18283 2133 18292
rect 576 18164 5952 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 5952 18164
rect 576 18100 5952 18124
rect 74016 18164 80736 18188
rect 74016 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 80736 18164
rect 74016 18100 80736 18124
rect 5059 17912 5117 17913
rect 5059 17872 5068 17912
rect 5108 17872 5117 17912
rect 5059 17871 5117 17872
rect 2467 17828 2525 17829
rect 2467 17788 2476 17828
rect 2516 17788 2525 17828
rect 2467 17787 2525 17788
rect 3043 17744 3101 17745
rect 3043 17704 3052 17744
rect 3092 17704 3101 17744
rect 3043 17703 3101 17704
rect 3907 17744 3965 17745
rect 3907 17704 3916 17744
rect 3956 17704 3965 17744
rect 3907 17703 3965 17704
rect 2667 17660 2709 17669
rect 2667 17620 2668 17660
rect 2708 17620 2709 17660
rect 2667 17611 2709 17620
rect 643 17576 701 17577
rect 643 17536 652 17576
rect 692 17536 701 17576
rect 643 17535 701 17536
rect 2283 17576 2325 17585
rect 2283 17536 2284 17576
rect 2324 17536 2325 17576
rect 2283 17527 2325 17536
rect 576 17408 5952 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 5952 17408
rect 576 17344 5952 17368
rect 74016 17408 80736 17432
rect 74016 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80736 17408
rect 74016 17344 80736 17368
rect 643 17240 701 17241
rect 643 17200 652 17240
rect 692 17200 701 17240
rect 643 17199 701 17200
rect 2667 17156 2709 17165
rect 2667 17116 2668 17156
rect 2708 17116 2709 17156
rect 2667 17107 2709 17116
rect 2275 17072 2333 17073
rect 2275 17032 2284 17072
rect 2324 17032 2333 17072
rect 2275 17031 2333 17032
rect 2571 17072 2613 17081
rect 2571 17032 2572 17072
rect 2612 17032 2613 17072
rect 2571 17023 2613 17032
rect 78219 17072 78261 17081
rect 78219 17032 78220 17072
rect 78260 17032 78261 17072
rect 78219 17023 78261 17032
rect 78595 17072 78653 17073
rect 78595 17032 78604 17072
rect 78644 17032 78653 17072
rect 78595 17031 78653 17032
rect 79459 17072 79517 17073
rect 79459 17032 79468 17072
rect 79508 17032 79517 17072
rect 79459 17031 79517 17032
rect 3235 16988 3293 16989
rect 3235 16948 3244 16988
rect 3284 16948 3293 16988
rect 3235 16947 3293 16948
rect 2947 16904 3005 16905
rect 2947 16864 2956 16904
rect 2996 16864 3005 16904
rect 2947 16863 3005 16864
rect 3435 16820 3477 16829
rect 3435 16780 3436 16820
rect 3476 16780 3477 16820
rect 3435 16771 3477 16780
rect 80611 16820 80669 16821
rect 80611 16780 80620 16820
rect 80660 16780 80669 16820
rect 80611 16779 80669 16780
rect 576 16652 5952 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 5952 16652
rect 576 16588 5952 16612
rect 74016 16652 80736 16676
rect 74016 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 80736 16652
rect 74016 16588 80736 16612
rect 3235 16484 3293 16485
rect 3235 16444 3244 16484
rect 3284 16444 3293 16484
rect 3235 16443 3293 16444
rect 5827 16484 5885 16485
rect 5827 16444 5836 16484
rect 5876 16444 5885 16484
rect 5827 16443 5885 16444
rect 78115 16484 78173 16485
rect 78115 16444 78124 16484
rect 78164 16444 78173 16484
rect 78115 16443 78173 16444
rect 1219 16232 1277 16233
rect 1219 16192 1228 16232
rect 1268 16192 1277 16232
rect 1219 16191 1277 16192
rect 2083 16232 2141 16233
rect 2083 16192 2092 16232
rect 2132 16192 2141 16232
rect 2083 16191 2141 16192
rect 3811 16232 3869 16233
rect 3811 16192 3820 16232
rect 3860 16192 3869 16232
rect 3811 16191 3869 16192
rect 4675 16232 4733 16233
rect 4675 16192 4684 16232
rect 4724 16192 4733 16232
rect 4675 16191 4733 16192
rect 78411 16232 78453 16241
rect 78411 16192 78412 16232
rect 78452 16192 78453 16232
rect 78411 16183 78453 16192
rect 78507 16232 78549 16241
rect 78507 16192 78508 16232
rect 78548 16192 78549 16232
rect 78507 16183 78549 16192
rect 78787 16232 78845 16233
rect 78787 16192 78796 16232
rect 78836 16192 78845 16232
rect 78787 16191 78845 16192
rect 843 16148 885 16157
rect 843 16108 844 16148
rect 884 16108 885 16148
rect 843 16099 885 16108
rect 3435 16148 3477 16157
rect 3435 16108 3436 16148
rect 3476 16108 3477 16148
rect 3435 16099 3477 16108
rect 5827 16064 5885 16065
rect 5827 16024 5836 16064
rect 5876 16024 5885 16064
rect 5827 16023 5885 16024
rect 576 15896 5952 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 5952 15896
rect 576 15832 5952 15856
rect 74016 15896 80736 15920
rect 74016 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80736 15896
rect 74016 15832 80736 15856
rect 643 15728 701 15729
rect 643 15688 652 15728
rect 692 15688 701 15728
rect 643 15687 701 15688
rect 1803 15644 1845 15653
rect 1803 15604 1804 15644
rect 1844 15604 1845 15644
rect 1803 15595 1845 15604
rect 4491 15644 4533 15653
rect 4491 15604 4492 15644
rect 4532 15604 4533 15644
rect 4491 15595 4533 15604
rect 1899 15560 1941 15569
rect 1899 15520 1900 15560
rect 1940 15520 1941 15560
rect 1899 15511 1941 15520
rect 2179 15560 2237 15561
rect 2179 15520 2188 15560
rect 2228 15520 2237 15560
rect 2179 15519 2237 15520
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 4867 15560 4925 15561
rect 4867 15520 4876 15560
rect 4916 15520 4925 15560
rect 4867 15519 4925 15520
rect 1219 15476 1277 15477
rect 1219 15436 1228 15476
rect 1268 15436 1277 15476
rect 1219 15435 1277 15436
rect 1507 15392 1565 15393
rect 1507 15352 1516 15392
rect 1556 15352 1565 15392
rect 1507 15351 1565 15352
rect 4195 15392 4253 15393
rect 4195 15352 4204 15392
rect 4244 15352 4253 15392
rect 4195 15351 4253 15352
rect 1035 15308 1077 15317
rect 1035 15268 1036 15308
rect 1076 15268 1077 15308
rect 1035 15259 1077 15268
rect 576 15140 5952 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 5952 15140
rect 576 15076 5952 15100
rect 74016 15140 80736 15164
rect 74016 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 80736 15140
rect 74016 15076 80736 15100
rect 5827 14972 5885 14973
rect 5827 14932 5836 14972
rect 5876 14932 5885 14972
rect 5827 14931 5885 14932
rect 3235 14888 3293 14889
rect 3235 14848 3244 14888
rect 3284 14848 3293 14888
rect 3235 14847 3293 14848
rect 1219 14720 1277 14721
rect 1219 14680 1228 14720
rect 1268 14680 1277 14720
rect 1219 14679 1277 14680
rect 2083 14720 2141 14721
rect 2083 14680 2092 14720
rect 2132 14680 2141 14720
rect 2083 14679 2141 14680
rect 3811 14720 3869 14721
rect 3811 14680 3820 14720
rect 3860 14680 3869 14720
rect 3811 14679 3869 14680
rect 4675 14720 4733 14721
rect 4675 14680 4684 14720
rect 4724 14680 4733 14720
rect 4675 14679 4733 14680
rect 843 14636 885 14645
rect 843 14596 844 14636
rect 884 14596 885 14636
rect 843 14587 885 14596
rect 3435 14636 3477 14645
rect 3435 14596 3436 14636
rect 3476 14596 3477 14636
rect 3435 14587 3477 14596
rect 576 14384 5952 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 5952 14384
rect 576 14320 5952 14344
rect 74016 14384 80736 14408
rect 74016 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80736 14384
rect 74016 14320 80736 14344
rect 1611 14132 1653 14141
rect 1611 14092 1612 14132
rect 1652 14092 1653 14132
rect 1611 14083 1653 14092
rect 3819 14132 3861 14141
rect 3819 14092 3820 14132
rect 3860 14092 3861 14132
rect 3819 14083 3861 14092
rect 1707 14048 1749 14057
rect 1707 14008 1708 14048
rect 1748 14008 1749 14048
rect 1707 13999 1749 14008
rect 1987 14048 2045 14049
rect 1987 14008 1996 14048
rect 2036 14008 2045 14048
rect 1987 14007 2045 14008
rect 3915 14048 3957 14057
rect 3915 14008 3916 14048
rect 3956 14008 3957 14048
rect 3915 13999 3957 14008
rect 4195 14048 4253 14049
rect 4195 14008 4204 14048
rect 4244 14008 4253 14048
rect 4195 14007 4253 14008
rect 835 13964 893 13965
rect 835 13924 844 13964
rect 884 13924 893 13964
rect 835 13923 893 13924
rect 651 13880 693 13889
rect 651 13840 652 13880
rect 692 13840 693 13880
rect 651 13831 693 13840
rect 1315 13880 1373 13881
rect 1315 13840 1324 13880
rect 1364 13840 1373 13880
rect 1315 13839 1373 13840
rect 3523 13880 3581 13881
rect 3523 13840 3532 13880
rect 3572 13840 3581 13880
rect 3523 13839 3581 13840
rect 576 13628 5952 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 5952 13628
rect 576 13564 5952 13588
rect 74016 13628 80736 13652
rect 74016 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 80736 13628
rect 74016 13564 80736 13588
rect 1219 13208 1277 13209
rect 1219 13168 1228 13208
rect 1268 13168 1277 13208
rect 1219 13167 1277 13168
rect 2083 13208 2141 13209
rect 2083 13168 2092 13208
rect 2132 13168 2141 13208
rect 2083 13167 2141 13168
rect 3811 13208 3869 13209
rect 3811 13168 3820 13208
rect 3860 13168 3869 13208
rect 3811 13167 3869 13168
rect 4675 13208 4733 13209
rect 4675 13168 4684 13208
rect 4724 13168 4733 13208
rect 4675 13167 4733 13168
rect 843 13124 885 13133
rect 843 13084 844 13124
rect 884 13084 885 13124
rect 843 13075 885 13084
rect 3435 13124 3477 13133
rect 3435 13084 3436 13124
rect 3476 13084 3477 13124
rect 3435 13075 3477 13084
rect 3235 13040 3293 13041
rect 3235 13000 3244 13040
rect 3284 13000 3293 13040
rect 3235 12999 3293 13000
rect 5827 13040 5885 13041
rect 5827 13000 5836 13040
rect 5876 13000 5885 13040
rect 5827 12999 5885 13000
rect 576 12872 5952 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 5952 12872
rect 576 12808 5952 12832
rect 74016 12872 80736 12896
rect 74016 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80736 12872
rect 74016 12808 80736 12832
rect 651 12704 693 12713
rect 651 12664 652 12704
rect 692 12664 693 12704
rect 651 12655 693 12664
rect 3819 12620 3861 12629
rect 3819 12580 3820 12620
rect 3860 12580 3861 12620
rect 3819 12571 3861 12580
rect 1707 12536 1749 12545
rect 1707 12496 1708 12536
rect 1748 12496 1749 12536
rect 1707 12487 1749 12496
rect 1803 12536 1845 12545
rect 1803 12496 1804 12536
rect 1844 12496 1845 12536
rect 1803 12487 1845 12496
rect 2083 12536 2141 12537
rect 2083 12496 2092 12536
rect 2132 12496 2141 12536
rect 2083 12495 2141 12496
rect 3915 12536 3957 12545
rect 3915 12496 3916 12536
rect 3956 12496 3957 12536
rect 3915 12487 3957 12496
rect 4195 12536 4253 12537
rect 4195 12496 4204 12536
rect 4244 12496 4253 12536
rect 4195 12495 4253 12496
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 1219 12452 1277 12453
rect 1219 12412 1228 12452
rect 1268 12412 1277 12452
rect 1219 12411 1277 12412
rect 1035 12368 1077 12377
rect 1035 12328 1036 12368
rect 1076 12328 1077 12368
rect 1035 12319 1077 12328
rect 1411 12368 1469 12369
rect 1411 12328 1420 12368
rect 1460 12328 1469 12368
rect 1411 12327 1469 12328
rect 3523 12368 3581 12369
rect 3523 12328 3532 12368
rect 3572 12328 3581 12368
rect 3523 12327 3581 12328
rect 576 12116 5952 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 5952 12116
rect 576 12052 5952 12076
rect 74016 12116 80736 12140
rect 74016 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 80736 12116
rect 74016 12052 80736 12076
rect 5827 11948 5885 11949
rect 5827 11908 5836 11948
rect 5876 11908 5885 11948
rect 5827 11907 5885 11908
rect 3235 11864 3293 11865
rect 3235 11824 3244 11864
rect 3284 11824 3293 11864
rect 3235 11823 3293 11824
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 2859 11738 2901 11747
rect 2859 11698 2860 11738
rect 2900 11698 2901 11738
rect 2563 11696 2621 11697
rect 2563 11656 2572 11696
rect 2612 11656 2621 11696
rect 2859 11689 2901 11698
rect 2955 11696 2997 11705
rect 2563 11655 2621 11656
rect 2955 11656 2956 11696
rect 2996 11656 2997 11696
rect 2955 11647 2997 11656
rect 3435 11696 3477 11705
rect 3435 11656 3436 11696
rect 3476 11656 3477 11696
rect 3435 11647 3477 11656
rect 3811 11696 3869 11697
rect 3811 11656 3820 11696
rect 3860 11656 3869 11696
rect 3811 11655 3869 11656
rect 4675 11696 4733 11697
rect 4675 11656 4684 11696
rect 4724 11656 4733 11696
rect 4675 11655 4733 11656
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 576 11360 5952 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 5952 11360
rect 576 11296 5952 11320
rect 74016 11360 80736 11384
rect 74016 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80736 11360
rect 74016 11296 80736 11320
rect 4867 11192 4925 11193
rect 4867 11152 4876 11192
rect 4916 11152 4925 11192
rect 4867 11151 4925 11152
rect 2475 11024 2517 11033
rect 2475 10984 2476 11024
rect 2516 10984 2517 11024
rect 2475 10975 2517 10984
rect 2907 11024 2949 11033
rect 2907 10984 2908 11024
rect 2948 10984 2949 11024
rect 2907 10975 2949 10984
rect 3715 11024 3773 11025
rect 3715 10984 3724 11024
rect 3764 10984 3773 11024
rect 3715 10983 3773 10984
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 576 10604 5952 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 5952 10604
rect 576 10540 5952 10564
rect 74016 10604 80736 10628
rect 74016 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 80736 10604
rect 74016 10540 80736 10564
rect 2275 10436 2333 10437
rect 2275 10396 2284 10436
rect 2324 10396 2333 10436
rect 2275 10395 2333 10396
rect 3907 10352 3965 10353
rect 3907 10312 3916 10352
rect 3956 10312 3965 10352
rect 3907 10311 3965 10312
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 2571 10184 2613 10193
rect 2571 10144 2572 10184
rect 2612 10144 2613 10184
rect 2571 10135 2613 10144
rect 2667 10184 2709 10193
rect 2667 10144 2668 10184
rect 2708 10144 2709 10184
rect 2667 10135 2709 10144
rect 2947 10184 3005 10185
rect 2947 10144 2956 10184
rect 2996 10144 3005 10184
rect 2947 10143 3005 10144
rect 4299 10184 4341 10193
rect 4299 10144 4300 10184
rect 4340 10144 4341 10184
rect 4299 10135 4341 10144
rect 4579 10184 4637 10185
rect 4579 10144 4588 10184
rect 4628 10144 4637 10184
rect 4579 10143 4637 10144
rect 4203 10100 4245 10109
rect 4203 10060 4204 10100
rect 4244 10060 4245 10100
rect 4203 10051 4245 10060
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 576 9848 5952 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 5952 9848
rect 576 9784 5952 9808
rect 74016 9848 80736 9872
rect 74016 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80736 9848
rect 74016 9784 80736 9808
rect 5827 9680 5885 9681
rect 5827 9640 5836 9680
rect 5876 9640 5885 9680
rect 5827 9639 5885 9640
rect 3435 9596 3477 9605
rect 3435 9556 3436 9596
rect 3476 9556 3477 9596
rect 3435 9547 3477 9556
rect 3811 9512 3869 9513
rect 3811 9472 3820 9512
rect 3860 9472 3869 9512
rect 3811 9471 3869 9472
rect 4675 9512 4733 9513
rect 4675 9472 4684 9512
rect 4724 9472 4733 9512
rect 4675 9471 4733 9472
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 651 9260 693 9269
rect 651 9220 652 9260
rect 692 9220 693 9260
rect 651 9211 693 9220
rect 5827 9260 5885 9261
rect 5827 9220 5836 9260
rect 5876 9220 5885 9260
rect 5827 9219 5885 9220
rect 576 9092 5952 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 5952 9092
rect 576 9028 5952 9052
rect 74016 9092 80736 9116
rect 74016 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 80736 9092
rect 74016 9028 80736 9052
rect 643 8504 701 8505
rect 643 8464 652 8504
rect 692 8464 701 8504
rect 643 8463 701 8464
rect 576 8336 5952 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 5952 8336
rect 576 8272 5952 8296
rect 74016 8336 80736 8360
rect 74016 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80736 8336
rect 74016 8272 80736 8296
rect 643 8168 701 8169
rect 643 8128 652 8168
rect 692 8128 701 8168
rect 643 8127 701 8128
rect 5827 8168 5885 8169
rect 5827 8128 5836 8168
rect 5876 8128 5885 8168
rect 5827 8127 5885 8128
rect 3435 8000 3477 8009
rect 3435 7960 3436 8000
rect 3476 7960 3477 8000
rect 3435 7951 3477 7960
rect 3811 8000 3869 8001
rect 3811 7960 3820 8000
rect 3860 7960 3869 8000
rect 3811 7959 3869 7960
rect 4675 8000 4733 8001
rect 4675 7960 4684 8000
rect 4724 7960 4733 8000
rect 4675 7959 4733 7960
rect 576 7580 5952 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 5952 7580
rect 576 7516 5952 7540
rect 74016 7580 80736 7604
rect 74016 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 80736 7580
rect 74016 7516 80736 7540
rect 4291 7412 4349 7413
rect 4291 7372 4300 7412
rect 4340 7372 4349 7412
rect 4291 7371 4349 7372
rect 4587 7160 4629 7169
rect 4587 7120 4588 7160
rect 4628 7120 4629 7160
rect 4587 7111 4629 7120
rect 4683 7160 4725 7169
rect 4683 7120 4684 7160
rect 4724 7120 4725 7160
rect 4683 7111 4725 7120
rect 4963 7160 5021 7161
rect 4963 7120 4972 7160
rect 5012 7120 5021 7160
rect 4963 7119 5021 7120
rect 643 6992 701 6993
rect 643 6952 652 6992
rect 692 6952 701 6992
rect 643 6951 701 6952
rect 576 6824 5952 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 5952 6824
rect 576 6760 5952 6784
rect 74016 6824 80736 6848
rect 74016 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80736 6824
rect 74016 6760 80736 6784
rect 80523 6656 80565 6665
rect 80523 6616 80524 6656
rect 80564 6616 80565 6656
rect 80523 6607 80565 6616
rect 78499 6488 78557 6489
rect 78499 6448 78508 6488
rect 78548 6448 78557 6488
rect 78499 6447 78557 6448
rect 576 6068 5952 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 5952 6068
rect 576 6004 5952 6028
rect 74016 6068 80736 6092
rect 74016 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 80736 6068
rect 74016 6004 80736 6028
rect 643 5480 701 5481
rect 643 5440 652 5480
rect 692 5440 701 5480
rect 643 5439 701 5440
rect 576 5312 80736 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80736 5312
rect 576 5248 80736 5272
rect 643 5144 701 5145
rect 643 5104 652 5144
rect 692 5104 701 5144
rect 643 5103 701 5104
rect 21571 5144 21629 5145
rect 21571 5104 21580 5144
rect 21620 5104 21629 5144
rect 21571 5103 21629 5104
rect 25707 5144 25749 5153
rect 25707 5104 25708 5144
rect 25748 5104 25749 5144
rect 25707 5095 25749 5104
rect 35875 5144 35933 5145
rect 35875 5104 35884 5144
rect 35924 5104 35933 5144
rect 35875 5103 35933 5104
rect 39435 5144 39477 5153
rect 39435 5104 39436 5144
rect 39476 5104 39477 5144
rect 39435 5095 39477 5104
rect 44523 5144 44565 5153
rect 44523 5104 44524 5144
rect 44564 5104 44565 5144
rect 44523 5095 44565 5104
rect 49987 5144 50045 5145
rect 49987 5104 49996 5144
rect 50036 5104 50045 5144
rect 49987 5103 50045 5104
rect 17547 5060 17589 5069
rect 17547 5020 17548 5060
rect 17588 5020 17589 5060
rect 17547 5011 17589 5020
rect 18699 5060 18741 5069
rect 18699 5020 18700 5060
rect 18740 5020 18741 5060
rect 18699 5011 18741 5020
rect 23307 5060 23349 5069
rect 23307 5020 23308 5060
rect 23348 5020 23349 5060
rect 23307 5011 23349 5020
rect 24651 5060 24693 5069
rect 24651 5020 24652 5060
rect 24692 5020 24693 5060
rect 24651 5011 24693 5020
rect 31755 5060 31797 5069
rect 31755 5020 31756 5060
rect 31796 5020 31797 5060
rect 31755 5011 31797 5020
rect 46347 5060 46389 5069
rect 46347 5020 46348 5060
rect 46388 5020 46389 5060
rect 46347 5011 46389 5020
rect 49419 5060 49461 5069
rect 49419 5020 49420 5060
rect 49460 5020 49461 5060
rect 49419 5011 49461 5020
rect 17643 4976 17685 4985
rect 17643 4936 17644 4976
rect 17684 4936 17685 4976
rect 17643 4927 17685 4936
rect 17923 4976 17981 4977
rect 17923 4936 17932 4976
rect 17972 4936 17981 4976
rect 17923 4935 17981 4936
rect 18307 4976 18365 4977
rect 18307 4936 18316 4976
rect 18356 4936 18365 4976
rect 18307 4935 18365 4936
rect 18603 4976 18645 4985
rect 18603 4936 18604 4976
rect 18644 4936 18645 4976
rect 18603 4927 18645 4936
rect 19179 4976 19221 4985
rect 19179 4936 19180 4976
rect 19220 4936 19221 4976
rect 19179 4927 19221 4936
rect 19555 4976 19613 4977
rect 19555 4936 19564 4976
rect 19604 4936 19613 4976
rect 19555 4935 19613 4936
rect 20419 4976 20477 4977
rect 20419 4936 20428 4976
rect 20468 4936 20477 4976
rect 20419 4935 20477 4936
rect 22915 4976 22973 4977
rect 22915 4936 22924 4976
rect 22964 4936 22973 4976
rect 22915 4935 22973 4936
rect 23211 4976 23253 4985
rect 23211 4936 23212 4976
rect 23252 4936 23253 4976
rect 23211 4927 23253 4936
rect 24747 4976 24789 4985
rect 24747 4936 24748 4976
rect 24788 4936 24789 4976
rect 24747 4927 24789 4936
rect 25027 4976 25085 4977
rect 25027 4936 25036 4976
rect 25076 4936 25085 4976
rect 25027 4935 25085 4936
rect 31651 4976 31709 4977
rect 31651 4936 31660 4976
rect 31700 4936 31709 4976
rect 31651 4935 31709 4936
rect 31851 4976 31893 4985
rect 31851 4936 31852 4976
rect 31892 4936 31893 4976
rect 31851 4927 31893 4936
rect 32707 4976 32765 4977
rect 32707 4936 32716 4976
rect 32756 4936 32765 4976
rect 32707 4935 32765 4936
rect 32907 4976 32949 4985
rect 32907 4936 32908 4976
rect 32948 4936 32949 4976
rect 32907 4927 32949 4936
rect 33091 4976 33149 4977
rect 33091 4936 33100 4976
rect 33140 4936 33149 4976
rect 33091 4935 33149 4936
rect 33483 4976 33525 4985
rect 33483 4936 33484 4976
rect 33524 4936 33525 4976
rect 33483 4927 33525 4936
rect 35011 4976 35069 4977
rect 35011 4936 35020 4976
rect 35060 4936 35069 4976
rect 35011 4935 35069 4936
rect 35115 4976 35157 4985
rect 35115 4936 35116 4976
rect 35156 4936 35157 4976
rect 35115 4927 35157 4936
rect 35211 4976 35253 4985
rect 35211 4936 35212 4976
rect 35252 4936 35253 4976
rect 35211 4927 35253 4936
rect 35403 4976 35445 4985
rect 35403 4936 35404 4976
rect 35444 4936 35445 4976
rect 35403 4927 35445 4936
rect 35499 4976 35541 4985
rect 35499 4936 35500 4976
rect 35540 4936 35541 4976
rect 35499 4927 35541 4936
rect 35595 4976 35637 4985
rect 35595 4936 35596 4976
rect 35636 4936 35637 4976
rect 35595 4927 35637 4936
rect 35691 4976 35733 4985
rect 35691 4936 35692 4976
rect 35732 4936 35733 4976
rect 35691 4927 35733 4936
rect 36075 4976 36117 4985
rect 36075 4936 36076 4976
rect 36116 4936 36117 4976
rect 36075 4927 36117 4936
rect 36171 4976 36213 4985
rect 36171 4936 36172 4976
rect 36212 4936 36213 4976
rect 36171 4927 36213 4936
rect 37603 4976 37661 4977
rect 37603 4936 37612 4976
rect 37652 4936 37661 4976
rect 37603 4935 37661 4936
rect 37995 4976 38037 4985
rect 37995 4936 37996 4976
rect 38036 4936 38037 4976
rect 40099 4976 40157 4977
rect 37995 4927 38037 4936
rect 39627 4962 39669 4971
rect 39627 4922 39628 4962
rect 39668 4922 39669 4962
rect 40099 4936 40108 4976
rect 40148 4936 40157 4976
rect 40099 4935 40157 4936
rect 40587 4976 40629 4985
rect 40587 4936 40588 4976
rect 40628 4936 40629 4976
rect 40587 4927 40629 4936
rect 41067 4976 41109 4985
rect 41067 4936 41068 4976
rect 41108 4936 41109 4976
rect 41067 4927 41109 4936
rect 41163 4976 41205 4985
rect 41163 4936 41164 4976
rect 41204 4936 41205 4976
rect 41163 4927 41205 4936
rect 42883 4976 42941 4977
rect 42883 4936 42892 4976
rect 42932 4936 42941 4976
rect 42883 4935 42941 4936
rect 46443 4976 46485 4985
rect 46443 4936 46444 4976
rect 46484 4936 46485 4976
rect 46443 4927 46485 4936
rect 46723 4976 46781 4977
rect 46723 4936 46732 4976
rect 46772 4936 46781 4976
rect 46723 4935 46781 4936
rect 49323 4976 49365 4985
rect 49323 4936 49324 4976
rect 49364 4936 49365 4976
rect 49323 4927 49365 4936
rect 49507 4976 49565 4977
rect 49507 4936 49516 4976
rect 49556 4936 49565 4976
rect 49507 4935 49565 4936
rect 49891 4976 49949 4977
rect 49891 4936 49900 4976
rect 49940 4936 49949 4976
rect 49891 4935 49949 4936
rect 52195 4976 52253 4977
rect 52195 4936 52204 4976
rect 52244 4936 52253 4976
rect 52195 4935 52253 4936
rect 52491 4976 52533 4985
rect 52491 4936 52492 4976
rect 52532 4936 52533 4976
rect 52491 4927 52533 4936
rect 52587 4976 52629 4985
rect 52587 4936 52588 4976
rect 52628 4936 52629 4976
rect 52587 4927 52629 4936
rect 39627 4913 39669 4922
rect 22435 4892 22493 4893
rect 22435 4852 22444 4892
rect 22484 4852 22493 4892
rect 22435 4851 22493 4852
rect 25891 4892 25949 4893
rect 25891 4852 25900 4892
rect 25940 4852 25949 4892
rect 25891 4851 25949 4852
rect 26275 4892 26333 4893
rect 26275 4852 26284 4892
rect 26324 4852 26333 4892
rect 26275 4851 26333 4852
rect 33195 4892 33237 4901
rect 33195 4852 33196 4892
rect 33236 4852 33237 4892
rect 33195 4843 33237 4852
rect 33387 4892 33429 4901
rect 33387 4852 33388 4892
rect 33428 4852 33429 4892
rect 33387 4843 33429 4852
rect 37707 4892 37749 4901
rect 37707 4852 37708 4892
rect 37748 4852 37749 4892
rect 37707 4843 37749 4852
rect 37899 4892 37941 4901
rect 37899 4852 37900 4892
rect 37940 4852 37941 4892
rect 37899 4843 37941 4852
rect 40683 4892 40725 4901
rect 40683 4852 40684 4892
rect 40724 4852 40725 4892
rect 40683 4843 40725 4852
rect 42403 4892 42461 4893
rect 42403 4852 42412 4892
rect 42452 4852 42461 4892
rect 42403 4851 42461 4852
rect 45187 4892 45245 4893
rect 45187 4852 45196 4892
rect 45236 4852 45245 4892
rect 45187 4851 45245 4852
rect 18979 4808 19037 4809
rect 18979 4768 18988 4808
rect 19028 4768 19037 4808
rect 18979 4767 19037 4768
rect 32811 4808 32853 4817
rect 32811 4768 32812 4808
rect 32852 4768 32853 4808
rect 32811 4759 32853 4768
rect 33291 4808 33333 4817
rect 33291 4768 33292 4808
rect 33332 4768 33333 4808
rect 33291 4759 33333 4768
rect 37803 4808 37845 4817
rect 37803 4768 37804 4808
rect 37844 4768 37845 4808
rect 37803 4759 37845 4768
rect 39243 4808 39285 4817
rect 39243 4768 39244 4808
rect 39284 4768 39285 4808
rect 39243 4759 39285 4768
rect 22635 4724 22677 4733
rect 22635 4684 22636 4724
rect 22676 4684 22677 4724
rect 17251 4682 17309 4683
rect 17251 4642 17260 4682
rect 17300 4642 17309 4682
rect 22635 4675 22677 4684
rect 23587 4724 23645 4725
rect 23587 4684 23596 4724
rect 23636 4684 23645 4724
rect 23587 4683 23645 4684
rect 24355 4724 24413 4725
rect 24355 4684 24364 4724
rect 24404 4684 24413 4724
rect 24355 4683 24413 4684
rect 25707 4724 25749 4733
rect 25707 4684 25708 4724
rect 25748 4684 25749 4724
rect 25707 4675 25749 4684
rect 26091 4724 26133 4733
rect 26091 4684 26092 4724
rect 26132 4684 26133 4724
rect 26091 4675 26133 4684
rect 42219 4724 42261 4733
rect 42219 4684 42220 4724
rect 42260 4684 42261 4724
rect 42219 4675 42261 4684
rect 45387 4724 45429 4733
rect 45387 4684 45388 4724
rect 45428 4684 45429 4724
rect 45387 4675 45429 4684
rect 46051 4724 46109 4725
rect 46051 4684 46060 4724
rect 46100 4684 46109 4724
rect 46051 4683 46109 4684
rect 49699 4724 49757 4725
rect 49699 4684 49708 4724
rect 49748 4684 49757 4724
rect 49699 4683 49757 4684
rect 52867 4724 52925 4725
rect 52867 4684 52876 4724
rect 52916 4684 52925 4724
rect 52867 4683 52925 4684
rect 17251 4641 17309 4642
rect 576 4556 80736 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 80736 4556
rect 576 4492 80736 4516
rect 21099 4304 21141 4313
rect 21099 4264 21100 4304
rect 21140 4264 21141 4304
rect 21099 4255 21141 4264
rect 31851 4304 31893 4313
rect 31851 4264 31852 4304
rect 31892 4264 31893 4304
rect 31851 4255 31893 4264
rect 32419 4304 32477 4305
rect 32419 4264 32428 4304
rect 32468 4264 32477 4304
rect 32419 4263 32477 4264
rect 35787 4304 35829 4313
rect 35787 4264 35788 4304
rect 35828 4264 35829 4304
rect 35787 4255 35829 4264
rect 36939 4304 36981 4313
rect 36939 4264 36940 4304
rect 36980 4264 36981 4304
rect 36939 4255 36981 4264
rect 42595 4304 42653 4305
rect 42595 4264 42604 4304
rect 42644 4264 42653 4304
rect 42595 4263 42653 4264
rect 48355 4304 48413 4305
rect 48355 4264 48364 4304
rect 48404 4264 48413 4304
rect 48355 4263 48413 4264
rect 19275 4220 19317 4229
rect 19275 4180 19276 4220
rect 19316 4180 19317 4220
rect 19275 4171 19317 4180
rect 20899 4220 20957 4221
rect 20899 4180 20908 4220
rect 20948 4180 20957 4220
rect 20899 4179 20957 4180
rect 27147 4220 27189 4229
rect 27147 4180 27148 4220
rect 27188 4180 27189 4220
rect 27147 4171 27189 4180
rect 31755 4220 31797 4229
rect 31755 4180 31756 4220
rect 31796 4180 31797 4220
rect 31755 4171 31797 4180
rect 31947 4220 31989 4229
rect 31947 4180 31948 4220
rect 31988 4180 31989 4220
rect 31947 4171 31989 4180
rect 36843 4220 36885 4229
rect 36843 4180 36844 4220
rect 36884 4180 36885 4220
rect 36843 4171 36885 4180
rect 37035 4220 37077 4229
rect 37035 4180 37036 4220
rect 37076 4180 37077 4220
rect 37035 4171 37077 4180
rect 37611 4220 37653 4229
rect 37611 4180 37612 4220
rect 37652 4180 37653 4220
rect 37611 4171 37653 4180
rect 45195 4220 45237 4229
rect 45195 4180 45196 4220
rect 45236 4180 45237 4220
rect 45195 4171 45237 4180
rect 16875 4136 16917 4145
rect 16875 4096 16876 4136
rect 16916 4096 16917 4136
rect 18115 4136 18173 4137
rect 16875 4087 16917 4096
rect 17251 4123 17309 4124
rect 17251 4083 17260 4123
rect 17300 4083 17309 4123
rect 18115 4096 18124 4136
rect 18164 4096 18173 4136
rect 18115 4095 18173 4096
rect 21667 4136 21725 4137
rect 21667 4096 21676 4136
rect 21716 4096 21725 4136
rect 21667 4095 21725 4096
rect 22531 4136 22589 4137
rect 22531 4096 22540 4136
rect 22580 4096 22589 4136
rect 22531 4095 22589 4096
rect 24747 4136 24789 4145
rect 24747 4096 24748 4136
rect 24788 4096 24789 4136
rect 24747 4087 24789 4096
rect 25123 4136 25181 4137
rect 25123 4096 25132 4136
rect 25172 4096 25181 4136
rect 25123 4095 25181 4096
rect 25987 4136 26045 4137
rect 25987 4096 25996 4136
rect 26036 4096 26045 4136
rect 25987 4095 26045 4096
rect 27715 4136 27773 4137
rect 27715 4096 27724 4136
rect 27764 4096 27773 4136
rect 27715 4095 27773 4096
rect 28579 4136 28637 4137
rect 28579 4096 28588 4136
rect 28628 4096 28637 4136
rect 28579 4095 28637 4096
rect 29923 4136 29981 4137
rect 29923 4096 29932 4136
rect 29972 4096 29981 4136
rect 29923 4095 29981 4096
rect 31171 4136 31229 4137
rect 31171 4096 31180 4136
rect 31220 4096 31229 4136
rect 31171 4095 31229 4096
rect 31651 4136 31709 4137
rect 31651 4096 31660 4136
rect 31700 4096 31709 4136
rect 31651 4095 31709 4096
rect 32043 4136 32085 4145
rect 32043 4096 32044 4136
rect 32084 4096 32085 4136
rect 32043 4087 32085 4096
rect 32611 4136 32669 4137
rect 32611 4096 32620 4136
rect 32660 4096 32669 4136
rect 32611 4095 32669 4096
rect 34635 4136 34677 4145
rect 34635 4096 34636 4136
rect 34676 4096 34677 4136
rect 34635 4087 34677 4096
rect 34731 4136 34773 4145
rect 34731 4096 34732 4136
rect 34772 4096 34773 4136
rect 34731 4087 34773 4096
rect 34827 4136 34869 4145
rect 34827 4096 34828 4136
rect 34868 4096 34869 4136
rect 34827 4087 34869 4096
rect 34923 4136 34965 4145
rect 34923 4096 34924 4136
rect 34964 4096 34965 4136
rect 34923 4087 34965 4096
rect 35595 4136 35637 4145
rect 35595 4096 35596 4136
rect 35636 4096 35637 4136
rect 35595 4087 35637 4096
rect 35787 4136 35829 4145
rect 35787 4096 35788 4136
rect 35828 4096 35829 4136
rect 35787 4087 35829 4096
rect 35979 4136 36021 4145
rect 35979 4096 35980 4136
rect 36020 4096 36021 4136
rect 35979 4087 36021 4096
rect 36171 4136 36213 4145
rect 36171 4096 36172 4136
rect 36212 4096 36213 4136
rect 36171 4087 36213 4096
rect 36259 4136 36317 4137
rect 36259 4096 36268 4136
rect 36308 4096 36317 4136
rect 36259 4095 36317 4096
rect 36739 4136 36797 4137
rect 36739 4096 36748 4136
rect 36788 4096 36797 4136
rect 36739 4095 36797 4096
rect 37131 4136 37173 4145
rect 37131 4096 37132 4136
rect 37172 4096 37173 4136
rect 37131 4087 37173 4096
rect 37515 4136 37557 4145
rect 37515 4096 37516 4136
rect 37556 4096 37557 4136
rect 37515 4087 37557 4096
rect 37707 4136 37749 4145
rect 37707 4096 37708 4136
rect 37748 4096 37749 4136
rect 37707 4087 37749 4096
rect 38859 4136 38901 4145
rect 38859 4096 38860 4136
rect 38900 4096 38901 4136
rect 38859 4087 38901 4096
rect 39147 4136 39189 4145
rect 39147 4096 39148 4136
rect 39188 4096 39189 4136
rect 39147 4087 39189 4096
rect 41923 4136 41981 4137
rect 41923 4096 41932 4136
rect 41972 4096 41981 4136
rect 41923 4095 41981 4096
rect 42219 4136 42261 4145
rect 42219 4096 42220 4136
rect 42260 4096 42261 4136
rect 42219 4087 42261 4096
rect 42315 4136 42357 4145
rect 42315 4096 42316 4136
rect 42356 4096 42357 4136
rect 42315 4087 42357 4096
rect 42795 4136 42837 4145
rect 42795 4096 42796 4136
rect 42836 4096 42837 4136
rect 42795 4087 42837 4096
rect 43171 4136 43229 4137
rect 43171 4096 43180 4136
rect 43220 4096 43229 4136
rect 43171 4095 43229 4096
rect 44035 4136 44093 4137
rect 44035 4096 44044 4136
rect 44084 4096 44093 4136
rect 44035 4095 44093 4096
rect 45963 4136 46005 4145
rect 45963 4096 45964 4136
rect 46004 4096 46005 4136
rect 45963 4087 46005 4096
rect 46339 4136 46397 4137
rect 46339 4096 46348 4136
rect 46388 4096 46397 4136
rect 46339 4095 46397 4096
rect 47203 4136 47261 4137
rect 47203 4096 47212 4136
rect 47252 4096 47261 4136
rect 47203 4095 47261 4096
rect 48931 4136 48989 4137
rect 48931 4096 48940 4136
rect 48980 4096 48989 4136
rect 48931 4095 48989 4096
rect 49795 4136 49853 4137
rect 49795 4096 49804 4136
rect 49844 4096 49853 4136
rect 49795 4095 49853 4096
rect 51523 4136 51581 4137
rect 51523 4096 51532 4136
rect 51572 4096 51581 4136
rect 51523 4095 51581 4096
rect 52387 4136 52445 4137
rect 52387 4096 52396 4136
rect 52436 4096 52445 4136
rect 52387 4095 52445 4096
rect 17251 4082 17309 4083
rect 21291 4052 21333 4061
rect 21291 4012 21292 4052
rect 21332 4012 21333 4052
rect 21291 4003 21333 4012
rect 27339 4052 27381 4061
rect 27339 4012 27340 4052
rect 27380 4012 27381 4052
rect 27339 4003 27381 4012
rect 31371 4052 31413 4061
rect 31371 4012 31372 4052
rect 31412 4012 31413 4052
rect 31371 4003 31413 4012
rect 36075 4052 36117 4061
rect 36075 4012 36076 4052
rect 36116 4012 36117 4052
rect 36075 4003 36117 4012
rect 48555 4052 48597 4061
rect 48555 4012 48556 4052
rect 48596 4012 48597 4052
rect 48555 4003 48597 4012
rect 51147 4052 51189 4061
rect 51147 4012 51148 4052
rect 51188 4012 51189 4052
rect 51147 4003 51189 4012
rect 643 3968 701 3969
rect 643 3928 652 3968
rect 692 3928 701 3968
rect 643 3927 701 3928
rect 23683 3968 23741 3969
rect 23683 3928 23692 3968
rect 23732 3928 23741 3968
rect 23683 3927 23741 3928
rect 29731 3968 29789 3969
rect 29731 3928 29740 3968
rect 29780 3928 29789 3968
rect 29731 3927 29789 3928
rect 32707 3968 32765 3969
rect 32707 3928 32716 3968
rect 32756 3928 32765 3968
rect 32707 3927 32765 3928
rect 39051 3968 39093 3977
rect 39051 3928 39052 3968
rect 39092 3928 39093 3968
rect 39051 3919 39093 3928
rect 50947 3968 51005 3969
rect 50947 3928 50956 3968
rect 50996 3928 51005 3968
rect 50947 3927 51005 3928
rect 53539 3968 53597 3969
rect 53539 3928 53548 3968
rect 53588 3928 53597 3968
rect 53539 3927 53597 3928
rect 576 3800 80736 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80736 3800
rect 576 3736 80736 3760
rect 643 3632 701 3633
rect 643 3592 652 3632
rect 692 3592 701 3632
rect 643 3591 701 3592
rect 25699 3632 25757 3633
rect 25699 3592 25708 3632
rect 25748 3592 25757 3632
rect 25699 3591 25757 3592
rect 32715 3632 32757 3641
rect 32715 3592 32716 3632
rect 32756 3592 32757 3632
rect 32715 3583 32757 3592
rect 42883 3632 42941 3633
rect 42883 3592 42892 3632
rect 42932 3592 42941 3632
rect 42883 3591 42941 3592
rect 44707 3632 44765 3633
rect 44707 3592 44716 3632
rect 44756 3592 44765 3632
rect 44707 3591 44765 3592
rect 49027 3632 49085 3633
rect 49027 3592 49036 3632
rect 49076 3592 49085 3632
rect 49027 3591 49085 3592
rect 49315 3632 49373 3633
rect 49315 3592 49324 3632
rect 49364 3592 49373 3632
rect 49315 3591 49373 3592
rect 49507 3632 49565 3633
rect 49507 3592 49516 3632
rect 49556 3592 49565 3632
rect 49507 3591 49565 3592
rect 49795 3632 49853 3633
rect 49795 3592 49804 3632
rect 49844 3592 49853 3632
rect 49795 3591 49853 3592
rect 55075 3632 55133 3633
rect 55075 3592 55084 3632
rect 55124 3592 55133 3632
rect 55075 3591 55133 3592
rect 21579 3548 21621 3557
rect 21579 3508 21580 3548
rect 21620 3508 21621 3548
rect 21579 3499 21621 3508
rect 23307 3548 23349 3557
rect 23307 3508 23308 3548
rect 23348 3508 23349 3548
rect 23307 3499 23349 3508
rect 27243 3548 27285 3557
rect 27243 3508 27244 3548
rect 27284 3508 27285 3548
rect 27243 3499 27285 3508
rect 33867 3548 33909 3557
rect 33867 3508 33868 3548
rect 33908 3508 33909 3548
rect 27339 3491 27381 3500
rect 33867 3499 33909 3508
rect 35883 3548 35925 3557
rect 35883 3508 35884 3548
rect 35924 3508 35925 3548
rect 35883 3499 35925 3508
rect 40011 3548 40053 3557
rect 40011 3508 40012 3548
rect 40052 3508 40053 3548
rect 40011 3499 40053 3508
rect 44235 3548 44277 3557
rect 44235 3508 44236 3548
rect 44276 3508 44277 3548
rect 44235 3499 44277 3508
rect 50859 3548 50901 3557
rect 50859 3508 50860 3548
rect 50900 3508 50901 3548
rect 50859 3499 50901 3508
rect 52683 3548 52725 3557
rect 52683 3508 52684 3548
rect 52724 3508 52725 3548
rect 52683 3499 52725 3508
rect 21187 3464 21245 3465
rect 21187 3424 21196 3464
rect 21236 3424 21245 3464
rect 21187 3423 21245 3424
rect 21483 3464 21525 3473
rect 21483 3424 21484 3464
rect 21524 3424 21525 3464
rect 21483 3415 21525 3424
rect 23683 3464 23741 3465
rect 23683 3424 23692 3464
rect 23732 3424 23741 3464
rect 23683 3423 23741 3424
rect 24547 3464 24605 3465
rect 24547 3424 24556 3464
rect 24596 3424 24605 3464
rect 27339 3451 27340 3491
rect 27380 3451 27381 3491
rect 27339 3442 27381 3451
rect 27619 3464 27677 3465
rect 24547 3423 24605 3424
rect 27619 3424 27628 3464
rect 27668 3424 27677 3464
rect 27619 3423 27677 3424
rect 31267 3464 31325 3465
rect 31267 3424 31276 3464
rect 31316 3424 31325 3464
rect 31267 3423 31325 3424
rect 32515 3464 32573 3465
rect 32515 3424 32524 3464
rect 32564 3424 32573 3464
rect 32515 3423 32573 3424
rect 33475 3464 33533 3465
rect 33475 3424 33484 3464
rect 33524 3424 33533 3464
rect 33475 3423 33533 3424
rect 33771 3464 33813 3473
rect 33771 3424 33772 3464
rect 33812 3424 33813 3464
rect 33771 3415 33813 3424
rect 35491 3464 35549 3465
rect 35491 3424 35500 3464
rect 35540 3424 35549 3464
rect 35491 3423 35549 3424
rect 35787 3464 35829 3473
rect 35787 3424 35788 3464
rect 35828 3424 35829 3464
rect 35787 3415 35829 3424
rect 39051 3464 39093 3473
rect 39051 3424 39052 3464
rect 39092 3424 39093 3464
rect 39051 3415 39093 3424
rect 39147 3464 39189 3473
rect 39147 3424 39148 3464
rect 39188 3424 39189 3464
rect 39147 3415 39189 3424
rect 39235 3464 39293 3465
rect 39235 3424 39244 3464
rect 39284 3424 39293 3464
rect 39235 3423 39293 3424
rect 39619 3464 39677 3465
rect 39619 3424 39628 3464
rect 39668 3424 39677 3464
rect 39619 3423 39677 3424
rect 39915 3464 39957 3473
rect 39915 3424 39916 3464
rect 39956 3424 39957 3464
rect 39915 3415 39957 3424
rect 40491 3464 40533 3473
rect 40491 3424 40492 3464
rect 40532 3424 40533 3464
rect 40491 3415 40533 3424
rect 40867 3464 40925 3465
rect 40867 3424 40876 3464
rect 40916 3424 40925 3464
rect 40867 3423 40925 3424
rect 41731 3464 41789 3465
rect 41731 3424 41740 3464
rect 41780 3424 41789 3464
rect 41731 3423 41789 3424
rect 43843 3464 43901 3465
rect 43843 3424 43852 3464
rect 43892 3424 43901 3464
rect 43843 3423 43901 3424
rect 44139 3464 44181 3473
rect 44139 3424 44140 3464
rect 44180 3424 44181 3464
rect 44139 3415 44181 3424
rect 45859 3464 45917 3465
rect 45859 3424 45868 3464
rect 45908 3424 45917 3464
rect 45859 3423 45917 3424
rect 46723 3464 46781 3465
rect 46723 3424 46732 3464
rect 46772 3424 46781 3464
rect 46723 3423 46781 3424
rect 47115 3464 47157 3473
rect 47115 3424 47116 3464
rect 47156 3424 47157 3464
rect 47115 3415 47157 3424
rect 47971 3464 48029 3465
rect 47971 3424 47980 3464
rect 48020 3424 48029 3464
rect 47971 3423 48029 3424
rect 48267 3464 48309 3473
rect 48267 3424 48268 3464
rect 48308 3424 48309 3464
rect 48267 3415 48309 3424
rect 48363 3464 48405 3473
rect 48363 3424 48364 3464
rect 48404 3424 48405 3464
rect 48363 3415 48405 3424
rect 49219 3464 49277 3465
rect 49219 3424 49228 3464
rect 49268 3424 49277 3464
rect 49219 3423 49277 3424
rect 49699 3464 49757 3465
rect 49699 3424 49708 3464
rect 49748 3424 49757 3464
rect 49699 3423 49757 3424
rect 50467 3464 50525 3465
rect 50467 3424 50476 3464
rect 50516 3424 50525 3464
rect 50467 3423 50525 3424
rect 50763 3464 50805 3473
rect 50763 3424 50764 3464
rect 50804 3424 50805 3464
rect 50763 3415 50805 3424
rect 53059 3464 53117 3465
rect 53059 3424 53068 3464
rect 53108 3424 53117 3464
rect 53059 3423 53117 3424
rect 53923 3464 53981 3465
rect 53923 3424 53932 3464
rect 53972 3424 53981 3464
rect 53923 3423 53981 3424
rect 21859 3296 21917 3297
rect 21859 3256 21868 3296
rect 21908 3256 21917 3296
rect 21859 3255 21917 3256
rect 26947 3296 27005 3297
rect 26947 3256 26956 3296
rect 26996 3256 27005 3296
rect 26947 3255 27005 3256
rect 40291 3296 40349 3297
rect 40291 3256 40300 3296
rect 40340 3256 40349 3296
rect 40291 3255 40349 3256
rect 44515 3296 44573 3297
rect 44515 3256 44524 3296
rect 44564 3256 44573 3296
rect 44515 3255 44573 3256
rect 48643 3296 48701 3297
rect 48643 3256 48652 3296
rect 48692 3256 48701 3296
rect 48643 3255 48701 3256
rect 51139 3296 51197 3297
rect 51139 3256 51148 3296
rect 51188 3256 51197 3296
rect 51139 3255 51197 3256
rect 34147 3212 34205 3213
rect 34147 3172 34156 3212
rect 34196 3172 34205 3212
rect 34147 3171 34205 3172
rect 36163 3212 36221 3213
rect 36163 3172 36172 3212
rect 36212 3172 36221 3212
rect 36163 3171 36221 3172
rect 576 3044 80736 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 80736 3044
rect 576 2980 80736 3004
rect 22723 2876 22781 2877
rect 22723 2836 22732 2876
rect 22772 2836 22781 2876
rect 22723 2835 22781 2836
rect 35971 2876 36029 2877
rect 35971 2836 35980 2876
rect 36020 2836 36029 2876
rect 35971 2835 36029 2836
rect 39043 2876 39101 2877
rect 39043 2836 39052 2876
rect 39092 2836 39101 2876
rect 39043 2835 39101 2836
rect 28675 2792 28733 2793
rect 28675 2752 28684 2792
rect 28724 2752 28733 2792
rect 28675 2751 28733 2752
rect 30019 2792 30077 2793
rect 30019 2752 30028 2792
rect 30068 2752 30077 2792
rect 30019 2751 30077 2752
rect 40483 2792 40541 2793
rect 40483 2752 40492 2792
rect 40532 2752 40541 2792
rect 40483 2751 40541 2752
rect 44227 2792 44285 2793
rect 44227 2752 44236 2792
rect 44276 2752 44285 2792
rect 44227 2751 44285 2752
rect 45187 2792 45245 2793
rect 45187 2752 45196 2792
rect 45236 2752 45245 2792
rect 45187 2751 45245 2752
rect 48451 2792 48509 2793
rect 48451 2752 48460 2792
rect 48500 2752 48509 2792
rect 48451 2751 48509 2752
rect 23499 2708 23541 2717
rect 23499 2668 23500 2708
rect 23540 2668 23541 2708
rect 23499 2659 23541 2668
rect 32227 2708 32285 2709
rect 32227 2668 32236 2708
rect 32276 2668 32285 2708
rect 32227 2667 32285 2668
rect 44899 2666 44957 2667
rect 20707 2624 20765 2625
rect 20707 2584 20716 2624
rect 20756 2584 20765 2624
rect 20707 2583 20765 2584
rect 21571 2624 21629 2625
rect 21571 2584 21580 2624
rect 21620 2584 21629 2624
rect 21571 2583 21629 2584
rect 24643 2624 24701 2625
rect 24643 2584 24652 2624
rect 24692 2584 24701 2624
rect 24643 2583 24701 2584
rect 25507 2624 25565 2625
rect 25507 2584 25516 2624
rect 25556 2584 25565 2624
rect 25507 2583 25565 2584
rect 28003 2624 28061 2625
rect 28003 2584 28012 2624
rect 28052 2584 28061 2624
rect 28003 2583 28061 2584
rect 28299 2624 28341 2633
rect 28299 2584 28300 2624
rect 28340 2584 28341 2624
rect 28299 2575 28341 2584
rect 30411 2624 30453 2633
rect 30411 2584 30412 2624
rect 30452 2584 30453 2624
rect 30411 2575 30453 2584
rect 30691 2624 30749 2625
rect 30691 2584 30700 2624
rect 30740 2584 30749 2624
rect 30691 2583 30749 2584
rect 33579 2624 33621 2633
rect 33579 2584 33580 2624
rect 33620 2584 33621 2624
rect 33579 2575 33621 2584
rect 33955 2624 34013 2625
rect 33955 2584 33964 2624
rect 34004 2584 34013 2624
rect 33955 2583 34013 2584
rect 34819 2624 34877 2625
rect 34819 2584 34828 2624
rect 34868 2584 34877 2624
rect 34819 2583 34877 2584
rect 36651 2624 36693 2633
rect 36651 2584 36652 2624
rect 36692 2584 36693 2624
rect 36651 2575 36693 2584
rect 37027 2624 37085 2625
rect 37027 2584 37036 2624
rect 37076 2584 37085 2624
rect 37027 2583 37085 2584
rect 37891 2624 37949 2625
rect 37891 2584 37900 2624
rect 37940 2584 37949 2624
rect 37891 2583 37949 2584
rect 39811 2624 39869 2625
rect 39811 2584 39820 2624
rect 39860 2584 39869 2624
rect 39811 2583 39869 2584
rect 40107 2624 40149 2633
rect 40107 2584 40108 2624
rect 40148 2584 40149 2624
rect 40107 2575 40149 2584
rect 40203 2624 40245 2633
rect 40203 2584 40204 2624
rect 40244 2584 40245 2624
rect 40203 2575 40245 2584
rect 43555 2624 43613 2625
rect 43555 2584 43564 2624
rect 43604 2584 43613 2624
rect 43555 2583 43613 2584
rect 43851 2624 43893 2633
rect 43851 2584 43852 2624
rect 43892 2584 43893 2624
rect 43851 2575 43893 2584
rect 44515 2624 44573 2625
rect 44515 2584 44524 2624
rect 44564 2584 44573 2624
rect 44515 2583 44573 2584
rect 44811 2624 44853 2633
rect 44899 2626 44908 2666
rect 44948 2626 44957 2666
rect 44899 2625 44957 2626
rect 44811 2584 44812 2624
rect 44852 2584 44853 2624
rect 44811 2575 44853 2584
rect 47779 2624 47837 2625
rect 47779 2584 47788 2624
rect 47828 2584 47837 2624
rect 47779 2583 47837 2584
rect 48075 2624 48117 2633
rect 48075 2584 48076 2624
rect 48116 2584 48117 2624
rect 48075 2575 48117 2584
rect 48171 2624 48213 2633
rect 48171 2584 48172 2624
rect 48212 2584 48213 2624
rect 48171 2575 48213 2584
rect 20331 2540 20373 2549
rect 20331 2500 20332 2540
rect 20372 2500 20373 2540
rect 20331 2491 20373 2500
rect 25899 2540 25941 2549
rect 25899 2500 25900 2540
rect 25940 2500 25941 2540
rect 25899 2491 25941 2500
rect 28395 2540 28437 2549
rect 28395 2500 28396 2540
rect 28436 2500 28437 2540
rect 28395 2491 28437 2500
rect 30315 2540 30357 2549
rect 30315 2500 30316 2540
rect 30356 2500 30357 2540
rect 30315 2491 30357 2500
rect 43947 2540 43989 2549
rect 43947 2500 43948 2540
rect 43988 2500 43989 2540
rect 43947 2491 43989 2500
rect 643 2456 701 2457
rect 643 2416 652 2456
rect 692 2416 701 2456
rect 643 2415 701 2416
rect 32427 2456 32469 2465
rect 32427 2416 32428 2456
rect 32468 2416 32469 2456
rect 32427 2407 32469 2416
rect 576 2288 80736 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80736 2288
rect 576 2224 80736 2248
rect 29251 2120 29309 2121
rect 29251 2080 29260 2120
rect 29300 2080 29309 2120
rect 29251 2079 29309 2080
rect 32035 2120 32093 2121
rect 32035 2080 32044 2120
rect 32084 2080 32093 2120
rect 32035 2079 32093 2080
rect 34627 2120 34685 2121
rect 34627 2080 34636 2120
rect 34676 2080 34685 2120
rect 34627 2079 34685 2080
rect 34915 2120 34973 2121
rect 34915 2080 34924 2120
rect 34964 2080 34973 2120
rect 34915 2079 34973 2080
rect 44227 2120 44285 2121
rect 44227 2080 44236 2120
rect 44276 2080 44285 2120
rect 44227 2079 44285 2080
rect 45091 2120 45149 2121
rect 45091 2080 45100 2120
rect 45140 2080 45149 2120
rect 45091 2079 45149 2080
rect 20619 2036 20661 2045
rect 20619 1996 20620 2036
rect 20660 1996 20661 2036
rect 20619 1987 20661 1996
rect 24267 2036 24309 2045
rect 24267 1996 24268 2036
rect 24308 1996 24309 2036
rect 24267 1987 24309 1996
rect 29643 2036 29685 2045
rect 29643 1996 29644 2036
rect 29684 1996 29685 2036
rect 29643 1987 29685 1996
rect 41355 2036 41397 2045
rect 41355 1996 41356 2036
rect 41396 1996 41397 2036
rect 41355 1987 41397 1996
rect 47499 2036 47541 2045
rect 47499 1996 47500 2036
rect 47540 1996 47541 2036
rect 47499 1987 47541 1996
rect 50859 2036 50901 2045
rect 50859 1996 50860 2036
rect 50900 1996 50901 2036
rect 50859 1987 50901 1996
rect 20715 1952 20757 1961
rect 20715 1912 20716 1952
rect 20756 1912 20757 1952
rect 20715 1903 20757 1912
rect 20995 1952 21053 1953
rect 20995 1912 21004 1952
rect 21044 1912 21053 1952
rect 20995 1911 21053 1912
rect 24363 1952 24405 1961
rect 24363 1912 24364 1952
rect 24404 1912 24405 1952
rect 24363 1903 24405 1912
rect 24643 1952 24701 1953
rect 24643 1912 24652 1952
rect 24692 1912 24701 1952
rect 24643 1911 24701 1912
rect 26859 1952 26901 1961
rect 26859 1912 26860 1952
rect 26900 1912 26901 1952
rect 26859 1903 26901 1912
rect 27235 1952 27293 1953
rect 27235 1912 27244 1952
rect 27284 1912 27293 1952
rect 27235 1911 27293 1912
rect 28099 1952 28157 1953
rect 28099 1912 28108 1952
rect 28148 1912 28157 1952
rect 28099 1911 28157 1912
rect 30019 1952 30077 1953
rect 30019 1912 30028 1952
rect 30068 1912 30077 1952
rect 30019 1911 30077 1912
rect 30883 1952 30941 1953
rect 30883 1912 30892 1952
rect 30932 1912 30941 1952
rect 30883 1911 30941 1912
rect 32235 1952 32277 1961
rect 36931 1957 36989 1958
rect 32235 1912 32236 1952
rect 32276 1912 32277 1952
rect 32235 1903 32277 1912
rect 32611 1952 32669 1953
rect 32611 1912 32620 1952
rect 32660 1912 32669 1952
rect 32611 1911 32669 1912
rect 33475 1952 33533 1953
rect 33475 1912 33484 1952
rect 33524 1912 33533 1952
rect 33475 1911 33533 1912
rect 36067 1952 36125 1953
rect 36067 1912 36076 1952
rect 36116 1912 36125 1952
rect 36931 1917 36940 1957
rect 36980 1917 36989 1957
rect 36931 1916 36989 1917
rect 37323 1952 37365 1961
rect 36067 1911 36125 1912
rect 37323 1912 37324 1952
rect 37364 1912 37365 1952
rect 37323 1903 37365 1912
rect 38851 1952 38909 1953
rect 38851 1912 38860 1952
rect 38900 1912 38909 1952
rect 38851 1911 38909 1912
rect 39715 1952 39773 1953
rect 39715 1912 39724 1952
rect 39764 1912 39773 1952
rect 39715 1911 39773 1912
rect 40107 1952 40149 1961
rect 40107 1912 40108 1952
rect 40148 1912 40149 1952
rect 40107 1903 40149 1912
rect 40963 1952 41021 1953
rect 40963 1912 40972 1952
rect 41012 1912 41021 1952
rect 40963 1911 41021 1912
rect 41259 1952 41301 1961
rect 41259 1912 41260 1952
rect 41300 1912 41301 1952
rect 41259 1903 41301 1912
rect 41835 1952 41877 1961
rect 41835 1912 41836 1952
rect 41876 1912 41877 1952
rect 41835 1903 41877 1912
rect 42211 1952 42269 1953
rect 42211 1912 42220 1952
rect 42260 1912 42269 1952
rect 42211 1911 42269 1912
rect 43075 1952 43133 1953
rect 43075 1912 43084 1952
rect 43124 1912 43133 1952
rect 43075 1911 43133 1912
rect 46243 1952 46301 1953
rect 46243 1912 46252 1952
rect 46292 1912 46301 1952
rect 46243 1911 46301 1912
rect 47107 1952 47165 1953
rect 47107 1912 47116 1952
rect 47156 1912 47165 1952
rect 47107 1911 47165 1912
rect 49603 1952 49661 1953
rect 49603 1912 49612 1952
rect 49652 1912 49661 1952
rect 49603 1911 49661 1912
rect 50467 1952 50525 1953
rect 50467 1912 50476 1952
rect 50516 1912 50525 1952
rect 50467 1911 50525 1912
rect 48459 1868 48501 1877
rect 48459 1828 48460 1868
rect 48500 1828 48501 1868
rect 48459 1819 48501 1828
rect 20323 1784 20381 1785
rect 20323 1744 20332 1784
rect 20372 1744 20381 1784
rect 20323 1743 20381 1744
rect 23971 1784 24029 1785
rect 23971 1744 23980 1784
rect 24020 1744 24029 1784
rect 23971 1743 24029 1744
rect 41635 1784 41693 1785
rect 41635 1744 41644 1784
rect 41684 1744 41693 1784
rect 41635 1743 41693 1744
rect 34627 1700 34685 1701
rect 34627 1660 34636 1700
rect 34676 1660 34685 1700
rect 34627 1659 34685 1660
rect 37699 1700 37757 1701
rect 37699 1660 37708 1700
rect 37748 1660 37757 1700
rect 37699 1659 37757 1660
rect 576 1532 80736 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 80736 1532
rect 576 1468 80736 1492
rect 26659 1364 26717 1365
rect 26659 1324 26668 1364
rect 26708 1324 26717 1364
rect 26659 1323 26717 1324
rect 30787 1364 30845 1365
rect 30787 1324 30796 1364
rect 30836 1324 30845 1364
rect 30787 1323 30845 1324
rect 32035 1364 32093 1365
rect 32035 1324 32044 1364
rect 32084 1324 32093 1364
rect 32035 1323 32093 1324
rect 35587 1364 35645 1365
rect 35587 1324 35596 1364
rect 35636 1324 35645 1364
rect 35587 1323 35645 1324
rect 38851 1364 38909 1365
rect 38851 1324 38860 1364
rect 38900 1324 38909 1364
rect 38851 1323 38909 1324
rect 40195 1364 40253 1365
rect 40195 1324 40204 1364
rect 40244 1324 40253 1364
rect 40195 1323 40253 1324
rect 44131 1364 44189 1365
rect 44131 1324 44140 1364
rect 44180 1324 44189 1364
rect 44131 1323 44189 1324
rect 47779 1364 47837 1365
rect 47779 1324 47788 1364
rect 47828 1324 47837 1364
rect 47779 1323 47837 1324
rect 47587 1280 47645 1281
rect 47587 1240 47596 1280
rect 47636 1240 47645 1280
rect 47587 1239 47645 1240
rect 27331 1129 27389 1130
rect 26955 1112 26997 1121
rect 26955 1072 26956 1112
rect 26996 1072 26997 1112
rect 26955 1063 26997 1072
rect 27051 1112 27093 1121
rect 27051 1072 27052 1112
rect 27092 1072 27093 1112
rect 27331 1089 27340 1129
rect 27380 1089 27389 1129
rect 27331 1088 27389 1089
rect 28395 1112 28437 1121
rect 27051 1063 27093 1072
rect 28395 1072 28396 1112
rect 28436 1072 28437 1112
rect 28395 1063 28437 1072
rect 28771 1112 28829 1113
rect 28771 1072 28780 1112
rect 28820 1072 28829 1112
rect 28771 1071 28829 1072
rect 29635 1112 29693 1113
rect 29635 1072 29644 1112
rect 29684 1072 29693 1112
rect 29635 1071 29693 1072
rect 32331 1112 32373 1121
rect 32331 1072 32332 1112
rect 32372 1072 32373 1112
rect 32331 1063 32373 1072
rect 32427 1112 32469 1121
rect 32427 1072 32428 1112
rect 32468 1072 32469 1112
rect 34915 1112 34973 1113
rect 32427 1063 32469 1072
rect 32725 1097 32783 1098
rect 32725 1057 32734 1097
rect 32774 1057 32783 1097
rect 34915 1072 34924 1112
rect 34964 1072 34973 1112
rect 34915 1071 34973 1072
rect 35211 1112 35253 1121
rect 35211 1072 35212 1112
rect 35252 1072 35253 1112
rect 35211 1063 35253 1072
rect 35307 1112 35349 1121
rect 35307 1072 35308 1112
rect 35348 1072 35349 1112
rect 35307 1063 35349 1072
rect 38179 1112 38237 1113
rect 38179 1072 38188 1112
rect 38228 1072 38237 1112
rect 38179 1071 38237 1072
rect 38475 1112 38517 1121
rect 38475 1072 38476 1112
rect 38516 1072 38517 1112
rect 38475 1063 38517 1072
rect 38571 1112 38613 1121
rect 38571 1072 38572 1112
rect 38612 1072 38613 1112
rect 38571 1063 38613 1072
rect 41347 1112 41405 1113
rect 41347 1072 41356 1112
rect 41396 1072 41405 1112
rect 41347 1071 41405 1072
rect 42211 1112 42269 1113
rect 42211 1072 42220 1112
rect 42260 1072 42269 1112
rect 42211 1071 42269 1072
rect 42603 1112 42645 1121
rect 42603 1072 42604 1112
rect 42644 1072 42645 1112
rect 42603 1063 42645 1072
rect 45283 1112 45341 1113
rect 45283 1072 45292 1112
rect 45332 1072 45341 1112
rect 45283 1071 45341 1072
rect 46147 1112 46205 1113
rect 46147 1072 46156 1112
rect 46196 1072 46205 1112
rect 46147 1071 46205 1072
rect 46539 1112 46581 1121
rect 46539 1072 46540 1112
rect 46580 1072 46581 1112
rect 46539 1063 46581 1072
rect 46915 1112 46973 1113
rect 46915 1072 46924 1112
rect 46964 1072 46973 1112
rect 46915 1071 46973 1072
rect 47211 1112 47253 1121
rect 47211 1072 47212 1112
rect 47252 1072 47253 1112
rect 47211 1063 47253 1072
rect 47307 1112 47349 1121
rect 47307 1072 47308 1112
rect 47348 1072 47349 1112
rect 47307 1063 47349 1072
rect 48931 1112 48989 1113
rect 48931 1072 48940 1112
rect 48980 1072 48989 1112
rect 48931 1071 48989 1072
rect 49795 1112 49853 1113
rect 49795 1072 49804 1112
rect 49844 1072 49853 1112
rect 49795 1071 49853 1072
rect 50187 1112 50229 1121
rect 50187 1072 50188 1112
rect 50228 1072 50229 1112
rect 50187 1063 50229 1072
rect 32725 1056 32783 1057
rect 576 776 80736 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80736 776
rect 576 712 80736 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 22060 38368 22100 38408
rect 26572 38368 26612 38408
rect 27532 38368 27572 38408
rect 27628 38284 27668 38324
rect 29452 38284 29492 38324
rect 33676 38284 33716 38324
rect 21964 38200 22004 38240
rect 25996 38200 26036 38240
rect 26476 38200 26516 38240
rect 26668 38200 26708 38240
rect 27724 38200 27764 38240
rect 27820 38200 27860 38240
rect 28972 38200 29012 38240
rect 29260 38200 29300 38240
rect 29740 38200 29780 38240
rect 29932 38200 29972 38240
rect 33292 38200 33332 38240
rect 33580 38200 33620 38240
rect 37516 38200 37556 38240
rect 37420 38158 37460 38198
rect 37804 38200 37844 38240
rect 652 38116 692 38156
rect 22732 38116 22772 38156
rect 23692 38116 23732 38156
rect 24268 38116 24308 38156
rect 24652 38116 24692 38156
rect 24460 38032 24500 38072
rect 844 37948 884 37988
rect 21772 37948 21812 37988
rect 22540 37948 22580 37988
rect 23884 37948 23924 37988
rect 24076 37948 24116 37988
rect 26092 37948 26132 37988
rect 27532 37948 27572 37988
rect 29836 37948 29876 37988
rect 33964 37948 34004 37988
rect 37132 37948 37172 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 26668 37612 26708 37652
rect 19756 37444 19796 37484
rect 32908 37444 32948 37484
rect 20620 37360 20660 37400
rect 20716 37360 20756 37400
rect 21004 37360 21044 37400
rect 21388 37360 21428 37400
rect 22252 37360 22292 37400
rect 23980 37360 24020 37400
rect 24844 37360 24884 37400
rect 26380 37360 26420 37400
rect 26476 37360 26516 37400
rect 26668 37360 26708 37400
rect 26860 37360 26900 37400
rect 27244 37360 27284 37400
rect 28108 37360 28148 37400
rect 29740 37360 29780 37400
rect 29836 37360 29876 37400
rect 30604 37360 30644 37400
rect 31468 37360 31508 37400
rect 34444 37360 34484 37400
rect 35308 37360 35348 37400
rect 35692 37360 35732 37400
rect 36652 37360 36692 37400
rect 36940 37360 36980 37400
rect 37324 37360 37364 37400
rect 37708 37360 37748 37400
rect 38572 37360 38612 37400
rect 41068 37360 41108 37400
rect 41932 37360 41972 37400
rect 23596 37276 23636 37316
rect 30220 37276 30260 37316
rect 36556 37276 36596 37316
rect 42316 37276 42356 37316
rect 19564 37192 19604 37232
rect 20428 37192 20468 37232
rect 23404 37192 23444 37232
rect 25996 37192 26036 37232
rect 29260 37192 29300 37232
rect 30028 37192 30068 37232
rect 32620 37192 32660 37232
rect 33100 37192 33140 37232
rect 33292 37192 33332 37232
rect 39724 37192 39764 37232
rect 39916 37192 39956 37232
rect 36268 37150 36308 37190
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 22540 36914 22580 36954
rect 21100 36856 21140 36896
rect 23404 36856 23444 36896
rect 24844 36856 24884 36896
rect 25132 36856 25172 36896
rect 25612 36856 25652 36896
rect 28108 36856 28148 36896
rect 32044 36856 32084 36896
rect 38476 36856 38516 36896
rect 25324 36772 25364 36812
rect 26284 36772 26324 36812
rect 29644 36772 29684 36812
rect 32716 36772 32756 36812
rect 36076 36772 36116 36812
rect 40012 36772 40052 36812
rect 18700 36688 18740 36728
rect 19084 36688 19124 36728
rect 19948 36688 19988 36728
rect 21388 36688 21428 36728
rect 22348 36688 22388 36728
rect 22444 36688 22484 36728
rect 23020 36688 23060 36728
rect 23116 36688 23156 36728
rect 23884 36688 23924 36728
rect 23980 36688 24020 36728
rect 24172 36688 24212 36728
rect 24364 36688 24404 36728
rect 24460 36688 24500 36728
rect 24652 36688 24692 36728
rect 24940 36688 24980 36728
rect 25516 36688 25556 36728
rect 25612 36688 25652 36728
rect 26380 36688 26420 36728
rect 26764 36688 26804 36728
rect 27148 36688 27188 36728
rect 27244 36688 27284 36728
rect 27340 36688 27380 36728
rect 27436 36688 27476 36728
rect 28012 36688 28052 36728
rect 30028 36688 30068 36728
rect 30892 36688 30932 36728
rect 33100 36701 33140 36741
rect 33964 36688 34004 36728
rect 35308 36688 35348 36728
rect 35500 36688 35540 36728
rect 35692 36688 35732 36728
rect 35884 36688 35924 36728
rect 36460 36688 36500 36728
rect 37324 36688 37364 36728
rect 39628 36688 39668 36728
rect 39916 36688 39956 36728
rect 41548 36688 41588 36728
rect 41932 36688 41972 36728
rect 42796 36688 42836 36728
rect 32524 36604 32564 36644
rect 35788 36604 35828 36644
rect 22060 36520 22100 36560
rect 24172 36520 24212 36560
rect 27628 36520 27668 36560
rect 27820 36520 27860 36560
rect 40300 36520 40340 36560
rect 21292 36436 21332 36476
rect 24652 36436 24692 36476
rect 32332 36436 32372 36476
rect 35116 36436 35156 36476
rect 35308 36436 35348 36476
rect 43948 36436 43988 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 20524 36100 20564 36140
rect 21964 36100 22004 36140
rect 25708 36100 25748 36140
rect 32236 36100 32276 36140
rect 41644 36100 41684 36140
rect 16876 36016 16916 36056
rect 19180 36016 19220 36056
rect 20332 36016 20372 36056
rect 22924 36016 22964 36056
rect 27820 36016 27860 36056
rect 35116 36016 35156 36056
rect 36460 36016 36500 36056
rect 40588 36016 40628 36056
rect 43756 36016 43796 36056
rect 46252 36016 46292 36056
rect 49612 36016 49652 36056
rect 51340 36016 51380 36056
rect 52300 36016 52340 36056
rect 13900 35932 13940 35972
rect 35308 35932 35348 35972
rect 43948 35932 43988 35972
rect 44524 35932 44564 35972
rect 16204 35848 16244 35888
rect 16492 35848 16532 35888
rect 18508 35848 18548 35888
rect 18796 35848 18836 35888
rect 19660 35848 19700 35888
rect 19948 35848 19988 35888
rect 20812 35848 20852 35888
rect 20908 35848 20948 35888
rect 21196 35848 21236 35888
rect 21484 35848 21524 35888
rect 21676 35848 21716 35888
rect 21772 35848 21812 35888
rect 21964 35848 22004 35888
rect 22252 35848 22292 35888
rect 22540 35848 22580 35888
rect 23308 35848 23348 35888
rect 23692 35848 23732 35888
rect 24556 35848 24596 35888
rect 27100 35848 27140 35888
rect 27532 35848 27572 35888
rect 27724 35848 27764 35888
rect 27820 35848 27860 35888
rect 31564 35848 31604 35888
rect 31852 35848 31892 35888
rect 31948 35848 31988 35888
rect 32524 35848 32564 35888
rect 34828 35848 34868 35888
rect 34924 35848 34964 35888
rect 35116 35859 35156 35899
rect 35404 35848 35444 35888
rect 35596 35848 35636 35888
rect 35788 35848 35828 35888
rect 35980 35848 36020 35888
rect 36172 35848 36212 35888
rect 36268 35848 36308 35888
rect 36748 35848 36788 35888
rect 36844 35848 36884 35888
rect 37132 35848 37172 35888
rect 39916 35848 39956 35888
rect 40204 35848 40244 35888
rect 40300 35848 40340 35888
rect 40972 35848 41012 35888
rect 41260 35848 41300 35888
rect 41356 35848 41396 35888
rect 43084 35848 43124 35888
rect 43372 35848 43412 35888
rect 45580 35848 45620 35888
rect 45868 35848 45908 35888
rect 48940 35848 48980 35888
rect 49228 35848 49268 35888
rect 50668 35848 50708 35888
rect 50956 35848 50996 35888
rect 51628 35848 51668 35888
rect 51916 35848 51956 35888
rect 16588 35764 16628 35804
rect 18892 35764 18932 35804
rect 20044 35764 20084 35804
rect 22636 35764 22676 35804
rect 26188 35764 26228 35804
rect 43468 35764 43508 35804
rect 45964 35764 46004 35804
rect 49324 35764 49364 35804
rect 51052 35764 51092 35804
rect 52012 35764 52052 35804
rect 14092 35680 14132 35720
rect 21004 35676 21044 35716
rect 21388 35680 21428 35720
rect 34348 35680 34388 35720
rect 35692 35680 35732 35720
rect 36076 35680 36116 35720
rect 44140 35680 44180 35720
rect 44716 35680 44756 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 17548 35344 17588 35384
rect 28492 35344 28532 35384
rect 33388 35344 33428 35384
rect 38380 35344 38420 35384
rect 43276 35344 43316 35384
rect 44332 35344 44372 35384
rect 51916 35344 51956 35384
rect 19948 35260 19988 35300
rect 20716 35260 20756 35300
rect 26092 35260 26132 35300
rect 35788 35260 35828 35300
rect 35980 35260 36020 35300
rect 46732 35260 46772 35300
rect 49516 35260 49556 35300
rect 52108 35260 52148 35300
rect 13228 35176 13268 35216
rect 13324 35176 13364 35216
rect 13612 35176 13652 35216
rect 14092 35176 14132 35216
rect 14380 35176 14420 35216
rect 14476 35176 14516 35216
rect 14956 35176 14996 35216
rect 15340 35176 15380 35216
rect 16204 35176 16244 35216
rect 18700 35176 18740 35216
rect 19564 35176 19604 35216
rect 21100 35176 21140 35216
rect 21964 35176 22004 35216
rect 25036 35176 25076 35216
rect 26476 35176 26516 35216
rect 27340 35176 27380 35216
rect 30028 35176 30068 35216
rect 30412 35176 30452 35216
rect 31276 35176 31316 35216
rect 34540 35176 34580 35216
rect 35404 35176 35444 35216
rect 36364 35176 36404 35216
rect 37228 35176 37268 35216
rect 40012 35176 40052 35216
rect 40300 35176 40340 35216
rect 40396 35176 40436 35216
rect 40876 35176 40916 35216
rect 41260 35176 41300 35216
rect 42124 35176 42164 35216
rect 45484 35176 45524 35216
rect 46348 35176 46388 35216
rect 46924 35176 46964 35216
rect 47308 35176 47348 35216
rect 48172 35176 48212 35216
rect 49900 35176 49940 35216
rect 50764 35176 50804 35216
rect 52492 35176 52532 35216
rect 53356 35176 53396 35216
rect 64588 35176 64628 35216
rect 70156 35176 70196 35216
rect 10636 35092 10676 35132
rect 20332 35092 20372 35132
rect 43660 35092 43700 35132
rect 43948 35092 43988 35132
rect 14764 35008 14804 35048
rect 20140 35008 20180 35048
rect 40684 35008 40724 35048
rect 64396 35008 64436 35048
rect 10444 34924 10484 34964
rect 12940 34924 12980 34964
rect 17356 34924 17396 34964
rect 17548 34924 17588 34964
rect 23116 34924 23156 34964
rect 25228 34924 25268 34964
rect 32428 34924 32468 34964
rect 43468 34924 43508 34964
rect 44140 34924 44180 34964
rect 49324 34924 49364 34964
rect 51916 34924 51956 34964
rect 54508 34924 54548 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 19276 34588 19316 34628
rect 30220 34588 30260 34628
rect 46540 34588 46580 34628
rect 47980 34588 48020 34628
rect 7564 34504 7604 34544
rect 10636 34504 10676 34544
rect 26476 34504 26516 34544
rect 27436 34504 27476 34544
rect 31948 34504 31988 34544
rect 36940 34504 36980 34544
rect 70924 34504 70964 34544
rect 25516 34420 25556 34460
rect 26284 34420 26324 34460
rect 7852 34336 7892 34376
rect 9964 34336 10004 34376
rect 10252 34336 10292 34376
rect 10828 34336 10868 34376
rect 11212 34336 11252 34376
rect 12076 34336 12116 34376
rect 13420 34336 13460 34376
rect 13804 34336 13844 34376
rect 14668 34336 14708 34376
rect 16876 34336 16916 34376
rect 17308 34336 17348 34376
rect 18124 34336 18164 34376
rect 19564 34336 19604 34376
rect 20524 34336 20564 34376
rect 21004 34336 21044 34376
rect 21292 34336 21332 34376
rect 22252 34336 22292 34376
rect 23116 34336 23156 34376
rect 23500 34336 23540 34376
rect 24364 34336 24404 34376
rect 26764 34336 26804 34376
rect 27052 34336 27092 34376
rect 27628 34336 27668 34376
rect 28012 34336 28052 34376
rect 28876 34336 28916 34376
rect 30508 34336 30548 34376
rect 30604 34336 30644 34376
rect 30892 34336 30932 34376
rect 31276 34336 31316 34376
rect 31564 34336 31604 34376
rect 32140 34336 32180 34376
rect 32524 34336 32564 34376
rect 33388 34336 33428 34376
rect 35692 34336 35732 34376
rect 36268 34336 36308 34376
rect 36556 34336 36596 34376
rect 38092 34336 38132 34376
rect 39148 34336 39188 34376
rect 40012 34336 40052 34376
rect 42220 34336 42260 34376
rect 43660 34336 43700 34376
rect 43948 34336 43988 34376
rect 44332 34336 44372 34376
rect 45196 34336 45236 34376
rect 46828 34336 46868 34376
rect 46924 34336 46964 34376
rect 47212 34336 47252 34376
rect 49612 34336 49652 34376
rect 50860 34336 50900 34376
rect 52492 34336 52532 34376
rect 53164 34336 53204 34376
rect 54028 34336 54068 34376
rect 61516 34336 61556 34376
rect 62476 34336 62516 34376
rect 62764 34336 62804 34376
rect 64204 34336 64244 34376
rect 65452 34336 65492 34376
rect 66316 34336 66356 34376
rect 68044 34336 68084 34376
rect 68908 34336 68948 34376
rect 69292 34336 69332 34376
rect 70156 34336 70196 34376
rect 70636 34336 70676 34376
rect 10348 34252 10388 34292
rect 27148 34252 27188 34292
rect 31660 34252 31700 34292
rect 36652 34252 36692 34292
rect 38764 34252 38804 34292
rect 52780 34252 52820 34292
rect 7372 34168 7412 34208
rect 13228 34168 13268 34208
rect 15820 34168 15860 34208
rect 19276 34168 19316 34208
rect 30028 34168 30068 34208
rect 34540 34168 34580 34208
rect 35212 34168 35252 34208
rect 37612 34168 37652 34208
rect 41164 34168 41204 34208
rect 46348 34168 46388 34208
rect 50380 34168 50420 34208
rect 52012 34168 52052 34208
rect 55180 34168 55220 34208
rect 64588 34168 64628 34208
rect 68524 34168 68564 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 80812 33664 80852 33704
rect 81196 33664 81236 33704
rect 82060 33664 82100 33704
rect 83212 33412 83252 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 80524 33076 80564 33116
rect 5548 32908 5588 32948
rect 80140 32908 80180 32948
rect 82060 32908 82100 32948
rect 80812 32824 80852 32864
rect 80908 32824 80948 32864
rect 81196 32824 81236 32864
rect 5356 32656 5396 32696
rect 80332 32656 80372 32696
rect 81868 32656 81908 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 4588 32320 4628 32360
rect 5740 32152 5780 32192
rect 80812 32152 80852 32192
rect 81196 32152 81236 32192
rect 82060 32152 82100 32192
rect 4396 32068 4436 32108
rect 4588 31900 4628 31940
rect 5068 31900 5108 31940
rect 83212 31900 83252 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 5836 31564 5876 31604
rect 80716 31564 80756 31604
rect 80332 31396 80372 31436
rect 3820 31312 3860 31352
rect 4684 31312 4724 31352
rect 81100 31312 81140 31352
rect 81388 31312 81428 31352
rect 3436 31228 3476 31268
rect 81004 31228 81044 31268
rect 5836 31144 5876 31184
rect 80140 31144 80180 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 82924 30808 82964 30848
rect 4492 30724 4532 30764
rect 80044 30724 80084 30764
rect 4588 30640 4628 30680
rect 4876 30640 4916 30680
rect 79660 30640 79700 30680
rect 79948 30640 79988 30680
rect 80524 30640 80564 30680
rect 80908 30640 80948 30680
rect 81772 30640 81812 30680
rect 79180 30556 79220 30596
rect 4204 30472 4244 30512
rect 80332 30472 80372 30512
rect 79372 30388 79412 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 81388 29968 81428 30008
rect 79180 29800 79220 29840
rect 80044 29800 80084 29840
rect 81676 29800 81716 29840
rect 81772 29800 81812 29840
rect 82060 29800 82100 29840
rect 78796 29716 78836 29756
rect 81196 29632 81236 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 83212 29296 83252 29336
rect 79660 29212 79700 29252
rect 80812 29212 80852 29252
rect 4588 29128 4628 29168
rect 5452 29128 5492 29168
rect 5836 29128 5876 29168
rect 79756 29128 79796 29168
rect 80044 29128 80084 29168
rect 81196 29128 81236 29168
rect 82060 29128 82100 29168
rect 79372 28960 79412 29000
rect 3436 28876 3476 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 5164 28540 5204 28580
rect 83212 28540 83252 28580
rect 80620 28456 80660 28496
rect 4492 28288 4532 28328
rect 4780 28288 4820 28328
rect 74188 28288 74228 28328
rect 79948 28288 79988 28328
rect 80236 28288 80276 28328
rect 80332 28288 80372 28328
rect 80812 28288 80852 28328
rect 81196 28288 81236 28328
rect 82060 28288 82100 28328
rect 4876 28204 4916 28244
rect 75820 28120 75860 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 80524 27700 80564 27740
rect 80140 27616 80180 27656
rect 80428 27616 80468 27656
rect 80812 27364 80852 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 83212 27028 83252 27068
rect 79852 26944 79892 26984
rect 80236 26776 80276 26816
rect 80524 26776 80564 26816
rect 80812 26776 80852 26816
rect 81196 26776 81236 26816
rect 82060 26776 82100 26816
rect 80140 26692 80180 26732
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 5836 26272 5876 26312
rect 80236 26188 80276 26228
rect 3436 26104 3476 26144
rect 3820 26104 3860 26144
rect 4684 26104 4724 26144
rect 80620 26104 80660 26144
rect 81484 26104 81524 26144
rect 82636 25936 82676 25976
rect 5836 25852 5876 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 4204 25516 4244 25556
rect 80236 25432 80276 25472
rect 81196 25432 81236 25472
rect 652 25348 692 25388
rect 4492 25264 4532 25304
rect 4588 25264 4628 25304
rect 4876 25264 4916 25304
rect 80620 25264 80660 25304
rect 80908 25264 80948 25304
rect 81484 25264 81524 25304
rect 81580 25264 81620 25304
rect 81868 25264 81908 25304
rect 80524 25180 80564 25220
rect 844 25096 884 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 844 24760 884 24800
rect 80236 24676 80276 24716
rect 80620 24592 80660 24632
rect 81484 24592 81524 24632
rect 652 24508 692 24548
rect 82636 24508 82676 24548
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 844 24004 884 24044
rect 5836 24004 5876 24044
rect 83212 24004 83252 24044
rect 652 23836 692 23876
rect 3820 23752 3860 23792
rect 4684 23752 4724 23792
rect 80812 23752 80852 23792
rect 81196 23752 81236 23792
rect 82060 23752 82100 23792
rect 3436 23668 3476 23708
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 844 23248 884 23288
rect 4204 23290 4244 23330
rect 4492 23164 4532 23204
rect 3532 23080 3572 23120
rect 3628 23080 3668 23120
rect 3916 23080 3956 23120
rect 4588 23080 4628 23120
rect 4876 23080 4916 23120
rect 652 22996 692 23036
rect 3244 22828 3284 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 5836 22492 5876 22532
rect 3436 22240 3476 22280
rect 3820 22240 3860 22280
rect 4684 22240 4724 22280
rect 652 22072 692 22112
rect 5836 22072 5876 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3340 21652 3380 21692
rect 3436 21568 3476 21608
rect 3724 21568 3764 21608
rect 3052 21316 3092 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 5356 20980 5396 21020
rect 84460 20980 84500 21020
rect 81772 20896 81812 20936
rect 2956 20728 2996 20768
rect 3340 20728 3380 20768
rect 4204 20728 4244 20768
rect 81100 20728 81140 20768
rect 81388 20728 81428 20768
rect 81484 20728 81524 20768
rect 82444 20728 82484 20768
rect 83308 20728 83348 20768
rect 82060 20644 82100 20684
rect 652 20560 692 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 652 20224 692 20264
rect 3436 20056 3476 20096
rect 3820 20056 3860 20096
rect 4684 20056 4724 20096
rect 96748 20056 96788 20096
rect 5836 19972 5876 20012
rect 98572 19888 98612 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 3628 19468 3668 19508
rect 2860 19300 2900 19340
rect 3436 19300 3476 19340
rect 3916 19216 3956 19256
rect 4012 19216 4052 19256
rect 4300 19216 4340 19256
rect 652 19048 692 19088
rect 3052 19048 3092 19088
rect 3244 19048 3284 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 652 18712 692 18752
rect 2956 18628 2996 18668
rect 2572 18544 2612 18584
rect 2860 18544 2900 18584
rect 3436 18544 3476 18584
rect 3820 18544 3860 18584
rect 4684 18544 4724 18584
rect 2284 18460 2324 18500
rect 5836 18460 5876 18500
rect 3244 18376 3284 18416
rect 2092 18292 2132 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 5068 17872 5108 17912
rect 2476 17788 2516 17828
rect 3052 17704 3092 17744
rect 3916 17704 3956 17744
rect 2668 17620 2708 17660
rect 652 17536 692 17576
rect 2284 17536 2324 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 652 17200 692 17240
rect 2668 17116 2708 17156
rect 2284 17032 2324 17072
rect 2572 17032 2612 17072
rect 78220 17032 78260 17072
rect 78604 17032 78644 17072
rect 79468 17032 79508 17072
rect 3244 16948 3284 16988
rect 2956 16864 2996 16904
rect 3436 16780 3476 16820
rect 80620 16780 80660 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 3244 16444 3284 16484
rect 5836 16444 5876 16484
rect 78124 16444 78164 16484
rect 1228 16192 1268 16232
rect 2092 16192 2132 16232
rect 3820 16192 3860 16232
rect 4684 16192 4724 16232
rect 78412 16192 78452 16232
rect 78508 16192 78548 16232
rect 78796 16192 78836 16232
rect 844 16108 884 16148
rect 3436 16108 3476 16148
rect 5836 16024 5876 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 652 15688 692 15728
rect 1804 15604 1844 15644
rect 4492 15604 4532 15644
rect 1900 15520 1940 15560
rect 2188 15520 2228 15560
rect 4588 15520 4628 15560
rect 4876 15520 4916 15560
rect 1228 15436 1268 15476
rect 1516 15352 1556 15392
rect 4204 15352 4244 15392
rect 1036 15268 1076 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 5836 14932 5876 14972
rect 3244 14848 3284 14888
rect 1228 14680 1268 14720
rect 2092 14680 2132 14720
rect 3820 14680 3860 14720
rect 4684 14680 4724 14720
rect 844 14596 884 14636
rect 3436 14596 3476 14636
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 1612 14092 1652 14132
rect 3820 14092 3860 14132
rect 1708 14008 1748 14048
rect 1996 14008 2036 14048
rect 3916 14008 3956 14048
rect 4204 14008 4244 14048
rect 844 13924 884 13964
rect 652 13840 692 13880
rect 1324 13840 1364 13880
rect 3532 13840 3572 13880
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 1228 13168 1268 13208
rect 2092 13168 2132 13208
rect 3820 13168 3860 13208
rect 4684 13168 4724 13208
rect 844 13084 884 13124
rect 3436 13084 3476 13124
rect 3244 13000 3284 13040
rect 5836 13000 5876 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 652 12664 692 12704
rect 3820 12580 3860 12620
rect 1708 12496 1748 12536
rect 1804 12496 1844 12536
rect 2092 12496 2132 12536
rect 3916 12496 3956 12536
rect 4204 12496 4244 12536
rect 844 12412 884 12452
rect 1228 12412 1268 12452
rect 1036 12328 1076 12368
rect 1420 12328 1460 12368
rect 3532 12328 3572 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 5836 11908 5876 11948
rect 3244 11824 3284 11864
rect 844 11740 884 11780
rect 2860 11698 2900 11738
rect 2572 11656 2612 11696
rect 2956 11656 2996 11696
rect 3436 11656 3476 11696
rect 3820 11656 3860 11696
rect 4684 11656 4724 11696
rect 652 11488 692 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 4876 11152 4916 11192
rect 2476 10984 2516 11024
rect 2908 10984 2948 11024
rect 3724 10984 3764 11024
rect 844 10900 884 10940
rect 652 10732 692 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 2284 10396 2324 10436
rect 3916 10312 3956 10352
rect 844 10228 884 10268
rect 2572 10144 2612 10184
rect 2668 10144 2708 10184
rect 2956 10144 2996 10184
rect 4300 10144 4340 10184
rect 4588 10144 4628 10184
rect 4204 10060 4244 10100
rect 652 9976 692 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 5836 9640 5876 9680
rect 3436 9556 3476 9596
rect 3820 9472 3860 9512
rect 4684 9472 4724 9512
rect 844 9388 884 9428
rect 652 9220 692 9260
rect 5836 9220 5876 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 652 8464 692 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 652 8128 692 8168
rect 5836 8128 5876 8168
rect 3436 7960 3476 8000
rect 3820 7960 3860 8000
rect 4684 7960 4724 8000
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 4300 7372 4340 7412
rect 4588 7120 4628 7160
rect 4684 7120 4724 7160
rect 4972 7120 5012 7160
rect 652 6952 692 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 80524 6616 80564 6656
rect 78508 6448 78548 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 652 5440 692 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 652 5104 692 5144
rect 21580 5104 21620 5144
rect 25708 5104 25748 5144
rect 35884 5104 35924 5144
rect 39436 5104 39476 5144
rect 44524 5104 44564 5144
rect 49996 5104 50036 5144
rect 17548 5020 17588 5060
rect 18700 5020 18740 5060
rect 23308 5020 23348 5060
rect 24652 5020 24692 5060
rect 31756 5020 31796 5060
rect 46348 5020 46388 5060
rect 49420 5020 49460 5060
rect 17644 4936 17684 4976
rect 17932 4936 17972 4976
rect 18316 4936 18356 4976
rect 18604 4936 18644 4976
rect 19180 4936 19220 4976
rect 19564 4936 19604 4976
rect 20428 4936 20468 4976
rect 22924 4936 22964 4976
rect 23212 4936 23252 4976
rect 24748 4936 24788 4976
rect 25036 4936 25076 4976
rect 31660 4936 31700 4976
rect 31852 4936 31892 4976
rect 32716 4936 32756 4976
rect 32908 4936 32948 4976
rect 33100 4936 33140 4976
rect 33484 4936 33524 4976
rect 35020 4936 35060 4976
rect 35116 4936 35156 4976
rect 35212 4936 35252 4976
rect 35404 4936 35444 4976
rect 35500 4936 35540 4976
rect 35596 4936 35636 4976
rect 35692 4936 35732 4976
rect 36076 4936 36116 4976
rect 36172 4936 36212 4976
rect 37612 4936 37652 4976
rect 37996 4936 38036 4976
rect 39628 4922 39668 4962
rect 40108 4936 40148 4976
rect 40588 4936 40628 4976
rect 41068 4936 41108 4976
rect 41164 4936 41204 4976
rect 42892 4936 42932 4976
rect 46444 4936 46484 4976
rect 46732 4936 46772 4976
rect 49324 4936 49364 4976
rect 49516 4936 49556 4976
rect 49900 4936 49940 4976
rect 52204 4936 52244 4976
rect 52492 4936 52532 4976
rect 52588 4936 52628 4976
rect 22444 4852 22484 4892
rect 25900 4852 25940 4892
rect 26284 4852 26324 4892
rect 33196 4852 33236 4892
rect 33388 4852 33428 4892
rect 37708 4852 37748 4892
rect 37900 4852 37940 4892
rect 40684 4852 40724 4892
rect 42412 4852 42452 4892
rect 45196 4852 45236 4892
rect 18988 4768 19028 4808
rect 32812 4768 32852 4808
rect 33292 4768 33332 4808
rect 37804 4768 37844 4808
rect 39244 4768 39284 4808
rect 22636 4684 22676 4724
rect 17260 4642 17300 4682
rect 23596 4684 23636 4724
rect 24364 4684 24404 4724
rect 25708 4684 25748 4724
rect 26092 4684 26132 4724
rect 42220 4684 42260 4724
rect 45388 4684 45428 4724
rect 46060 4684 46100 4724
rect 49708 4684 49748 4724
rect 52876 4684 52916 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 21100 4264 21140 4304
rect 31852 4264 31892 4304
rect 32428 4264 32468 4304
rect 35788 4264 35828 4304
rect 36940 4264 36980 4304
rect 42604 4264 42644 4304
rect 48364 4264 48404 4304
rect 19276 4180 19316 4220
rect 20908 4180 20948 4220
rect 27148 4180 27188 4220
rect 31756 4180 31796 4220
rect 31948 4180 31988 4220
rect 36844 4180 36884 4220
rect 37036 4180 37076 4220
rect 37612 4180 37652 4220
rect 45196 4180 45236 4220
rect 16876 4096 16916 4136
rect 17260 4083 17300 4123
rect 18124 4096 18164 4136
rect 21676 4096 21716 4136
rect 22540 4096 22580 4136
rect 24748 4096 24788 4136
rect 25132 4096 25172 4136
rect 25996 4096 26036 4136
rect 27724 4096 27764 4136
rect 28588 4096 28628 4136
rect 29932 4096 29972 4136
rect 31180 4096 31220 4136
rect 31660 4096 31700 4136
rect 32044 4096 32084 4136
rect 32620 4096 32660 4136
rect 34636 4096 34676 4136
rect 34732 4096 34772 4136
rect 34828 4096 34868 4136
rect 34924 4096 34964 4136
rect 35596 4096 35636 4136
rect 35788 4096 35828 4136
rect 35980 4096 36020 4136
rect 36172 4096 36212 4136
rect 36268 4096 36308 4136
rect 36748 4096 36788 4136
rect 37132 4096 37172 4136
rect 37516 4096 37556 4136
rect 37708 4096 37748 4136
rect 38860 4096 38900 4136
rect 39148 4096 39188 4136
rect 41932 4096 41972 4136
rect 42220 4096 42260 4136
rect 42316 4096 42356 4136
rect 42796 4096 42836 4136
rect 43180 4096 43220 4136
rect 44044 4096 44084 4136
rect 45964 4096 46004 4136
rect 46348 4096 46388 4136
rect 47212 4096 47252 4136
rect 48940 4096 48980 4136
rect 49804 4096 49844 4136
rect 51532 4096 51572 4136
rect 52396 4096 52436 4136
rect 21292 4012 21332 4052
rect 27340 4012 27380 4052
rect 31372 4012 31412 4052
rect 36076 4012 36116 4052
rect 48556 4012 48596 4052
rect 51148 4012 51188 4052
rect 652 3928 692 3968
rect 23692 3928 23732 3968
rect 29740 3928 29780 3968
rect 32716 3928 32756 3968
rect 39052 3928 39092 3968
rect 50956 3928 50996 3968
rect 53548 3928 53588 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 652 3592 692 3632
rect 25708 3592 25748 3632
rect 32716 3592 32756 3632
rect 42892 3592 42932 3632
rect 44716 3592 44756 3632
rect 49036 3592 49076 3632
rect 49324 3592 49364 3632
rect 49516 3592 49556 3632
rect 49804 3592 49844 3632
rect 55084 3592 55124 3632
rect 21580 3508 21620 3548
rect 23308 3508 23348 3548
rect 27244 3508 27284 3548
rect 33868 3508 33908 3548
rect 35884 3508 35924 3548
rect 40012 3508 40052 3548
rect 44236 3508 44276 3548
rect 50860 3508 50900 3548
rect 52684 3508 52724 3548
rect 21196 3424 21236 3464
rect 21484 3424 21524 3464
rect 23692 3424 23732 3464
rect 24556 3424 24596 3464
rect 27340 3451 27380 3491
rect 27628 3424 27668 3464
rect 31276 3424 31316 3464
rect 32524 3424 32564 3464
rect 33484 3424 33524 3464
rect 33772 3424 33812 3464
rect 35500 3424 35540 3464
rect 35788 3424 35828 3464
rect 39052 3424 39092 3464
rect 39148 3424 39188 3464
rect 39244 3424 39284 3464
rect 39628 3424 39668 3464
rect 39916 3424 39956 3464
rect 40492 3424 40532 3464
rect 40876 3424 40916 3464
rect 41740 3424 41780 3464
rect 43852 3424 43892 3464
rect 44140 3424 44180 3464
rect 45868 3424 45908 3464
rect 46732 3424 46772 3464
rect 47116 3424 47156 3464
rect 47980 3424 48020 3464
rect 48268 3424 48308 3464
rect 48364 3424 48404 3464
rect 49228 3424 49268 3464
rect 49708 3424 49748 3464
rect 50476 3424 50516 3464
rect 50764 3424 50804 3464
rect 53068 3424 53108 3464
rect 53932 3424 53972 3464
rect 21868 3256 21908 3296
rect 26956 3256 26996 3296
rect 40300 3256 40340 3296
rect 44524 3256 44564 3296
rect 48652 3256 48692 3296
rect 51148 3256 51188 3296
rect 34156 3172 34196 3212
rect 36172 3172 36212 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 22732 2836 22772 2876
rect 35980 2836 36020 2876
rect 39052 2836 39092 2876
rect 28684 2752 28724 2792
rect 30028 2752 30068 2792
rect 40492 2752 40532 2792
rect 44236 2752 44276 2792
rect 45196 2752 45236 2792
rect 48460 2752 48500 2792
rect 23500 2668 23540 2708
rect 32236 2668 32276 2708
rect 20716 2584 20756 2624
rect 21580 2584 21620 2624
rect 24652 2584 24692 2624
rect 25516 2584 25556 2624
rect 28012 2584 28052 2624
rect 28300 2584 28340 2624
rect 30412 2584 30452 2624
rect 30700 2584 30740 2624
rect 33580 2584 33620 2624
rect 33964 2584 34004 2624
rect 34828 2584 34868 2624
rect 36652 2584 36692 2624
rect 37036 2584 37076 2624
rect 37900 2584 37940 2624
rect 39820 2584 39860 2624
rect 40108 2584 40148 2624
rect 40204 2584 40244 2624
rect 43564 2584 43604 2624
rect 43852 2584 43892 2624
rect 44524 2584 44564 2624
rect 44908 2626 44948 2666
rect 44812 2584 44852 2624
rect 47788 2584 47828 2624
rect 48076 2584 48116 2624
rect 48172 2584 48212 2624
rect 20332 2500 20372 2540
rect 25900 2500 25940 2540
rect 28396 2500 28436 2540
rect 30316 2500 30356 2540
rect 43948 2500 43988 2540
rect 652 2416 692 2456
rect 32428 2416 32468 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 29260 2080 29300 2120
rect 32044 2080 32084 2120
rect 34636 2080 34676 2120
rect 34924 2080 34964 2120
rect 44236 2080 44276 2120
rect 45100 2080 45140 2120
rect 20620 1996 20660 2036
rect 24268 1996 24308 2036
rect 29644 1996 29684 2036
rect 41356 1996 41396 2036
rect 47500 1996 47540 2036
rect 50860 1996 50900 2036
rect 20716 1912 20756 1952
rect 21004 1912 21044 1952
rect 24364 1912 24404 1952
rect 24652 1912 24692 1952
rect 26860 1912 26900 1952
rect 27244 1912 27284 1952
rect 28108 1912 28148 1952
rect 30028 1912 30068 1952
rect 30892 1912 30932 1952
rect 32236 1912 32276 1952
rect 32620 1912 32660 1952
rect 33484 1912 33524 1952
rect 36076 1912 36116 1952
rect 36940 1917 36980 1957
rect 37324 1912 37364 1952
rect 38860 1912 38900 1952
rect 39724 1912 39764 1952
rect 40108 1912 40148 1952
rect 40972 1912 41012 1952
rect 41260 1912 41300 1952
rect 41836 1912 41876 1952
rect 42220 1912 42260 1952
rect 43084 1912 43124 1952
rect 46252 1912 46292 1952
rect 47116 1912 47156 1952
rect 49612 1912 49652 1952
rect 50476 1912 50516 1952
rect 48460 1828 48500 1868
rect 20332 1744 20372 1784
rect 23980 1744 24020 1784
rect 41644 1744 41684 1784
rect 34636 1660 34676 1700
rect 37708 1660 37748 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 26668 1324 26708 1364
rect 30796 1324 30836 1364
rect 32044 1324 32084 1364
rect 35596 1324 35636 1364
rect 38860 1324 38900 1364
rect 40204 1324 40244 1364
rect 44140 1324 44180 1364
rect 47788 1324 47828 1364
rect 47596 1240 47636 1280
rect 26956 1072 26996 1112
rect 27052 1072 27092 1112
rect 27340 1089 27380 1129
rect 28396 1072 28436 1112
rect 28780 1072 28820 1112
rect 29644 1072 29684 1112
rect 32332 1072 32372 1112
rect 32428 1072 32468 1112
rect 32734 1057 32774 1097
rect 34924 1072 34964 1112
rect 35212 1072 35252 1112
rect 35308 1072 35348 1112
rect 38188 1072 38228 1112
rect 38476 1072 38516 1112
rect 38572 1072 38612 1112
rect 41356 1072 41396 1112
rect 42220 1072 42260 1112
rect 42604 1072 42644 1112
rect 45292 1072 45332 1112
rect 46156 1072 46196 1112
rect 46540 1072 46580 1112
rect 46924 1072 46964 1112
rect 47212 1072 47252 1112
rect 47308 1072 47348 1112
rect 48940 1072 48980 1112
rect 49804 1072 49844 1112
rect 50188 1072 50228 1112
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 22060 38408 22100 38417
rect 21868 38368 22060 38408
rect 652 38156 692 38165
rect 652 37577 692 38116
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 21772 37988 21812 37997
rect 844 37854 884 37939
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 651 37568 693 37577
rect 651 37528 652 37568
rect 692 37528 693 37568
rect 651 37519 693 37528
rect 19756 37493 19796 37578
rect 19755 37484 19797 37493
rect 19755 37444 19756 37484
rect 19796 37444 19797 37484
rect 19755 37435 19797 37444
rect 20427 37484 20469 37493
rect 20427 37444 20428 37484
rect 20468 37444 20469 37484
rect 20427 37435 20469 37444
rect 19564 37232 19604 37241
rect 20428 37232 20468 37435
rect 21772 37409 21812 37948
rect 19604 37192 20084 37232
rect 19564 37183 19604 37192
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 13899 36812 13941 36821
rect 13899 36772 13900 36812
rect 13940 36772 13941 36812
rect 20044 36812 20084 37192
rect 20428 37183 20468 37192
rect 20620 37400 20660 37409
rect 20044 36772 20276 36812
rect 13899 36763 13941 36772
rect 7083 36728 7125 36737
rect 7083 36688 7084 36728
rect 7124 36688 7125 36728
rect 7083 36679 7125 36688
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 7084 36065 7124 36679
rect 7083 36056 7125 36065
rect 7083 36016 7084 36056
rect 7124 36016 7125 36056
rect 7083 36007 7125 36016
rect 2379 35888 2421 35897
rect 2379 35848 2380 35888
rect 2420 35848 2421 35888
rect 2379 35839 2421 35848
rect 939 35468 981 35477
rect 939 35428 940 35468
rect 980 35428 981 35468
rect 939 35419 981 35428
rect 652 25388 692 25397
rect 652 24977 692 25348
rect 844 25136 884 25145
rect 748 25096 844 25136
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 652 24548 692 24557
rect 652 24137 692 24508
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 652 23876 692 23885
rect 652 23297 692 23836
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 652 23036 692 23045
rect 652 22457 692 22996
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 652 22112 692 22121
rect 652 21617 692 22072
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 652 20600 692 20719
rect 652 20551 692 20560
rect 652 20264 692 20273
rect 652 19937 692 20224
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18954 692 19039
rect 652 18752 692 18761
rect 652 18257 692 18712
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17576 692 17585
rect 652 17417 692 17536
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 17240 692 17249
rect 652 16577 692 17200
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 652 15594 692 15679
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 652 13880 692 13999
rect 652 13831 692 13840
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 12704 692 13159
rect 652 12655 692 12664
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 652 10638 692 10723
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9260 692 9269
rect 652 9017 692 9220
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 652 8504 692 8513
rect 556 8464 652 8504
rect 556 8177 596 8464
rect 652 8455 692 8464
rect 555 8168 597 8177
rect 555 8128 556 8168
rect 596 8128 597 8168
rect 555 8119 597 8128
rect 652 8168 692 8177
rect 652 7337 692 8128
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 652 5144 692 5153
rect 652 4817 692 5104
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 652 3632 692 3641
rect 652 3137 692 3592
rect 748 3389 788 25096
rect 844 25087 884 25096
rect 843 24800 885 24809
rect 843 24760 844 24800
rect 884 24760 885 24800
rect 843 24751 885 24760
rect 844 24666 884 24751
rect 843 24044 885 24053
rect 843 24004 844 24044
rect 884 24004 885 24044
rect 843 23995 885 24004
rect 844 23910 884 23995
rect 844 23288 884 23297
rect 940 23288 980 35419
rect 884 23248 980 23288
rect 844 23239 884 23248
rect 2283 18668 2325 18677
rect 2283 18628 2284 18668
rect 2324 18628 2325 18668
rect 2283 18619 2325 18628
rect 2187 18584 2229 18593
rect 2187 18544 2188 18584
rect 2228 18544 2229 18584
rect 2187 18535 2229 18544
rect 2092 18332 2132 18341
rect 2188 18332 2228 18535
rect 2284 18500 2324 18619
rect 2284 18451 2324 18460
rect 2132 18292 2228 18332
rect 2092 18283 2132 18292
rect 2091 17324 2133 17333
rect 2091 17284 2092 17324
rect 2132 17284 2133 17324
rect 2091 17275 2133 17284
rect 1323 17240 1365 17249
rect 1323 17200 1324 17240
rect 1364 17200 1365 17240
rect 1323 17191 1365 17200
rect 1228 16232 1268 16241
rect 1324 16232 1364 17191
rect 1803 16484 1845 16493
rect 1803 16444 1804 16484
rect 1844 16444 1845 16484
rect 1803 16435 1845 16444
rect 1268 16192 1364 16232
rect 1228 16183 1268 16192
rect 844 16148 884 16157
rect 844 15401 884 16108
rect 1227 15476 1269 15485
rect 1227 15436 1228 15476
rect 1268 15436 1269 15476
rect 1227 15427 1269 15436
rect 843 15392 885 15401
rect 843 15352 844 15392
rect 884 15352 885 15392
rect 843 15343 885 15352
rect 1228 15342 1268 15427
rect 1036 15308 1076 15317
rect 1036 14897 1076 15268
rect 1035 14888 1077 14897
rect 1035 14848 1036 14888
rect 1076 14848 1077 14888
rect 1035 14839 1077 14848
rect 1228 14720 1268 14729
rect 1324 14720 1364 16192
rect 1804 15644 1844 16435
rect 2092 16232 2132 17275
rect 2092 16183 2132 16192
rect 2188 17072 2228 18292
rect 2284 17576 2324 17585
rect 2284 17249 2324 17536
rect 2283 17240 2325 17249
rect 2283 17200 2284 17240
rect 2324 17200 2325 17240
rect 2283 17191 2325 17200
rect 2284 17072 2324 17081
rect 2188 17032 2284 17072
rect 1804 15595 1844 15604
rect 1900 15560 1940 15569
rect 2188 15560 2228 17032
rect 2284 17023 2324 17032
rect 1515 15392 1557 15401
rect 1515 15352 1516 15392
rect 1556 15352 1557 15392
rect 1515 15343 1557 15352
rect 1516 15258 1556 15343
rect 1900 14897 1940 15520
rect 1996 15520 2188 15560
rect 1611 14888 1653 14897
rect 1611 14848 1612 14888
rect 1652 14848 1653 14888
rect 1611 14839 1653 14848
rect 1899 14888 1941 14897
rect 1899 14848 1900 14888
rect 1940 14848 1941 14888
rect 1899 14839 1941 14848
rect 1268 14680 1460 14720
rect 1228 14671 1268 14680
rect 844 14636 884 14645
rect 884 14596 1172 14636
rect 844 14587 884 14596
rect 844 13964 884 13973
rect 884 13924 980 13964
rect 844 13915 884 13924
rect 844 13124 884 13133
rect 844 12629 884 13084
rect 940 12980 980 13924
rect 1132 13880 1172 14596
rect 1324 13880 1364 13889
rect 1132 13840 1324 13880
rect 1324 13831 1364 13840
rect 1420 13217 1460 14680
rect 1612 14132 1652 14839
rect 1612 14083 1652 14092
rect 1708 14048 1748 14057
rect 1227 13208 1269 13217
rect 1227 13168 1228 13208
rect 1268 13168 1269 13208
rect 1227 13159 1269 13168
rect 1419 13208 1461 13217
rect 1419 13168 1420 13208
rect 1460 13168 1461 13208
rect 1419 13159 1461 13168
rect 1228 13074 1268 13159
rect 940 12940 1172 12980
rect 843 12620 885 12629
rect 843 12580 844 12620
rect 884 12580 885 12620
rect 843 12571 885 12580
rect 844 12452 884 12461
rect 884 12412 980 12452
rect 844 12403 884 12412
rect 940 11864 980 12412
rect 1035 12368 1077 12377
rect 1035 12328 1036 12368
rect 1076 12328 1077 12368
rect 1035 12319 1077 12328
rect 1036 12234 1076 12319
rect 940 11824 1076 11864
rect 844 11780 884 11789
rect 884 11740 980 11780
rect 844 11731 884 11740
rect 843 10940 885 10949
rect 843 10900 844 10940
rect 884 10900 885 10940
rect 843 10891 885 10900
rect 844 10806 884 10891
rect 843 10268 885 10277
rect 843 10228 844 10268
rect 884 10228 885 10268
rect 843 10219 885 10228
rect 844 10134 884 10219
rect 843 9428 885 9437
rect 843 9388 844 9428
rect 884 9388 885 9428
rect 843 9379 885 9388
rect 844 9294 884 9379
rect 940 5489 980 11740
rect 939 5480 981 5489
rect 939 5440 940 5480
rect 980 5440 981 5480
rect 939 5431 981 5440
rect 1036 4817 1076 11824
rect 1132 5573 1172 12940
rect 1419 12620 1461 12629
rect 1419 12580 1420 12620
rect 1460 12580 1461 12620
rect 1419 12571 1461 12580
rect 1228 12452 1268 12461
rect 1228 11696 1268 12412
rect 1420 12368 1460 12571
rect 1420 12319 1460 12328
rect 1708 12536 1748 14008
rect 1996 14048 2036 15520
rect 2188 15511 2228 15520
rect 2091 14720 2133 14729
rect 2091 14680 2092 14720
rect 2132 14680 2133 14720
rect 2091 14671 2133 14680
rect 1996 13049 2036 14008
rect 2092 13208 2132 14671
rect 2092 13159 2132 13168
rect 1995 13040 2037 13049
rect 1995 13000 1996 13040
rect 2036 13000 2037 13040
rect 1995 12991 2037 13000
rect 1708 12293 1748 12496
rect 1803 12536 1845 12545
rect 1803 12496 1804 12536
rect 1844 12496 1845 12536
rect 1996 12536 2036 12991
rect 2380 12980 2420 35839
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 4971 34544 5013 34553
rect 4971 34504 4972 34544
rect 5012 34504 5013 34544
rect 4971 34495 5013 34504
rect 4875 34208 4917 34217
rect 4875 34168 4876 34208
rect 4916 34168 4917 34208
rect 4875 34159 4917 34168
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4876 33140 4916 34159
rect 4780 33100 4916 33140
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4587 32360 4629 32369
rect 4587 32320 4588 32360
rect 4628 32320 4629 32360
rect 4587 32311 4629 32320
rect 4588 32226 4628 32311
rect 2955 32108 2997 32117
rect 2955 32068 2956 32108
rect 2996 32068 2997 32108
rect 2955 32059 2997 32068
rect 4395 32108 4437 32117
rect 4395 32068 4396 32108
rect 4436 32068 4437 32108
rect 4395 32059 4437 32068
rect 2956 23060 2996 32059
rect 4396 31974 4436 32059
rect 4588 31940 4628 31949
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 4588 31361 4628 31900
rect 3819 31352 3861 31361
rect 3819 31312 3820 31352
rect 3860 31312 3861 31352
rect 3819 31303 3861 31312
rect 4587 31352 4629 31361
rect 4587 31312 4588 31352
rect 4628 31312 4629 31352
rect 4587 31303 4629 31312
rect 4684 31352 4724 31361
rect 4780 31352 4820 33100
rect 4972 32369 5012 34495
rect 5739 34376 5781 34385
rect 5739 34336 5740 34376
rect 5780 34336 5781 34376
rect 5739 34327 5781 34336
rect 5163 34040 5205 34049
rect 5163 34000 5164 34040
rect 5204 34000 5205 34040
rect 5163 33991 5205 34000
rect 5164 33140 5204 33991
rect 5068 33100 5204 33140
rect 4971 32360 5013 32369
rect 4971 32320 4972 32360
rect 5012 32320 5013 32360
rect 4971 32311 5013 32320
rect 5068 32108 5108 33100
rect 5547 32948 5589 32957
rect 5547 32908 5548 32948
rect 5588 32908 5589 32948
rect 5547 32899 5589 32908
rect 5548 32814 5588 32899
rect 5356 32696 5396 32705
rect 5259 32612 5301 32621
rect 5259 32572 5260 32612
rect 5300 32572 5301 32612
rect 5259 32563 5301 32572
rect 4724 31312 4820 31352
rect 4684 31303 4724 31312
rect 3436 31268 3476 31277
rect 3436 30521 3476 31228
rect 3435 30512 3477 30521
rect 3435 30472 3436 30512
rect 3476 30472 3477 30512
rect 3435 30463 3477 30472
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3436 28925 3476 29010
rect 3820 29009 3860 31303
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 4491 30764 4533 30773
rect 4491 30724 4492 30764
rect 4532 30724 4533 30764
rect 4491 30715 4533 30724
rect 4492 30630 4532 30715
rect 4587 30680 4629 30689
rect 4587 30640 4588 30680
rect 4628 30640 4629 30680
rect 4587 30631 4629 30640
rect 4588 30546 4628 30631
rect 4203 30512 4245 30521
rect 4203 30472 4204 30512
rect 4244 30472 4245 30512
rect 4203 30463 4245 30472
rect 4204 30378 4244 30463
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 4588 29168 4628 29177
rect 4780 29168 4820 31312
rect 4628 29128 4820 29168
rect 4876 32068 5108 32108
rect 4876 30680 4916 32068
rect 5068 31940 5108 31949
rect 4588 29119 4628 29128
rect 4491 29084 4533 29093
rect 4491 29044 4492 29084
rect 4532 29044 4533 29084
rect 4491 29035 4533 29044
rect 3819 29000 3861 29009
rect 3819 28960 3820 29000
rect 3860 28960 3861 29000
rect 3819 28951 3861 28960
rect 3435 28916 3477 28925
rect 3435 28876 3436 28916
rect 3476 28876 3477 28916
rect 3435 28867 3477 28876
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3435 26144 3477 26153
rect 3435 26104 3436 26144
rect 3476 26104 3477 26144
rect 3435 26095 3477 26104
rect 3820 26144 3860 28951
rect 4492 28328 4532 29035
rect 4492 28169 4532 28288
rect 4491 28160 4533 28169
rect 4491 28120 4492 28160
rect 4532 28120 4533 28160
rect 4684 28160 4724 29128
rect 4876 29093 4916 30640
rect 4972 31900 5068 31940
rect 4875 29084 4917 29093
rect 4875 29044 4876 29084
rect 4916 29044 4917 29084
rect 4875 29035 4917 29044
rect 4875 28916 4917 28925
rect 4875 28876 4876 28916
rect 4916 28876 4917 28916
rect 4875 28867 4917 28876
rect 4780 28337 4820 28422
rect 4779 28328 4821 28337
rect 4779 28288 4780 28328
rect 4820 28288 4821 28328
rect 4779 28279 4821 28288
rect 4876 28253 4916 28867
rect 4875 28244 4917 28253
rect 4875 28204 4876 28244
rect 4916 28204 4917 28244
rect 4875 28195 4917 28204
rect 4684 28120 4820 28160
rect 4491 28111 4533 28120
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3436 26010 3476 26095
rect 3627 25976 3669 25985
rect 3627 25936 3628 25976
rect 3668 25936 3669 25976
rect 3627 25927 3669 25936
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 3435 23708 3477 23717
rect 3435 23668 3436 23708
rect 3476 23668 3477 23708
rect 3435 23659 3477 23668
rect 3436 23574 3476 23659
rect 3532 23129 3572 23214
rect 3531 23120 3573 23129
rect 3531 23080 3532 23120
rect 3572 23080 3573 23120
rect 3531 23071 3573 23080
rect 3628 23120 3668 25927
rect 2860 23020 2996 23060
rect 2860 19340 2900 23020
rect 3244 22868 3284 22877
rect 3284 22828 3572 22868
rect 3244 22819 3284 22828
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 3339 22448 3381 22457
rect 3339 22408 3340 22448
rect 3380 22408 3381 22448
rect 3339 22399 3381 22408
rect 3340 21701 3380 22399
rect 3436 22280 3476 22289
rect 3532 22280 3572 22828
rect 3628 22457 3668 23080
rect 3820 23792 3860 26104
rect 4203 26144 4245 26153
rect 4203 26104 4204 26144
rect 4244 26104 4245 26144
rect 4203 26095 4245 26104
rect 4684 26144 4724 26153
rect 4780 26144 4820 28120
rect 4876 28110 4916 28195
rect 4875 27992 4917 28001
rect 4875 27952 4876 27992
rect 4916 27952 4917 27992
rect 4875 27943 4917 27952
rect 4724 26104 4820 26144
rect 4684 26095 4724 26104
rect 4204 25556 4244 26095
rect 4491 25892 4533 25901
rect 4491 25852 4492 25892
rect 4532 25852 4533 25892
rect 4491 25843 4533 25852
rect 4204 25507 4244 25516
rect 4492 25304 4532 25843
rect 4492 25255 4532 25264
rect 4587 25304 4629 25313
rect 4587 25264 4588 25304
rect 4628 25264 4629 25304
rect 4587 25255 4629 25264
rect 4588 25170 4628 25255
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 3627 22448 3669 22457
rect 3627 22408 3628 22448
rect 3668 22408 3669 22448
rect 3627 22399 3669 22408
rect 3820 22280 3860 23752
rect 4684 23792 4724 23801
rect 4780 23792 4820 26104
rect 4724 23752 4820 23792
rect 4684 23743 4724 23752
rect 4203 23708 4245 23717
rect 4203 23668 4204 23708
rect 4244 23668 4245 23708
rect 4203 23659 4245 23668
rect 3915 23372 3957 23381
rect 3915 23332 3916 23372
rect 3956 23332 3957 23372
rect 3915 23323 3957 23332
rect 4204 23330 4244 23659
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3476 22240 3572 22280
rect 3628 22240 3820 22280
rect 3436 22231 3476 22240
rect 3339 21692 3381 21701
rect 3339 21652 3340 21692
rect 3380 21652 3381 21692
rect 3339 21643 3381 21652
rect 3340 21558 3380 21643
rect 3435 21608 3477 21617
rect 3435 21568 3436 21608
rect 3476 21568 3477 21608
rect 3435 21559 3477 21568
rect 3436 21474 3476 21559
rect 3052 21356 3092 21365
rect 2956 21316 3052 21356
rect 2956 20768 2996 21316
rect 3052 21307 3092 21316
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 2956 20719 2996 20728
rect 3340 20768 3380 20777
rect 3628 20768 3668 22240
rect 3820 22231 3860 22240
rect 3916 23120 3956 23323
rect 4204 23281 4244 23290
rect 4587 23288 4629 23297
rect 4780 23288 4820 23752
rect 4876 25304 4916 27943
rect 4876 23549 4916 25264
rect 4875 23540 4917 23549
rect 4875 23500 4876 23540
rect 4916 23500 4917 23540
rect 4875 23491 4917 23500
rect 4587 23248 4588 23288
rect 4628 23248 4629 23288
rect 4587 23239 4629 23248
rect 4684 23248 4820 23288
rect 4491 23204 4533 23213
rect 4491 23164 4492 23204
rect 4532 23164 4533 23204
rect 4491 23155 4533 23164
rect 3724 21608 3764 21617
rect 3916 21608 3956 23080
rect 4492 23070 4532 23155
rect 4588 23129 4628 23239
rect 4587 23120 4629 23129
rect 4587 23080 4588 23120
rect 4628 23080 4629 23120
rect 4587 23071 4629 23080
rect 4684 22280 4724 23248
rect 4779 23120 4821 23129
rect 4779 23080 4780 23120
rect 4820 23080 4821 23120
rect 4779 23071 4821 23080
rect 4876 23120 4916 23491
rect 4876 23071 4916 23080
rect 4684 22231 4724 22240
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3764 21568 4052 21608
rect 3724 21559 3764 21568
rect 3380 20728 3860 20768
rect 3340 20719 3380 20728
rect 3436 20096 3476 20105
rect 3820 20096 3860 20728
rect 3476 20056 3572 20096
rect 3436 20047 3476 20056
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3532 19508 3572 20056
rect 3820 20047 3860 20056
rect 3915 20012 3957 20021
rect 3915 19972 3916 20012
rect 3956 19972 3957 20012
rect 3915 19963 3957 19972
rect 3628 19508 3668 19517
rect 3532 19468 3628 19508
rect 3628 19459 3668 19468
rect 2860 19291 2900 19300
rect 3436 19340 3476 19349
rect 3476 19300 3860 19340
rect 3436 19291 3476 19300
rect 2955 19088 2997 19097
rect 2955 19048 2956 19088
rect 2996 19048 2997 19088
rect 2955 19039 2997 19048
rect 3052 19088 3092 19097
rect 2956 18668 2996 19039
rect 2956 18619 2996 18628
rect 2571 18584 2613 18593
rect 2571 18544 2572 18584
rect 2612 18544 2613 18584
rect 2571 18535 2613 18544
rect 2860 18584 2900 18593
rect 2572 18450 2612 18535
rect 2860 17921 2900 18544
rect 3052 18332 3092 19048
rect 3244 19088 3284 19097
rect 3244 18677 3284 19048
rect 3820 18752 3860 19300
rect 3916 19256 3956 19963
rect 4012 19937 4052 21568
rect 4203 20768 4245 20777
rect 4203 20728 4204 20768
rect 4244 20728 4245 20768
rect 4203 20719 4245 20728
rect 4204 20180 4244 20719
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4204 20140 4724 20180
rect 4011 19928 4053 19937
rect 4011 19888 4012 19928
rect 4052 19888 4053 19928
rect 4011 19879 4053 19888
rect 3916 19207 3956 19216
rect 4012 19256 4052 19265
rect 4012 19097 4052 19216
rect 4011 19088 4053 19097
rect 4011 19048 4012 19088
rect 4052 19048 4053 19088
rect 4011 19039 4053 19048
rect 3820 18712 4148 18752
rect 3243 18668 3285 18677
rect 3243 18628 3244 18668
rect 3284 18628 3285 18668
rect 3243 18619 3285 18628
rect 3436 18584 3476 18593
rect 3244 18416 3284 18425
rect 3436 18416 3476 18544
rect 3284 18376 3476 18416
rect 3820 18584 3860 18593
rect 3244 18367 3284 18376
rect 2956 18292 3092 18332
rect 2571 17912 2613 17921
rect 2571 17872 2572 17912
rect 2612 17872 2613 17912
rect 2571 17863 2613 17872
rect 2859 17912 2901 17921
rect 2859 17872 2860 17912
rect 2900 17872 2901 17912
rect 2859 17863 2901 17872
rect 2475 17828 2517 17837
rect 2475 17788 2476 17828
rect 2516 17788 2517 17828
rect 2475 17779 2517 17788
rect 2476 17694 2516 17779
rect 2572 17300 2612 17863
rect 2668 17660 2708 17669
rect 2708 17620 2900 17660
rect 2668 17611 2708 17620
rect 2572 17260 2708 17300
rect 2668 17156 2708 17260
rect 2668 17107 2708 17116
rect 2572 17072 2612 17081
rect 2572 16493 2612 17032
rect 2860 16904 2900 17620
rect 2956 17072 2996 18292
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3820 17837 3860 18544
rect 3915 18584 3957 18593
rect 3915 18544 3916 18584
rect 3956 18544 3957 18584
rect 3915 18535 3957 18544
rect 3819 17828 3861 17837
rect 3819 17788 3820 17828
rect 3860 17788 3861 17828
rect 3819 17779 3861 17788
rect 3052 17744 3092 17753
rect 3052 17249 3092 17704
rect 3051 17240 3093 17249
rect 3051 17200 3052 17240
rect 3092 17200 3093 17240
rect 3051 17191 3093 17200
rect 2956 17032 3092 17072
rect 2956 16904 2996 16913
rect 2860 16864 2956 16904
rect 2956 16855 2996 16864
rect 3052 16778 3092 17032
rect 3244 16988 3284 16997
rect 3244 16778 3284 16948
rect 2956 16738 3284 16778
rect 3436 16820 3476 16829
rect 3820 16820 3860 17779
rect 3916 17744 3956 18535
rect 3916 17333 3956 17704
rect 3915 17324 3957 17333
rect 3915 17284 3916 17324
rect 3956 17284 3957 17324
rect 3915 17275 3957 17284
rect 3915 16904 3957 16913
rect 3915 16864 3916 16904
rect 3956 16864 3957 16904
rect 3915 16855 3957 16864
rect 3476 16780 3860 16820
rect 3436 16771 3476 16780
rect 2571 16484 2613 16493
rect 2571 16444 2572 16484
rect 2612 16444 2613 16484
rect 2571 16435 2613 16444
rect 2956 15401 2996 16738
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 3243 16484 3285 16493
rect 3243 16444 3244 16484
rect 3284 16444 3285 16484
rect 3243 16435 3285 16444
rect 3244 16350 3284 16435
rect 3820 16232 3860 16780
rect 3916 16493 3956 16855
rect 3915 16484 3957 16493
rect 3915 16444 3916 16484
rect 3956 16444 3957 16484
rect 3915 16435 3957 16444
rect 3860 16192 4052 16232
rect 3820 16183 3860 16192
rect 3436 16148 3476 16157
rect 3436 15485 3476 16108
rect 3435 15476 3477 15485
rect 3435 15436 3436 15476
rect 3476 15436 3477 15476
rect 3435 15427 3477 15436
rect 2955 15392 2997 15401
rect 2955 15352 2956 15392
rect 2996 15352 2997 15392
rect 2955 15343 2997 15352
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 3243 14888 3285 14897
rect 3243 14848 3244 14888
rect 3284 14848 3285 14888
rect 3243 14839 3285 14848
rect 3244 14754 3284 14839
rect 3820 14720 3860 14729
rect 3724 14680 3820 14720
rect 3436 14636 3476 14645
rect 3436 13880 3476 14596
rect 3532 13880 3572 13889
rect 3436 13840 3532 13880
rect 3532 13831 3572 13840
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 3724 13217 3764 14680
rect 3820 14671 3860 14680
rect 3819 14552 3861 14561
rect 3819 14512 3820 14552
rect 3860 14512 3861 14552
rect 3819 14503 3861 14512
rect 3820 14132 3860 14503
rect 3820 14083 3860 14092
rect 3916 14048 3956 14057
rect 3723 13208 3765 13217
rect 3820 13208 3860 13217
rect 3723 13168 3724 13208
rect 3764 13168 3820 13208
rect 3723 13159 3765 13168
rect 3820 13159 3860 13168
rect 3436 13124 3476 13133
rect 2571 13040 2613 13049
rect 2571 13000 2572 13040
rect 2612 13000 2613 13040
rect 2571 12991 2613 13000
rect 3244 13040 3284 13049
rect 2188 12940 2420 12980
rect 2092 12536 2132 12545
rect 1996 12496 2092 12536
rect 1803 12487 1845 12496
rect 2092 12487 2132 12496
rect 1804 12402 1844 12487
rect 1707 12284 1749 12293
rect 1707 12244 1708 12284
rect 1748 12244 1749 12284
rect 1707 12235 1749 12244
rect 1228 11656 1460 11696
rect 1420 6497 1460 11656
rect 1803 10940 1845 10949
rect 1803 10900 1804 10940
rect 1844 10900 1845 10940
rect 1803 10891 1845 10900
rect 1804 6749 1844 10891
rect 1899 10268 1941 10277
rect 1899 10228 1900 10268
rect 1940 10228 1941 10268
rect 1899 10219 1941 10228
rect 1803 6740 1845 6749
rect 1803 6700 1804 6740
rect 1844 6700 1845 6740
rect 1803 6691 1845 6700
rect 1900 6665 1940 10219
rect 2188 7169 2228 12940
rect 2475 12536 2517 12545
rect 2475 12496 2476 12536
rect 2516 12496 2517 12536
rect 2475 12487 2517 12496
rect 2476 11528 2516 12487
rect 2572 11696 2612 12991
rect 2763 12788 2805 12797
rect 2763 12748 2764 12788
rect 2804 12748 2805 12788
rect 2763 12739 2805 12748
rect 2764 12116 2804 12739
rect 2955 12368 2997 12377
rect 2955 12328 2956 12368
rect 2996 12328 2997 12368
rect 2955 12319 2997 12328
rect 2764 12076 2900 12116
rect 2860 11738 2900 12076
rect 2860 11689 2900 11698
rect 2956 11696 2996 12319
rect 3244 12293 3284 13000
rect 3436 12980 3476 13084
rect 3436 12940 3572 12980
rect 3532 12368 3572 12940
rect 3532 12319 3572 12328
rect 3243 12284 3285 12293
rect 3243 12244 3244 12284
rect 3284 12244 3285 12284
rect 3243 12235 3285 12244
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3244 11864 3284 11873
rect 3284 11824 3476 11864
rect 3244 11815 3284 11824
rect 2572 11647 2612 11656
rect 2956 11647 2996 11656
rect 3436 11696 3476 11824
rect 3724 11696 3764 13159
rect 3916 12713 3956 14008
rect 3915 12704 3957 12713
rect 3820 12664 3916 12704
rect 3956 12664 3957 12704
rect 3820 12620 3860 12664
rect 3915 12655 3957 12664
rect 3820 12571 3860 12580
rect 3916 12536 3956 12545
rect 3916 12377 3956 12496
rect 3915 12368 3957 12377
rect 3915 12328 3916 12368
rect 3956 12328 3957 12368
rect 3915 12319 3957 12328
rect 3820 11696 3860 11705
rect 3436 11647 3476 11656
rect 3628 11656 3820 11696
rect 2476 11488 2612 11528
rect 2476 11024 2516 11033
rect 2284 10436 2324 10445
rect 2476 10436 2516 10984
rect 2324 10396 2516 10436
rect 2284 10387 2324 10396
rect 2572 10184 2612 11488
rect 2908 11024 2948 11033
rect 3628 11024 3668 11656
rect 3820 11647 3860 11656
rect 3723 11528 3765 11537
rect 3723 11488 3724 11528
rect 3764 11488 3765 11528
rect 3723 11479 3765 11488
rect 2948 10984 3668 11024
rect 3724 11024 3764 11479
rect 2908 10975 2948 10984
rect 3724 10975 3764 10984
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3916 10352 3956 10361
rect 3436 10312 3916 10352
rect 2572 10135 2612 10144
rect 2667 10184 2709 10193
rect 2667 10144 2668 10184
rect 2708 10144 2709 10184
rect 2667 10135 2709 10144
rect 2955 10184 2997 10193
rect 2955 10144 2956 10184
rect 2996 10144 2997 10184
rect 2955 10135 2997 10144
rect 2668 10050 2708 10135
rect 2956 10050 2996 10135
rect 3436 9596 3476 10312
rect 3916 10303 3956 10312
rect 3436 9547 3476 9556
rect 3820 9512 3860 9521
rect 4012 9512 4052 16192
rect 4108 15644 4148 18712
rect 4204 18593 4244 20140
rect 4684 20096 4724 20140
rect 4684 20047 4724 20056
rect 4299 19928 4341 19937
rect 4299 19888 4300 19928
rect 4340 19888 4341 19928
rect 4299 19879 4341 19888
rect 4300 19256 4340 19879
rect 4300 19207 4340 19216
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4203 18584 4245 18593
rect 4203 18544 4204 18584
rect 4244 18544 4245 18584
rect 4203 18535 4245 18544
rect 4683 18584 4725 18593
rect 4683 18544 4684 18584
rect 4724 18544 4725 18584
rect 4683 18535 4725 18544
rect 4684 18450 4724 18535
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4658 17300 4700 17309
rect 4658 17260 4659 17300
rect 4699 17260 4724 17300
rect 4658 17251 4724 17260
rect 4684 16232 4724 17251
rect 4684 16183 4724 16192
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4491 15644 4533 15653
rect 4108 15604 4340 15644
rect 4203 15476 4245 15485
rect 4203 15436 4204 15476
rect 4244 15436 4245 15476
rect 4203 15427 4245 15436
rect 4107 15392 4149 15401
rect 4107 15352 4108 15392
rect 4148 15352 4149 15392
rect 4107 15343 4149 15352
rect 4204 15392 4244 15427
rect 3860 9472 4052 9512
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3435 8000 3477 8009
rect 3435 7960 3436 8000
rect 3476 7960 3477 8000
rect 3435 7951 3477 7960
rect 3820 8000 3860 9472
rect 3820 7951 3860 7960
rect 3436 7866 3476 7951
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 2187 7160 2229 7169
rect 2187 7120 2188 7160
rect 2228 7120 2229 7160
rect 2187 7111 2229 7120
rect 1899 6656 1941 6665
rect 1899 6616 1900 6656
rect 1940 6616 1941 6656
rect 1899 6607 1941 6616
rect 1419 6488 1461 6497
rect 1419 6448 1420 6488
rect 1460 6448 1461 6488
rect 1419 6439 1461 6448
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 1131 5564 1173 5573
rect 1131 5524 1132 5564
rect 1172 5524 1173 5564
rect 1131 5515 1173 5524
rect 1035 4808 1077 4817
rect 1035 4768 1036 4808
rect 1076 4768 1077 4808
rect 1035 4759 1077 4768
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 4108 3725 4148 15343
rect 4204 15341 4244 15352
rect 4300 15224 4340 15604
rect 4491 15604 4492 15644
rect 4532 15604 4533 15644
rect 4491 15595 4533 15604
rect 4492 15510 4532 15595
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 4204 15184 4340 15224
rect 4204 14225 4244 15184
rect 4588 14561 4628 15511
rect 4683 14720 4725 14729
rect 4683 14680 4684 14720
rect 4724 14680 4725 14720
rect 4683 14671 4725 14680
rect 4684 14586 4724 14671
rect 4587 14552 4629 14561
rect 4587 14512 4588 14552
rect 4628 14512 4629 14552
rect 4587 14503 4629 14512
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4203 14216 4245 14225
rect 4203 14176 4204 14216
rect 4244 14176 4245 14216
rect 4203 14167 4245 14176
rect 4204 14048 4244 14057
rect 4204 13049 4244 14008
rect 4683 13208 4725 13217
rect 4683 13168 4684 13208
rect 4724 13168 4725 13208
rect 4683 13159 4725 13168
rect 4684 13074 4724 13159
rect 4203 13040 4245 13049
rect 4203 13000 4204 13040
rect 4244 13000 4245 13040
rect 4203 12991 4245 13000
rect 4204 12536 4244 12991
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4204 12487 4244 12496
rect 4299 11696 4341 11705
rect 4299 11656 4300 11696
rect 4340 11656 4341 11696
rect 4299 11647 4341 11656
rect 4684 11696 4724 11705
rect 4300 11528 4340 11647
rect 4684 11537 4724 11656
rect 4204 11488 4340 11528
rect 4683 11528 4725 11537
rect 4683 11488 4684 11528
rect 4724 11488 4725 11528
rect 4204 11192 4244 11488
rect 4683 11479 4725 11488
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4204 11152 4340 11192
rect 4300 10184 4340 11152
rect 4300 10135 4340 10144
rect 4587 10184 4629 10193
rect 4587 10144 4588 10184
rect 4628 10144 4629 10184
rect 4587 10135 4629 10144
rect 4203 10100 4245 10109
rect 4203 10060 4204 10100
rect 4244 10060 4245 10100
rect 4203 10051 4245 10060
rect 4204 9966 4244 10051
rect 4588 10050 4628 10135
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4684 9512 4724 9521
rect 4780 9512 4820 23071
rect 4972 20777 5012 31900
rect 5068 31891 5108 31900
rect 5067 30680 5109 30689
rect 5067 30640 5068 30680
rect 5108 30640 5109 30680
rect 5067 30631 5109 30640
rect 5068 25472 5108 30631
rect 5163 29168 5205 29177
rect 5163 29128 5164 29168
rect 5204 29128 5205 29168
rect 5163 29119 5205 29128
rect 5164 28580 5204 29119
rect 5164 28531 5204 28540
rect 5068 25432 5204 25472
rect 5067 25304 5109 25313
rect 5067 25264 5068 25304
rect 5108 25264 5109 25304
rect 5067 25255 5109 25264
rect 5068 21953 5108 25255
rect 5164 24053 5204 25432
rect 5163 24044 5205 24053
rect 5163 24004 5164 24044
rect 5204 24004 5205 24044
rect 5163 23995 5205 24004
rect 5164 23381 5204 23995
rect 5163 23372 5205 23381
rect 5163 23332 5164 23372
rect 5204 23332 5205 23372
rect 5163 23323 5205 23332
rect 5260 23213 5300 32563
rect 5356 32117 5396 32656
rect 5740 32192 5780 34327
rect 6411 32444 6453 32453
rect 6411 32404 6412 32444
rect 6452 32404 6453 32444
rect 6411 32395 6453 32404
rect 5740 32143 5780 32152
rect 5355 32108 5397 32117
rect 5355 32068 5356 32108
rect 5396 32068 5397 32108
rect 5355 32059 5397 32068
rect 5835 31604 5877 31613
rect 5835 31564 5836 31604
rect 5876 31564 5877 31604
rect 5835 31555 5877 31564
rect 5836 31470 5876 31555
rect 5931 31520 5973 31529
rect 5931 31480 5932 31520
rect 5972 31480 5973 31520
rect 5931 31471 5973 31480
rect 5836 31184 5876 31193
rect 5836 30773 5876 31144
rect 5835 30764 5877 30773
rect 5835 30724 5836 30764
rect 5876 30724 5877 30764
rect 5835 30715 5877 30724
rect 5452 29168 5492 29177
rect 5452 29009 5492 29128
rect 5835 29168 5877 29177
rect 5835 29128 5836 29168
rect 5876 29128 5877 29168
rect 5835 29119 5877 29128
rect 5836 29034 5876 29119
rect 5451 29000 5493 29009
rect 5451 28960 5452 29000
rect 5492 28960 5493 29000
rect 5451 28951 5493 28960
rect 5355 28244 5397 28253
rect 5355 28204 5356 28244
rect 5396 28204 5397 28244
rect 5355 28195 5397 28204
rect 5259 23204 5301 23213
rect 5259 23164 5260 23204
rect 5300 23164 5301 23204
rect 5259 23155 5301 23164
rect 5356 23060 5396 28195
rect 5836 26312 5876 26321
rect 5932 26312 5972 31471
rect 5876 26272 5972 26312
rect 5836 26263 5876 26272
rect 5835 25892 5877 25901
rect 5835 25852 5836 25892
rect 5876 25852 5877 25892
rect 5835 25843 5877 25852
rect 5836 25758 5876 25843
rect 5835 24044 5877 24053
rect 5835 24004 5836 24044
rect 5876 24004 5877 24044
rect 5835 23995 5877 24004
rect 5836 23910 5876 23995
rect 5739 23372 5781 23381
rect 5739 23332 5740 23372
rect 5780 23332 5781 23372
rect 5739 23323 5781 23332
rect 5260 23020 5396 23060
rect 5067 21944 5109 21953
rect 5067 21904 5068 21944
rect 5108 21904 5109 21944
rect 5067 21895 5109 21904
rect 4971 20768 5013 20777
rect 4971 20728 4972 20768
rect 5012 20728 5013 20768
rect 4971 20719 5013 20728
rect 5068 20021 5108 21895
rect 5067 20012 5109 20021
rect 5067 19972 5068 20012
rect 5108 19972 5109 20012
rect 5067 19963 5109 19972
rect 4971 18668 5013 18677
rect 4971 18628 4972 18668
rect 5012 18628 5013 18668
rect 4971 18619 5013 18628
rect 4876 15560 4916 15569
rect 4972 15560 5012 18619
rect 5067 17912 5109 17921
rect 5067 17872 5068 17912
rect 5108 17872 5109 17912
rect 5067 17863 5109 17872
rect 5068 17778 5108 17863
rect 4916 15520 5204 15560
rect 4876 15511 4916 15520
rect 4875 14720 4917 14729
rect 4875 14680 4876 14720
rect 4916 14680 4917 14720
rect 4875 14671 4917 14680
rect 4876 13217 4916 14671
rect 5067 14216 5109 14225
rect 5067 14176 5068 14216
rect 5108 14176 5109 14216
rect 5067 14167 5109 14176
rect 4875 13208 4917 13217
rect 4875 13168 4876 13208
rect 4916 13168 4917 13208
rect 4875 13159 4917 13168
rect 4876 11537 4916 13159
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 4971 12487 5013 12496
rect 4875 11528 4917 11537
rect 4875 11488 4876 11528
rect 4916 11488 4917 11528
rect 4875 11479 4917 11488
rect 4876 11192 4916 11201
rect 4972 11192 5012 12487
rect 4916 11152 5012 11192
rect 4876 11143 4916 11152
rect 4971 10184 5013 10193
rect 4971 10144 4972 10184
rect 5012 10144 5013 10184
rect 4971 10135 5013 10144
rect 4724 9472 4820 9512
rect 4684 9463 4724 9472
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4587 8168 4629 8177
rect 4587 8128 4588 8168
rect 4628 8128 4629 8168
rect 4587 8119 4629 8128
rect 4299 8000 4341 8009
rect 4299 7960 4300 8000
rect 4340 7960 4341 8000
rect 4299 7951 4341 7960
rect 4300 7412 4340 7951
rect 4300 7363 4340 7372
rect 4588 7160 4628 8119
rect 4683 8000 4725 8009
rect 4780 8000 4820 9472
rect 4683 7960 4684 8000
rect 4724 7960 4820 8000
rect 4683 7951 4725 7960
rect 4684 7866 4724 7951
rect 4588 7111 4628 7120
rect 4684 7160 4724 7169
rect 4684 6992 4724 7120
rect 4972 7160 5012 10135
rect 4972 7111 5012 7120
rect 4684 6952 4820 6992
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 4780 5405 4820 6952
rect 4779 5396 4821 5405
rect 4779 5356 4780 5396
rect 4820 5356 4821 5396
rect 4779 5347 4821 5356
rect 5068 5321 5108 14167
rect 5164 10193 5204 15520
rect 5260 12041 5300 23020
rect 5355 21692 5397 21701
rect 5355 21652 5356 21692
rect 5396 21652 5397 21692
rect 5355 21643 5397 21652
rect 5356 21020 5396 21643
rect 5356 20971 5396 20980
rect 5740 20945 5780 23323
rect 5835 23288 5877 23297
rect 5835 23248 5836 23288
rect 5876 23248 5877 23288
rect 5835 23239 5877 23248
rect 5836 22532 5876 23239
rect 5836 22483 5876 22492
rect 5836 22112 5876 22121
rect 5876 22072 5972 22112
rect 5836 22063 5876 22072
rect 5739 20936 5781 20945
rect 5739 20896 5740 20936
rect 5780 20896 5781 20936
rect 5739 20887 5781 20896
rect 5835 20012 5877 20021
rect 5835 19972 5836 20012
rect 5876 19972 5877 20012
rect 5835 19963 5877 19972
rect 5836 19878 5876 19963
rect 5835 19088 5877 19097
rect 5835 19048 5836 19088
rect 5876 19048 5877 19088
rect 5835 19039 5877 19048
rect 5836 18500 5876 19039
rect 5932 18929 5972 22072
rect 5931 18920 5973 18929
rect 5931 18880 5932 18920
rect 5972 18880 5973 18920
rect 5931 18871 5973 18880
rect 5836 18451 5876 18460
rect 5835 16736 5877 16745
rect 5835 16696 5836 16736
rect 5876 16696 5877 16736
rect 5835 16687 5877 16696
rect 5836 16484 5876 16687
rect 5931 16568 5973 16577
rect 5931 16528 5932 16568
rect 5972 16528 5973 16568
rect 5931 16519 5973 16528
rect 5836 16435 5876 16444
rect 5836 16064 5876 16073
rect 5836 15653 5876 16024
rect 5835 15644 5877 15653
rect 5835 15604 5836 15644
rect 5876 15604 5877 15644
rect 5835 15595 5877 15604
rect 5932 15569 5972 16519
rect 5931 15560 5973 15569
rect 5931 15520 5932 15560
rect 5972 15520 5973 15560
rect 5931 15511 5973 15520
rect 5836 14972 5876 14981
rect 5932 14972 5972 15511
rect 5876 14932 5972 14972
rect 5836 14923 5876 14932
rect 6412 14729 6452 32395
rect 6411 14720 6453 14729
rect 6411 14680 6412 14720
rect 6452 14680 6453 14720
rect 6411 14671 6453 14680
rect 5836 13040 5876 13049
rect 5739 12788 5781 12797
rect 5739 12748 5740 12788
rect 5780 12748 5781 12788
rect 5739 12739 5781 12748
rect 5259 12032 5301 12041
rect 5259 11992 5260 12032
rect 5300 11992 5301 12032
rect 5259 11983 5301 11992
rect 5260 11705 5300 11983
rect 5259 11696 5301 11705
rect 5259 11656 5260 11696
rect 5300 11656 5301 11696
rect 5259 11647 5301 11656
rect 5163 10184 5205 10193
rect 5163 10144 5164 10184
rect 5204 10144 5205 10184
rect 5163 10135 5205 10144
rect 5740 8177 5780 12739
rect 5836 12713 5876 13000
rect 5835 12704 5877 12713
rect 5835 12664 5836 12704
rect 5876 12664 5877 12704
rect 5835 12655 5877 12664
rect 5835 12368 5877 12377
rect 5835 12328 5836 12368
rect 5876 12328 5877 12368
rect 5835 12319 5877 12328
rect 5836 11948 5876 12319
rect 5836 11899 5876 11908
rect 5835 10100 5877 10109
rect 5835 10060 5836 10100
rect 5876 10060 5877 10100
rect 5835 10051 5877 10060
rect 5836 9680 5876 10051
rect 5836 9631 5876 9640
rect 5836 9260 5876 9269
rect 5876 9220 5972 9260
rect 5836 9211 5876 9220
rect 5739 8168 5781 8177
rect 5836 8168 5876 8177
rect 5739 8128 5740 8168
rect 5780 8128 5836 8168
rect 5739 8119 5781 8128
rect 5836 8119 5876 8128
rect 5740 8034 5780 8119
rect 5163 8000 5205 8009
rect 5163 7960 5164 8000
rect 5204 7960 5205 8000
rect 5163 7951 5205 7960
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 5067 5312 5109 5321
rect 5067 5272 5068 5312
rect 5108 5272 5109 5312
rect 5067 5263 5109 5272
rect 5164 4145 5204 7951
rect 5932 7001 5972 9220
rect 5931 6992 5973 7001
rect 5931 6952 5932 6992
rect 5972 6952 5973 6992
rect 5931 6943 5973 6952
rect 7084 4985 7124 36007
rect 13900 35972 13940 36763
rect 18699 36728 18741 36737
rect 19084 36728 19124 36737
rect 18699 36688 18700 36728
rect 18740 36688 18741 36728
rect 18699 36679 18741 36688
rect 18988 36688 19084 36728
rect 18700 36594 18740 36679
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 13803 35720 13845 35729
rect 13803 35680 13804 35720
rect 13844 35680 13845 35720
rect 13803 35671 13845 35680
rect 8139 35636 8181 35645
rect 8139 35596 8140 35636
rect 8180 35596 8181 35636
rect 8139 35587 8181 35596
rect 7275 34544 7317 34553
rect 7275 34504 7276 34544
rect 7316 34504 7317 34544
rect 7275 34495 7317 34504
rect 7563 34544 7605 34553
rect 7563 34504 7564 34544
rect 7604 34504 7605 34544
rect 7563 34495 7605 34504
rect 7276 34133 7316 34495
rect 7564 34410 7604 34495
rect 7851 34376 7893 34385
rect 7851 34336 7852 34376
rect 7892 34336 7893 34376
rect 7851 34327 7893 34336
rect 7852 34242 7892 34327
rect 7371 34208 7413 34217
rect 7371 34168 7372 34208
rect 7412 34168 7413 34208
rect 7371 34159 7413 34168
rect 7275 34124 7317 34133
rect 7275 34084 7276 34124
rect 7316 34084 7317 34124
rect 7275 34075 7317 34084
rect 7372 34074 7412 34159
rect 7947 33704 7989 33713
rect 7947 33664 7948 33704
rect 7988 33664 7989 33704
rect 7947 33655 7989 33664
rect 7948 7085 7988 33655
rect 7947 7076 7989 7085
rect 7947 7036 7948 7076
rect 7988 7036 7989 7076
rect 7947 7027 7989 7036
rect 7083 4976 7125 4985
rect 7083 4936 7084 4976
rect 7124 4936 7125 4976
rect 7083 4927 7125 4936
rect 8140 4313 8180 35587
rect 13228 35216 13268 35225
rect 10635 35132 10677 35141
rect 10635 35092 10636 35132
rect 10676 35092 10677 35132
rect 10635 35083 10677 35092
rect 10444 34964 10484 34973
rect 9964 34376 10004 34385
rect 9964 34049 10004 34336
rect 10252 34376 10292 34385
rect 10252 34217 10292 34336
rect 10348 34292 10388 34301
rect 10251 34208 10293 34217
rect 10251 34168 10252 34208
rect 10292 34168 10293 34208
rect 10251 34159 10293 34168
rect 9963 34040 10005 34049
rect 9963 34000 9964 34040
rect 10004 34000 10005 34040
rect 9963 33991 10005 34000
rect 8331 33956 8373 33965
rect 8331 33916 8332 33956
rect 8372 33916 8373 33956
rect 8331 33907 8373 33916
rect 8235 33872 8277 33881
rect 8235 33832 8236 33872
rect 8276 33832 8277 33872
rect 8235 33823 8277 33832
rect 8139 4304 8181 4313
rect 8139 4264 8140 4304
rect 8180 4264 8181 4304
rect 8139 4255 8181 4264
rect 5163 4136 5205 4145
rect 5163 4096 5164 4136
rect 5204 4096 5205 4136
rect 5163 4087 5205 4096
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 4107 3716 4149 3725
rect 4107 3676 4108 3716
rect 4148 3676 4149 3716
rect 4107 3667 4149 3676
rect 8236 3473 8276 33823
rect 8235 3464 8277 3473
rect 8235 3424 8236 3464
rect 8276 3424 8277 3464
rect 8235 3415 8277 3424
rect 747 3380 789 3389
rect 747 3340 748 3380
rect 788 3340 789 3380
rect 747 3331 789 3340
rect 651 3128 693 3137
rect 651 3088 652 3128
rect 692 3088 693 3128
rect 651 3079 693 3088
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 8332 2885 8372 33907
rect 10348 33797 10388 34252
rect 10444 34049 10484 34924
rect 10636 34889 10676 35083
rect 12940 34964 12980 34973
rect 10635 34880 10677 34889
rect 10635 34840 10636 34880
rect 10676 34840 10677 34880
rect 10635 34831 10677 34840
rect 12940 34553 12980 34924
rect 13228 34628 13268 35176
rect 13324 35216 13364 35225
rect 13611 35216 13653 35225
rect 13364 35176 13556 35216
rect 13324 35167 13364 35176
rect 13228 34588 13364 34628
rect 10636 34544 10676 34553
rect 12075 34544 12117 34553
rect 10676 34504 10868 34544
rect 10636 34495 10676 34504
rect 10828 34376 10868 34504
rect 12075 34504 12076 34544
rect 12116 34504 12117 34544
rect 12075 34495 12117 34504
rect 12939 34544 12981 34553
rect 12939 34504 12940 34544
rect 12980 34504 12981 34544
rect 12939 34495 12981 34504
rect 10828 34327 10868 34336
rect 11212 34376 11252 34385
rect 11212 34133 11252 34336
rect 12076 34376 12116 34495
rect 12076 34327 12116 34336
rect 13324 34217 13364 34588
rect 13419 34544 13461 34553
rect 13419 34504 13420 34544
rect 13460 34504 13461 34544
rect 13419 34495 13461 34504
rect 13420 34376 13460 34495
rect 13420 34327 13460 34336
rect 13228 34208 13268 34217
rect 11211 34124 11253 34133
rect 11211 34084 11212 34124
rect 11252 34084 11253 34124
rect 11211 34075 11253 34084
rect 13228 34049 13268 34168
rect 13323 34208 13365 34217
rect 13323 34168 13324 34208
rect 13364 34168 13365 34208
rect 13323 34159 13365 34168
rect 13516 34049 13556 35176
rect 13611 35176 13612 35216
rect 13652 35176 13653 35216
rect 13611 35167 13653 35176
rect 13612 35082 13652 35167
rect 13804 34376 13844 35671
rect 13804 34327 13844 34336
rect 10443 34040 10485 34049
rect 10443 34000 10444 34040
rect 10484 34000 10485 34040
rect 10443 33991 10485 34000
rect 13227 34040 13269 34049
rect 13227 34000 13228 34040
rect 13268 34000 13269 34040
rect 13227 33991 13269 34000
rect 13515 34040 13557 34049
rect 13515 34000 13516 34040
rect 13556 34000 13557 34040
rect 13515 33991 13557 34000
rect 13228 33797 13268 33991
rect 10347 33788 10389 33797
rect 10347 33748 10348 33788
rect 10388 33748 10389 33788
rect 10347 33739 10389 33748
rect 13227 33788 13269 33797
rect 13227 33748 13228 33788
rect 13268 33748 13269 33788
rect 13227 33739 13269 33748
rect 13900 32117 13940 35932
rect 16876 36056 16916 36065
rect 14187 35888 14229 35897
rect 14187 35848 14188 35888
rect 14228 35848 14229 35888
rect 14187 35839 14229 35848
rect 16203 35888 16245 35897
rect 16203 35848 16204 35888
rect 16244 35848 16245 35888
rect 16203 35839 16245 35848
rect 16492 35888 16532 35897
rect 14091 35720 14133 35729
rect 14091 35680 14092 35720
rect 14132 35680 14133 35720
rect 14091 35671 14133 35680
rect 14092 35586 14132 35671
rect 14091 35216 14133 35225
rect 14188 35216 14228 35839
rect 16204 35754 16244 35839
rect 15339 35720 15381 35729
rect 15339 35680 15340 35720
rect 15380 35680 15381 35720
rect 15339 35671 15381 35680
rect 14091 35176 14092 35216
rect 14132 35176 14228 35216
rect 14380 35216 14420 35225
rect 14091 35167 14133 35176
rect 14092 35082 14132 35167
rect 14380 34217 14420 35176
rect 14476 35216 14516 35225
rect 14476 35057 14516 35176
rect 14667 35216 14709 35225
rect 14667 35176 14668 35216
rect 14708 35176 14709 35216
rect 14667 35167 14709 35176
rect 14956 35216 14996 35225
rect 14475 35048 14517 35057
rect 14475 35008 14476 35048
rect 14516 35008 14517 35048
rect 14475 34999 14517 35008
rect 14668 34376 14708 35167
rect 14764 35048 14804 35057
rect 14956 35048 14996 35176
rect 14804 35008 14996 35048
rect 15340 35216 15380 35671
rect 14764 34999 14804 35008
rect 15340 34973 15380 35176
rect 16203 35216 16245 35225
rect 16203 35176 16204 35216
rect 16244 35176 16245 35216
rect 16203 35167 16245 35176
rect 16204 35082 16244 35167
rect 15339 34964 15381 34973
rect 15339 34924 15340 34964
rect 15380 34924 15381 34964
rect 15339 34915 15381 34924
rect 14668 34327 14708 34336
rect 14379 34208 14421 34217
rect 14379 34168 14380 34208
rect 14420 34168 14421 34208
rect 14379 34159 14421 34168
rect 15819 34208 15861 34217
rect 15819 34168 15820 34208
rect 15860 34168 15861 34208
rect 15819 34159 15861 34168
rect 15820 33797 15860 34159
rect 16011 34040 16053 34049
rect 16011 34000 16012 34040
rect 16052 34000 16053 34040
rect 16011 33991 16053 34000
rect 15819 33788 15861 33797
rect 15819 33748 15820 33788
rect 15860 33748 15861 33788
rect 15819 33739 15861 33748
rect 16012 33713 16052 33991
rect 16011 33704 16053 33713
rect 16011 33664 16012 33704
rect 16052 33664 16053 33704
rect 16011 33655 16053 33664
rect 13899 32108 13941 32117
rect 13899 32068 13900 32108
rect 13940 32068 13941 32108
rect 13899 32059 13941 32068
rect 15160 31604 15202 31613
rect 15160 31564 15161 31604
rect 15201 31564 15202 31604
rect 15160 31555 15202 31564
rect 15161 31374 15201 31555
rect 16492 31529 16532 35848
rect 16588 35804 16628 35813
rect 16588 34637 16628 35764
rect 16587 34628 16629 34637
rect 16587 34588 16588 34628
rect 16628 34588 16629 34628
rect 16587 34579 16629 34588
rect 16876 34376 16916 36016
rect 18507 35888 18549 35897
rect 18507 35848 18508 35888
rect 18548 35848 18549 35888
rect 18507 35839 18549 35848
rect 18796 35888 18836 35897
rect 17547 35804 17589 35813
rect 17547 35764 17548 35804
rect 17588 35764 17589 35804
rect 17547 35755 17589 35764
rect 17548 35384 17588 35755
rect 18508 35754 18548 35839
rect 18796 35729 18836 35848
rect 18891 35804 18933 35813
rect 18891 35764 18892 35804
rect 18932 35764 18933 35804
rect 18891 35755 18933 35764
rect 18795 35720 18837 35729
rect 18795 35680 18796 35720
rect 18836 35680 18837 35720
rect 18795 35671 18837 35680
rect 18892 35670 18932 35755
rect 17548 35335 17588 35344
rect 18123 35216 18165 35225
rect 18123 35176 18124 35216
rect 18164 35176 18165 35216
rect 18123 35167 18165 35176
rect 18699 35216 18741 35225
rect 18699 35176 18700 35216
rect 18740 35176 18741 35216
rect 18699 35167 18741 35176
rect 17451 35132 17493 35141
rect 17451 35092 17452 35132
rect 17492 35092 17493 35132
rect 17451 35083 17493 35092
rect 17259 35048 17301 35057
rect 17259 35008 17260 35048
rect 17300 35008 17396 35048
rect 17259 34999 17301 35008
rect 17260 34980 17300 34999
rect 17356 34964 17396 35008
rect 17356 34805 17396 34924
rect 17355 34796 17397 34805
rect 17355 34756 17356 34796
rect 17396 34756 17397 34796
rect 17355 34747 17397 34756
rect 17452 34628 17492 35083
rect 16876 34327 16916 34336
rect 17308 34588 17492 34628
rect 17548 34964 17588 34973
rect 17308 34376 17348 34588
rect 17308 34327 17348 34336
rect 17548 31697 17588 34924
rect 18027 34796 18069 34805
rect 18027 34756 18028 34796
rect 18068 34756 18069 34796
rect 18027 34747 18069 34756
rect 18028 31772 18068 34747
rect 18124 34376 18164 35167
rect 18700 35082 18740 35167
rect 18988 35141 19028 36688
rect 19084 36679 19124 36688
rect 19948 36728 19988 36737
rect 19988 36688 20180 36728
rect 19948 36679 19988 36688
rect 19180 36056 19220 36065
rect 19083 35888 19125 35897
rect 19083 35848 19084 35888
rect 19124 35848 19125 35888
rect 19083 35839 19125 35848
rect 18987 35132 19029 35141
rect 18987 35092 18988 35132
rect 19028 35092 19029 35132
rect 18987 35083 19029 35092
rect 19084 35057 19124 35839
rect 19180 35720 19220 36016
rect 19660 35897 19700 35982
rect 19948 35897 19988 35982
rect 19659 35888 19701 35897
rect 19659 35848 19660 35888
rect 19700 35848 19701 35888
rect 19659 35839 19701 35848
rect 19947 35888 19989 35897
rect 19947 35848 19948 35888
rect 19988 35848 19989 35888
rect 19947 35839 19989 35848
rect 20044 35804 20084 35813
rect 20044 35729 20084 35764
rect 20043 35720 20085 35729
rect 19180 35680 19988 35720
rect 19275 35552 19317 35561
rect 19275 35512 19276 35552
rect 19316 35512 19317 35552
rect 19275 35503 19317 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 19083 35048 19125 35057
rect 19083 35008 19084 35048
rect 19124 35008 19125 35048
rect 19083 34999 19125 35008
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 19276 34637 19316 35503
rect 19948 35300 19988 35680
rect 20043 35680 20044 35720
rect 20084 35680 20085 35720
rect 20043 35671 20085 35680
rect 19948 35251 19988 35260
rect 19564 35216 19604 35227
rect 19564 35141 19604 35176
rect 19563 35132 19605 35141
rect 19563 35092 19564 35132
rect 19604 35092 19605 35132
rect 19563 35083 19605 35092
rect 20044 34973 20084 35671
rect 20140 35225 20180 36688
rect 20139 35216 20181 35225
rect 20139 35176 20140 35216
rect 20180 35176 20181 35216
rect 20139 35167 20181 35176
rect 20236 35132 20276 36772
rect 20523 36728 20565 36737
rect 20523 36688 20524 36728
rect 20564 36688 20565 36728
rect 20523 36679 20565 36688
rect 20524 36140 20564 36679
rect 20524 36091 20564 36100
rect 20332 36056 20372 36065
rect 20332 35636 20372 36016
rect 20620 35897 20660 37360
rect 20716 37400 20756 37409
rect 21003 37400 21045 37409
rect 20756 37360 20948 37400
rect 20716 37351 20756 37360
rect 20908 36980 20948 37360
rect 21003 37360 21004 37400
rect 21044 37360 21045 37400
rect 21003 37351 21045 37360
rect 21388 37400 21428 37409
rect 21771 37400 21813 37409
rect 21428 37360 21620 37400
rect 21388 37351 21428 37360
rect 21004 37266 21044 37351
rect 20812 36940 21140 36980
rect 20619 35888 20661 35897
rect 20619 35848 20620 35888
rect 20660 35848 20661 35888
rect 20619 35839 20661 35848
rect 20812 35888 20852 36940
rect 21100 36896 21140 36940
rect 21140 36856 21524 36896
rect 21100 36847 21140 36856
rect 21388 36728 21428 36737
rect 21388 36569 21428 36688
rect 21387 36560 21429 36569
rect 21387 36520 21388 36560
rect 21428 36520 21429 36560
rect 21387 36511 21429 36520
rect 21292 36476 21332 36485
rect 20812 35839 20852 35848
rect 20907 35888 20949 35897
rect 21196 35888 21236 35897
rect 20907 35848 20908 35888
rect 20948 35848 21196 35888
rect 20907 35839 20949 35848
rect 21196 35839 21236 35848
rect 20332 35596 20756 35636
rect 20716 35300 20756 35596
rect 20908 35393 20948 35839
rect 21004 35720 21044 35725
rect 21292 35720 21332 36436
rect 21484 35888 21524 36856
rect 21484 35839 21524 35848
rect 21004 35716 21332 35720
rect 21044 35680 21332 35716
rect 21388 35720 21428 35729
rect 21004 35667 21044 35676
rect 20907 35384 20949 35393
rect 20907 35344 20908 35384
rect 20948 35344 20949 35384
rect 20907 35335 20949 35344
rect 21099 35384 21141 35393
rect 21099 35344 21100 35384
rect 21140 35344 21141 35384
rect 21099 35335 21141 35344
rect 20716 35251 20756 35260
rect 20523 35216 20565 35225
rect 20523 35176 20524 35216
rect 20564 35176 20565 35216
rect 20523 35167 20565 35176
rect 21100 35216 21140 35335
rect 20332 35132 20372 35141
rect 20236 35092 20332 35132
rect 20139 35048 20181 35057
rect 20139 35008 20140 35048
rect 20180 35008 20181 35048
rect 20139 34999 20181 35008
rect 20043 34964 20085 34973
rect 20043 34924 20044 34964
rect 20084 34924 20085 34964
rect 20043 34915 20085 34924
rect 20140 34914 20180 34999
rect 20332 34889 20372 35092
rect 20331 34880 20373 34889
rect 20331 34840 20332 34880
rect 20372 34840 20373 34880
rect 20331 34831 20373 34840
rect 19275 34628 19317 34637
rect 19275 34588 19276 34628
rect 19316 34588 19317 34628
rect 19275 34579 19317 34588
rect 19276 34494 19316 34579
rect 19563 34460 19605 34469
rect 19563 34420 19564 34460
rect 19604 34420 19605 34460
rect 19563 34411 19605 34420
rect 18124 34327 18164 34336
rect 19564 34376 19604 34411
rect 19564 34325 19604 34336
rect 20524 34376 20564 35167
rect 21100 35141 21140 35176
rect 21099 35132 21141 35141
rect 21099 35092 21100 35132
rect 21140 35092 21141 35132
rect 21099 35083 21141 35092
rect 21100 35052 21140 35083
rect 21388 35057 21428 35680
rect 21580 35393 21620 37360
rect 21771 37360 21772 37400
rect 21812 37360 21813 37400
rect 21771 37351 21813 37360
rect 21868 36737 21908 38368
rect 22060 38359 22100 38368
rect 26572 38408 26612 38417
rect 27532 38408 27572 38417
rect 26612 38368 26900 38408
rect 26572 38359 26612 38368
rect 21964 38240 22004 38249
rect 25996 38240 26036 38249
rect 21964 37460 22004 38200
rect 25900 38200 25996 38240
rect 22732 38156 22772 38165
rect 22540 37988 22580 37997
rect 22540 37460 22580 37948
rect 21964 37420 22100 37460
rect 21867 36728 21909 36737
rect 21867 36688 21868 36728
rect 21908 36688 21909 36728
rect 21867 36679 21909 36688
rect 21675 36560 21717 36569
rect 21675 36520 21676 36560
rect 21716 36520 21717 36560
rect 21675 36511 21717 36520
rect 21676 35888 21716 36511
rect 21771 36224 21813 36233
rect 21771 36184 21772 36224
rect 21812 36184 21813 36224
rect 21771 36175 21813 36184
rect 21676 35839 21716 35848
rect 21772 35888 21812 36175
rect 21868 36140 21908 36679
rect 22060 36560 22100 37420
rect 22444 37420 22580 37460
rect 22251 37400 22293 37409
rect 22251 37360 22252 37400
rect 22292 37360 22293 37400
rect 22251 37351 22293 37360
rect 22252 37266 22292 37351
rect 22347 37232 22389 37241
rect 22347 37192 22348 37232
rect 22388 37192 22389 37232
rect 22347 37183 22389 37192
rect 22348 36728 22388 37183
rect 22060 36511 22100 36520
rect 22156 36688 22348 36728
rect 21964 36140 22004 36149
rect 21868 36100 21964 36140
rect 21964 36091 22004 36100
rect 21772 35839 21812 35848
rect 21964 35888 22004 35897
rect 22156 35888 22196 36688
rect 22348 36679 22388 36688
rect 22444 36728 22484 37420
rect 22539 37316 22581 37325
rect 22539 37276 22540 37316
rect 22580 37276 22581 37316
rect 22539 37267 22581 37276
rect 22444 36653 22484 36688
rect 22540 36954 22580 37267
rect 22443 36644 22485 36653
rect 22443 36604 22444 36644
rect 22484 36604 22485 36644
rect 22443 36595 22485 36604
rect 22444 36233 22484 36595
rect 22540 36569 22580 36914
rect 22539 36560 22581 36569
rect 22539 36520 22540 36560
rect 22580 36520 22581 36560
rect 22539 36511 22581 36520
rect 22443 36224 22485 36233
rect 22443 36184 22444 36224
rect 22484 36184 22485 36224
rect 22443 36175 22485 36184
rect 22004 35848 22196 35888
rect 22252 35888 22292 35897
rect 22444 35888 22484 36175
rect 22292 35848 22484 35888
rect 22540 35888 22580 35897
rect 21964 35839 22004 35848
rect 22252 35839 22292 35848
rect 21579 35384 21621 35393
rect 21579 35344 21580 35384
rect 21620 35344 21621 35384
rect 21579 35335 21621 35344
rect 21963 35216 22005 35225
rect 21963 35176 21964 35216
rect 22004 35176 22005 35216
rect 21963 35167 22005 35176
rect 21964 35082 22004 35167
rect 21387 35048 21429 35057
rect 21387 35008 21388 35048
rect 21428 35008 21429 35048
rect 21387 34999 21429 35008
rect 22540 34469 22580 35848
rect 22635 35804 22677 35813
rect 22635 35764 22636 35804
rect 22676 35764 22677 35804
rect 22635 35755 22677 35764
rect 22636 35670 22676 35755
rect 22732 35057 22772 38116
rect 23692 38156 23732 38165
rect 23596 37316 23636 37325
rect 23500 37276 23596 37316
rect 23403 37232 23445 37241
rect 23403 37192 23404 37232
rect 23444 37192 23445 37232
rect 23403 37183 23445 37192
rect 23404 37098 23444 37183
rect 23115 37064 23157 37073
rect 23115 37024 23116 37064
rect 23156 37024 23157 37064
rect 23115 37015 23157 37024
rect 23019 36728 23061 36737
rect 23019 36688 23020 36728
rect 23060 36688 23061 36728
rect 23019 36679 23061 36688
rect 23116 36728 23156 37015
rect 23404 36896 23444 36905
rect 23500 36896 23540 37276
rect 23596 37267 23636 37276
rect 23444 36856 23540 36896
rect 23404 36847 23444 36856
rect 23692 36821 23732 38116
rect 24268 38156 24308 38165
rect 24268 38072 24308 38116
rect 24652 38156 24692 38165
rect 24460 38072 24500 38081
rect 24268 38032 24460 38072
rect 23883 37988 23925 37997
rect 23883 37948 23884 37988
rect 23924 37948 23925 37988
rect 23883 37939 23925 37948
rect 24076 37988 24116 37997
rect 23884 37854 23924 37939
rect 23980 37400 24020 37409
rect 24076 37400 24116 37948
rect 24460 37577 24500 38032
rect 24652 37997 24692 38116
rect 24651 37988 24693 37997
rect 24651 37948 24652 37988
rect 24692 37948 24693 37988
rect 24651 37939 24693 37948
rect 24459 37568 24501 37577
rect 24459 37528 24460 37568
rect 24500 37528 24501 37568
rect 24459 37519 24501 37528
rect 24020 37360 24116 37400
rect 23980 37351 24020 37360
rect 24076 37157 24116 37360
rect 24555 37400 24597 37409
rect 24555 37360 24556 37400
rect 24596 37360 24597 37400
rect 24555 37351 24597 37360
rect 24843 37400 24885 37409
rect 24843 37360 24844 37400
rect 24884 37360 24885 37400
rect 24843 37351 24885 37360
rect 24171 37232 24213 37241
rect 24171 37192 24172 37232
rect 24212 37192 24213 37232
rect 24171 37183 24213 37192
rect 23787 37148 23829 37157
rect 23787 37108 23788 37148
rect 23828 37108 23829 37148
rect 23787 37099 23829 37108
rect 24075 37148 24117 37157
rect 24075 37108 24076 37148
rect 24116 37108 24117 37148
rect 24075 37099 24117 37108
rect 23691 36812 23733 36821
rect 23691 36772 23692 36812
rect 23732 36772 23733 36812
rect 23691 36763 23733 36772
rect 23116 36679 23156 36688
rect 23020 36594 23060 36679
rect 23307 36476 23349 36485
rect 23307 36436 23308 36476
rect 23348 36436 23349 36476
rect 23307 36427 23349 36436
rect 22924 36056 22964 36065
rect 22731 35048 22773 35057
rect 22731 35008 22732 35048
rect 22772 35008 22773 35048
rect 22731 34999 22773 35008
rect 21291 34460 21333 34469
rect 21291 34420 21292 34460
rect 21332 34420 21333 34460
rect 21291 34411 21333 34420
rect 22539 34460 22581 34469
rect 22539 34420 22540 34460
rect 22580 34420 22581 34460
rect 22539 34411 22581 34420
rect 20524 34327 20564 34336
rect 21004 34376 21044 34387
rect 21004 34301 21044 34336
rect 21292 34376 21332 34411
rect 21292 34325 21332 34336
rect 22251 34376 22293 34385
rect 22251 34336 22252 34376
rect 22292 34336 22293 34376
rect 22924 34376 22964 36016
rect 23308 35888 23348 36427
rect 23692 35888 23732 35897
rect 23788 35888 23828 37099
rect 23979 37064 24021 37073
rect 23979 37024 23980 37064
rect 24020 37024 24021 37064
rect 23979 37015 24021 37024
rect 23884 36728 23924 36739
rect 23884 36653 23924 36688
rect 23980 36728 24020 37015
rect 24172 36905 24212 37183
rect 24459 36980 24501 36989
rect 24459 36940 24460 36980
rect 24500 36940 24501 36980
rect 24459 36931 24501 36940
rect 24171 36896 24213 36905
rect 24171 36856 24172 36896
rect 24212 36856 24213 36896
rect 24171 36847 24213 36856
rect 23980 36679 24020 36688
rect 24172 36728 24212 36847
rect 24172 36679 24212 36688
rect 24364 36728 24404 36737
rect 23883 36644 23925 36653
rect 23883 36604 23884 36644
rect 23924 36604 23925 36644
rect 23883 36595 23925 36604
rect 24172 36560 24212 36569
rect 24364 36560 24404 36688
rect 24460 36728 24500 36931
rect 24460 36679 24500 36688
rect 24212 36520 24404 36560
rect 24172 36511 24212 36520
rect 24556 35888 24596 37351
rect 24844 37266 24884 37351
rect 25611 37064 25653 37073
rect 25611 37024 25612 37064
rect 25652 37024 25653 37064
rect 25611 37015 25653 37024
rect 24843 36896 24885 36905
rect 24843 36856 24844 36896
rect 24884 36856 24885 36896
rect 24843 36847 24885 36856
rect 25131 36896 25173 36905
rect 25131 36856 25132 36896
rect 25172 36856 25173 36896
rect 25131 36847 25173 36856
rect 25515 36896 25557 36905
rect 25515 36856 25516 36896
rect 25556 36856 25557 36896
rect 25515 36847 25557 36856
rect 25612 36896 25652 37015
rect 25900 36896 25940 38200
rect 25996 38191 26036 38200
rect 26476 38240 26516 38249
rect 26668 38240 26708 38249
rect 26516 38200 26612 38240
rect 26476 38191 26516 38200
rect 26092 37988 26132 37997
rect 25996 37232 26036 37241
rect 25996 37073 26036 37192
rect 25995 37064 26037 37073
rect 25995 37024 25996 37064
rect 26036 37024 26037 37064
rect 25995 37015 26037 37024
rect 25612 36847 25652 36856
rect 25708 36856 25940 36896
rect 24651 36812 24693 36821
rect 24651 36772 24652 36812
rect 24692 36772 24693 36812
rect 24651 36763 24693 36772
rect 24652 36728 24692 36763
rect 24844 36762 24884 36847
rect 25132 36762 25172 36847
rect 25323 36812 25365 36821
rect 25323 36772 25324 36812
rect 25364 36772 25365 36812
rect 25323 36763 25365 36772
rect 24652 36677 24692 36688
rect 24939 36728 24981 36737
rect 24939 36688 24940 36728
rect 24980 36688 24981 36728
rect 24939 36679 24981 36688
rect 24940 36594 24980 36679
rect 25324 36678 25364 36763
rect 25516 36728 25556 36847
rect 25516 36679 25556 36688
rect 25612 36728 25652 36739
rect 25708 36737 25748 36856
rect 25612 36653 25652 36688
rect 25707 36728 25749 36737
rect 25707 36688 25708 36728
rect 25748 36688 25749 36728
rect 25707 36679 25749 36688
rect 25611 36644 25653 36653
rect 25611 36604 25612 36644
rect 25652 36604 25653 36644
rect 25611 36595 25653 36604
rect 24651 36476 24693 36485
rect 24651 36436 24652 36476
rect 24692 36436 24693 36476
rect 24651 36427 24693 36436
rect 24652 36342 24692 36427
rect 25708 36140 25748 36679
rect 25996 36653 26036 37015
rect 26092 36989 26132 37948
rect 26572 37652 26612 38200
rect 26668 37829 26708 38200
rect 26667 37820 26709 37829
rect 26667 37780 26668 37820
rect 26708 37780 26709 37820
rect 26667 37771 26709 37780
rect 26668 37652 26708 37661
rect 26572 37612 26668 37652
rect 26668 37603 26708 37612
rect 26380 37400 26420 37409
rect 26091 36980 26133 36989
rect 26091 36940 26092 36980
rect 26132 36940 26133 36980
rect 26091 36931 26133 36940
rect 26380 36821 26420 37360
rect 26476 37400 26516 37409
rect 26284 36812 26324 36821
rect 26092 36772 26284 36812
rect 25995 36644 26037 36653
rect 25995 36604 25996 36644
rect 26036 36604 26037 36644
rect 25995 36595 26037 36604
rect 25708 36091 25748 36100
rect 23308 35839 23348 35848
rect 23500 35848 23692 35888
rect 23732 35848 23828 35888
rect 24460 35848 24556 35888
rect 23115 34964 23157 34973
rect 23115 34924 23116 34964
rect 23156 34924 23157 34964
rect 23115 34915 23157 34924
rect 23116 34830 23156 34915
rect 23116 34376 23156 34385
rect 22924 34336 23116 34376
rect 22251 34327 22293 34336
rect 23116 34327 23156 34336
rect 23500 34376 23540 35848
rect 23692 35839 23732 35848
rect 23787 34964 23829 34973
rect 23787 34924 23788 34964
rect 23828 34924 23829 34964
rect 23787 34915 23829 34924
rect 23500 34327 23540 34336
rect 21003 34292 21045 34301
rect 21003 34252 21004 34292
rect 21044 34252 21045 34292
rect 21003 34243 21045 34252
rect 22252 34242 22292 34327
rect 18795 34208 18837 34217
rect 18795 34168 18796 34208
rect 18836 34168 18837 34208
rect 18795 34159 18837 34168
rect 19276 34208 19316 34217
rect 18796 31772 18836 34159
rect 19276 31772 19316 34168
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 23788 31772 23828 34915
rect 24363 34376 24405 34385
rect 24460 34376 24500 35848
rect 24556 35839 24596 35848
rect 25035 35888 25077 35897
rect 25035 35848 25036 35888
rect 25076 35848 25077 35888
rect 25035 35839 25077 35848
rect 25036 35216 25076 35839
rect 26092 35300 26132 36772
rect 26284 36763 26324 36772
rect 26379 36812 26421 36821
rect 26379 36772 26380 36812
rect 26420 36772 26421 36812
rect 26379 36763 26421 36772
rect 26380 36728 26420 36763
rect 26476 36728 26516 37360
rect 26668 37400 26708 37409
rect 26668 37157 26708 37360
rect 26860 37400 26900 38368
rect 27436 38368 27532 38408
rect 26860 37351 26900 37360
rect 27244 37400 27284 37409
rect 26667 37148 26709 37157
rect 26667 37108 26668 37148
rect 26708 37108 26709 37148
rect 26667 37099 26709 37108
rect 27244 37073 27284 37360
rect 27436 37157 27476 38368
rect 27532 38359 27572 38368
rect 33196 38368 33716 38408
rect 27628 38324 27668 38333
rect 27532 37988 27572 37997
rect 27532 37325 27572 37948
rect 27531 37316 27573 37325
rect 27531 37276 27532 37316
rect 27572 37276 27573 37316
rect 27531 37267 27573 37276
rect 27628 37241 27668 38284
rect 29452 38324 29492 38333
rect 29492 38284 29684 38324
rect 29452 38275 29492 38284
rect 27724 38240 27764 38249
rect 27724 37988 27764 38200
rect 27820 38240 27860 38249
rect 28972 38240 29012 38249
rect 27860 38200 27956 38240
rect 27820 38191 27860 38200
rect 27724 37948 27860 37988
rect 27723 37820 27765 37829
rect 27723 37780 27724 37820
rect 27764 37780 27765 37820
rect 27723 37771 27765 37780
rect 27627 37232 27669 37241
rect 27627 37192 27628 37232
rect 27668 37192 27669 37232
rect 27627 37183 27669 37192
rect 27435 37148 27477 37157
rect 27435 37108 27436 37148
rect 27476 37108 27477 37148
rect 27435 37099 27477 37108
rect 26859 37064 26901 37073
rect 26859 37024 26860 37064
rect 26900 37024 26901 37064
rect 26859 37015 26901 37024
rect 27243 37064 27285 37073
rect 27243 37024 27244 37064
rect 27284 37024 27285 37064
rect 27243 37015 27285 37024
rect 26764 36728 26804 36737
rect 26476 36688 26764 36728
rect 26380 36678 26420 36688
rect 26475 36308 26517 36317
rect 26475 36268 26476 36308
rect 26516 36268 26517 36308
rect 26475 36259 26517 36268
rect 26092 35251 26132 35260
rect 26188 35804 26228 35813
rect 25036 34637 25076 35176
rect 25228 34964 25268 34973
rect 25035 34628 25077 34637
rect 25035 34588 25036 34628
rect 25076 34588 25077 34628
rect 25035 34579 25077 34588
rect 24363 34336 24364 34376
rect 24404 34336 24500 34376
rect 24363 34327 24405 34336
rect 24364 34242 24404 34327
rect 25228 33965 25268 34924
rect 25516 34460 25556 34471
rect 25516 34385 25556 34420
rect 25515 34376 25557 34385
rect 25515 34336 25516 34376
rect 25556 34336 25557 34376
rect 25515 34327 25557 34336
rect 25227 33956 25269 33965
rect 25227 33916 25228 33956
rect 25268 33916 25269 33956
rect 25227 33907 25269 33916
rect 26188 33881 26228 35764
rect 26476 35216 26516 36259
rect 26764 36233 26804 36688
rect 26860 36317 26900 37015
rect 27339 36980 27381 36989
rect 27339 36940 27340 36980
rect 27380 36940 27381 36980
rect 27339 36931 27381 36940
rect 27243 36812 27285 36821
rect 27243 36772 27244 36812
rect 27284 36772 27285 36812
rect 27243 36763 27285 36772
rect 27148 36728 27188 36739
rect 27148 36653 27188 36688
rect 27244 36728 27284 36763
rect 27244 36677 27284 36688
rect 27340 36728 27380 36931
rect 27340 36679 27380 36688
rect 27436 36728 27476 36737
rect 27147 36644 27189 36653
rect 27147 36604 27148 36644
rect 27188 36604 27189 36644
rect 27147 36595 27189 36604
rect 27436 36569 27476 36688
rect 27531 36644 27573 36653
rect 27531 36604 27532 36644
rect 27572 36604 27573 36644
rect 27531 36595 27573 36604
rect 27435 36560 27477 36569
rect 27435 36520 27436 36560
rect 27476 36520 27477 36560
rect 27435 36511 27477 36520
rect 26859 36308 26901 36317
rect 26859 36268 26860 36308
rect 26900 36268 26901 36308
rect 26859 36259 26901 36268
rect 26763 36224 26805 36233
rect 26763 36184 26764 36224
rect 26804 36184 26805 36224
rect 26763 36175 26805 36184
rect 27099 35888 27141 35897
rect 27099 35848 27100 35888
rect 27140 35848 27141 35888
rect 27099 35839 27141 35848
rect 27532 35888 27572 36595
rect 27628 36560 27668 36569
rect 27724 36560 27764 37771
rect 27820 36989 27860 37948
rect 27819 36980 27861 36989
rect 27819 36940 27820 36980
rect 27860 36940 27861 36980
rect 27819 36931 27861 36940
rect 27668 36520 27764 36560
rect 27819 36560 27861 36569
rect 27819 36520 27820 36560
rect 27860 36520 27861 36560
rect 27628 36511 27668 36520
rect 27819 36511 27861 36520
rect 27820 36426 27860 36511
rect 27723 36224 27765 36233
rect 27723 36184 27724 36224
rect 27764 36184 27765 36224
rect 27723 36175 27765 36184
rect 27532 35839 27572 35848
rect 27724 35888 27764 36175
rect 27820 36056 27860 36065
rect 27916 36056 27956 38200
rect 28972 37409 29012 38200
rect 29259 38240 29301 38249
rect 29259 38200 29260 38240
rect 29300 38200 29301 38240
rect 29259 38191 29301 38200
rect 29260 37829 29300 38191
rect 29259 37820 29301 37829
rect 29259 37780 29260 37820
rect 29300 37780 29301 37820
rect 29259 37771 29301 37780
rect 28107 37400 28149 37409
rect 28107 37360 28108 37400
rect 28148 37360 28149 37400
rect 28107 37351 28149 37360
rect 28971 37400 29013 37409
rect 28971 37360 28972 37400
rect 29012 37360 29013 37400
rect 28971 37351 29013 37360
rect 28108 37266 28148 37351
rect 28011 37148 28053 37157
rect 28011 37108 28012 37148
rect 28052 37108 28053 37148
rect 28011 37099 28053 37108
rect 28012 36737 28052 37099
rect 28203 37064 28245 37073
rect 28203 37024 28204 37064
rect 28244 37024 28245 37064
rect 28203 37015 28245 37024
rect 28108 36896 28148 36905
rect 28011 36728 28053 36737
rect 28011 36688 28012 36728
rect 28052 36688 28053 36728
rect 28011 36679 28053 36688
rect 28012 36594 28052 36679
rect 28011 36476 28053 36485
rect 28011 36436 28012 36476
rect 28052 36436 28053 36476
rect 28011 36427 28053 36436
rect 27860 36016 27956 36056
rect 27820 36007 27860 36016
rect 27724 35839 27764 35848
rect 27820 35888 27860 35897
rect 28012 35888 28052 36427
rect 28108 36233 28148 36856
rect 28107 36224 28149 36233
rect 28107 36184 28108 36224
rect 28148 36184 28149 36224
rect 28107 36175 28149 36184
rect 27860 35848 28052 35888
rect 27820 35839 27860 35848
rect 27100 35754 27140 35839
rect 28204 35804 28244 37015
rect 28972 36485 29012 37351
rect 29260 37232 29300 37241
rect 29260 36737 29300 37192
rect 29644 36812 29684 38284
rect 29739 38240 29781 38249
rect 29739 38200 29740 38240
rect 29780 38200 29781 38240
rect 29739 38191 29781 38200
rect 29932 38240 29972 38249
rect 29740 38106 29780 38191
rect 29836 37988 29876 37997
rect 29740 37400 29780 37409
rect 29740 37241 29780 37360
rect 29836 37400 29876 37948
rect 29932 37409 29972 38200
rect 30411 37568 30453 37577
rect 30411 37528 30412 37568
rect 30452 37528 30453 37568
rect 30411 37519 30453 37528
rect 32907 37568 32949 37577
rect 32907 37528 32908 37568
rect 32948 37528 32949 37568
rect 32907 37519 32949 37528
rect 29836 37351 29876 37360
rect 29931 37400 29973 37409
rect 29931 37360 29932 37400
rect 29972 37360 29973 37400
rect 29931 37351 29973 37360
rect 30220 37316 30260 37325
rect 29739 37232 29781 37241
rect 29739 37192 29740 37232
rect 29780 37192 29781 37232
rect 29739 37183 29781 37192
rect 30028 37232 30068 37241
rect 30220 37232 30260 37276
rect 30068 37192 30260 37232
rect 30028 37183 30068 37192
rect 30027 37064 30069 37073
rect 30027 37024 30028 37064
rect 30068 37024 30069 37064
rect 30027 37015 30069 37024
rect 29644 36763 29684 36772
rect 30028 36737 30068 37015
rect 29259 36728 29301 36737
rect 29259 36688 29260 36728
rect 29300 36688 29301 36728
rect 29259 36679 29301 36688
rect 30027 36728 30069 36737
rect 30027 36688 30028 36728
rect 30068 36688 30069 36728
rect 30027 36679 30069 36688
rect 30028 36594 30068 36679
rect 28971 36476 29013 36485
rect 28971 36436 28972 36476
rect 29012 36436 29013 36476
rect 28971 36427 29013 36436
rect 28491 36224 28533 36233
rect 28491 36184 28492 36224
rect 28532 36184 28533 36224
rect 28491 36175 28533 36184
rect 28012 35764 28244 35804
rect 26476 35167 26516 35176
rect 27340 35216 27380 35225
rect 26283 34880 26325 34889
rect 26283 34840 26284 34880
rect 26324 34840 26325 34880
rect 26283 34831 26325 34840
rect 26284 34460 26324 34831
rect 26475 34712 26517 34721
rect 26475 34672 26476 34712
rect 26516 34672 26517 34712
rect 26475 34663 26517 34672
rect 26763 34712 26805 34721
rect 26763 34672 26764 34712
rect 26804 34672 26805 34712
rect 26763 34663 26805 34672
rect 26476 34544 26516 34663
rect 26476 34495 26516 34504
rect 26284 34411 26324 34420
rect 26764 34376 26804 34663
rect 27340 34637 27380 35176
rect 27339 34628 27381 34637
rect 27339 34588 27340 34628
rect 27380 34588 27381 34628
rect 27339 34579 27381 34588
rect 27436 34544 27476 34553
rect 27476 34504 27668 34544
rect 27436 34495 27476 34504
rect 26764 34327 26804 34336
rect 27051 34376 27093 34385
rect 27051 34336 27052 34376
rect 27092 34336 27093 34376
rect 27051 34327 27093 34336
rect 27628 34376 27668 34504
rect 27628 34327 27668 34336
rect 28012 34376 28052 35764
rect 28492 35384 28532 36175
rect 28492 35335 28532 35344
rect 30028 35216 30068 35225
rect 28875 34628 28917 34637
rect 28875 34588 28876 34628
rect 28916 34588 28917 34628
rect 30028 34628 30068 35176
rect 30412 35216 30452 37519
rect 32908 37484 32948 37519
rect 30604 37400 30644 37409
rect 30604 36737 30644 37360
rect 30891 37400 30933 37409
rect 30891 37360 30892 37400
rect 30932 37360 30933 37400
rect 30891 37351 30933 37360
rect 31467 37400 31509 37409
rect 31467 37360 31468 37400
rect 31508 37360 31509 37400
rect 31467 37351 31509 37360
rect 30603 36728 30645 36737
rect 30603 36688 30604 36728
rect 30644 36688 30645 36728
rect 30603 36679 30645 36688
rect 30892 36728 30932 37351
rect 31468 37266 31508 37351
rect 32043 37316 32085 37325
rect 32043 37276 32044 37316
rect 32084 37276 32085 37316
rect 32043 37267 32085 37276
rect 32044 36896 32084 37267
rect 32619 37232 32661 37241
rect 32619 37192 32620 37232
rect 32660 37192 32661 37232
rect 32619 37183 32661 37192
rect 32620 37098 32660 37183
rect 32044 36847 32084 36856
rect 32716 36812 32756 36821
rect 32428 36772 32716 36812
rect 32428 36728 32468 36772
rect 32716 36763 32756 36772
rect 30892 36679 30932 36688
rect 32236 36688 32468 36728
rect 31563 36476 31605 36485
rect 31563 36436 31564 36476
rect 31604 36436 31605 36476
rect 31563 36427 31605 36436
rect 31564 35888 31604 36427
rect 31947 36224 31989 36233
rect 31947 36184 31948 36224
rect 31988 36184 31989 36224
rect 31947 36175 31989 36184
rect 31468 35848 31564 35888
rect 30412 35167 30452 35176
rect 31276 35216 31316 35225
rect 30891 34712 30933 34721
rect 30891 34672 30892 34712
rect 30932 34672 30933 34712
rect 30891 34663 30933 34672
rect 30220 34628 30260 34637
rect 30028 34588 30220 34628
rect 28875 34579 28917 34588
rect 30220 34579 30260 34588
rect 28012 34327 28052 34336
rect 28876 34376 28916 34579
rect 28876 34327 28916 34336
rect 29547 34376 29589 34385
rect 29547 34336 29548 34376
rect 29588 34336 29589 34376
rect 29547 34327 29589 34336
rect 30507 34376 30549 34385
rect 30507 34336 30508 34376
rect 30548 34336 30549 34376
rect 30507 34327 30549 34336
rect 30604 34376 30644 34387
rect 27052 34242 27092 34327
rect 27147 34292 27189 34301
rect 27147 34252 27148 34292
rect 27188 34252 27189 34292
rect 27147 34243 27189 34252
rect 27148 34158 27188 34243
rect 26187 33872 26229 33881
rect 26187 33832 26188 33872
rect 26228 33832 26229 33872
rect 26187 33823 26229 33832
rect 23979 33788 24021 33797
rect 23979 33748 23980 33788
rect 24020 33748 24021 33788
rect 23979 33739 24021 33748
rect 23980 31772 24020 33739
rect 29548 31772 29588 34327
rect 29739 34292 29781 34301
rect 29739 34252 29740 34292
rect 29780 34252 29781 34292
rect 29739 34243 29781 34252
rect 30027 34292 30069 34301
rect 30027 34252 30028 34292
rect 30068 34252 30069 34292
rect 30027 34243 30069 34252
rect 29740 31772 29780 34243
rect 30028 34208 30068 34243
rect 30508 34242 30548 34327
rect 30604 34301 30644 34336
rect 30892 34376 30932 34663
rect 31276 34637 31316 35176
rect 31275 34628 31317 34637
rect 31275 34588 31276 34628
rect 31316 34588 31317 34628
rect 31275 34579 31317 34588
rect 30892 34327 30932 34336
rect 31276 34376 31316 34385
rect 31468 34376 31508 35848
rect 31564 35839 31604 35848
rect 31852 35888 31892 35897
rect 31852 35141 31892 35848
rect 31948 35888 31988 36175
rect 32236 36140 32276 36688
rect 32524 36644 32564 36653
rect 32332 36485 32372 36570
rect 32331 36476 32373 36485
rect 32331 36436 32332 36476
rect 32372 36436 32373 36476
rect 32331 36427 32373 36436
rect 32524 36224 32564 36604
rect 32908 36569 32948 37444
rect 33099 37232 33141 37241
rect 33099 37192 33100 37232
rect 33140 37192 33141 37232
rect 33099 37183 33141 37192
rect 33196 37232 33236 38368
rect 33676 38324 33716 38368
rect 33676 38275 33716 38284
rect 33291 38240 33333 38249
rect 33291 38200 33292 38240
rect 33332 38200 33333 38240
rect 33291 38191 33333 38200
rect 33580 38240 33620 38249
rect 33292 38106 33332 38191
rect 33580 37988 33620 38200
rect 33867 38240 33909 38249
rect 33867 38200 33868 38240
rect 33908 38200 33909 38240
rect 37516 38240 37556 38249
rect 33867 38191 33909 38200
rect 37420 38198 37460 38207
rect 33580 37948 33812 37988
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 33292 37232 33332 37260
rect 33196 37192 33292 37232
rect 33100 36741 33140 37183
rect 33100 36692 33140 36701
rect 32907 36560 32949 36569
rect 32907 36520 32908 36560
rect 32948 36520 32949 36560
rect 32907 36511 32949 36520
rect 32524 36184 32756 36224
rect 32236 36091 32276 36100
rect 32523 36056 32565 36065
rect 32523 36016 32524 36056
rect 32564 36016 32565 36056
rect 32523 36007 32565 36016
rect 31948 35839 31988 35848
rect 32524 35888 32564 36007
rect 32524 35839 32564 35848
rect 31851 35132 31893 35141
rect 31851 35092 31852 35132
rect 31892 35092 31893 35132
rect 31851 35083 31893 35092
rect 32428 34964 32468 34973
rect 31948 34544 31988 34553
rect 31988 34504 32180 34544
rect 31948 34495 31988 34504
rect 31316 34336 31508 34376
rect 31563 34376 31605 34385
rect 31563 34336 31564 34376
rect 31604 34336 31605 34376
rect 31276 34327 31316 34336
rect 31563 34327 31605 34336
rect 32043 34376 32085 34385
rect 32043 34336 32044 34376
rect 32084 34336 32085 34376
rect 32043 34327 32085 34336
rect 32140 34376 32180 34504
rect 32428 34385 32468 34924
rect 32523 34880 32565 34889
rect 32523 34840 32524 34880
rect 32564 34840 32565 34880
rect 32523 34831 32565 34840
rect 32140 34327 32180 34336
rect 32427 34376 32469 34385
rect 32427 34336 32428 34376
rect 32468 34336 32469 34376
rect 32427 34327 32469 34336
rect 32524 34376 32564 34831
rect 32716 34721 32756 36184
rect 32811 35132 32853 35141
rect 32811 35092 32812 35132
rect 32852 35092 32853 35132
rect 32811 35083 32853 35092
rect 32715 34712 32757 34721
rect 32715 34672 32716 34712
rect 32756 34672 32757 34712
rect 32715 34663 32757 34672
rect 32524 34327 32564 34336
rect 30603 34292 30645 34301
rect 30603 34252 30604 34292
rect 30644 34252 30645 34292
rect 30603 34243 30645 34252
rect 31564 34242 31604 34327
rect 31660 34292 31700 34303
rect 31660 34217 31700 34252
rect 30028 34157 30068 34168
rect 31659 34208 31701 34217
rect 31659 34168 31660 34208
rect 31700 34168 31701 34208
rect 31659 34159 31701 34168
rect 30219 34124 30261 34133
rect 30219 34084 30220 34124
rect 30260 34084 30261 34124
rect 30219 34075 30261 34084
rect 30220 31772 30260 34075
rect 31660 31772 31700 34159
rect 18028 31732 18081 31772
rect 18796 31732 18849 31772
rect 19276 31732 19617 31772
rect 23788 31732 23841 31772
rect 23980 31732 24033 31772
rect 29548 31732 29601 31772
rect 29740 31732 29793 31772
rect 17547 31688 17589 31697
rect 17547 31648 17548 31688
rect 17588 31648 17589 31688
rect 17547 31639 17589 31648
rect 16312 31520 16354 31529
rect 16312 31480 16313 31520
rect 16353 31480 16354 31520
rect 16312 31471 16354 31480
rect 16491 31520 16533 31529
rect 16491 31480 16492 31520
rect 16532 31480 16533 31520
rect 16491 31471 16533 31480
rect 16313 31374 16353 31471
rect 18041 31374 18081 31732
rect 18232 31688 18274 31697
rect 18232 31648 18233 31688
rect 18273 31648 18274 31688
rect 18232 31639 18274 31648
rect 18233 31374 18273 31639
rect 18809 31374 18849 31732
rect 19577 31374 19617 31732
rect 23801 31374 23841 31732
rect 23993 31374 24033 31732
rect 29561 31374 29601 31732
rect 29753 31374 29793 31732
rect 30175 31732 30260 31772
rect 31519 31732 31700 31772
rect 32044 31772 32084 34327
rect 32812 31772 32852 35083
rect 32908 34889 32948 36511
rect 33003 36224 33045 36233
rect 33003 36184 33004 36224
rect 33044 36184 33045 36224
rect 33003 36175 33045 36184
rect 32907 34880 32949 34889
rect 32907 34840 32908 34880
rect 32948 34840 32949 34880
rect 32907 34831 32949 34840
rect 33004 31772 33044 36175
rect 33196 34049 33236 37192
rect 33292 37183 33332 37192
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 33772 36149 33812 37948
rect 33868 36485 33908 38191
rect 33963 37988 34005 37997
rect 33963 37948 33964 37988
rect 34004 37948 34005 37988
rect 33963 37939 34005 37948
rect 35691 37988 35733 37997
rect 35691 37948 35692 37988
rect 35732 37948 35733 37988
rect 35691 37939 35733 37948
rect 37132 37988 37172 37997
rect 33964 37854 34004 37939
rect 34443 37400 34485 37409
rect 34443 37360 34444 37400
rect 34484 37360 34485 37400
rect 34443 37351 34485 37360
rect 35308 37400 35348 37409
rect 33963 37316 34005 37325
rect 33963 37276 33964 37316
rect 34004 37276 34005 37316
rect 33963 37267 34005 37276
rect 33964 36728 34004 37267
rect 33867 36476 33909 36485
rect 33867 36436 33868 36476
rect 33908 36436 33909 36476
rect 33867 36427 33909 36436
rect 33771 36140 33813 36149
rect 33771 36100 33772 36140
rect 33812 36100 33813 36140
rect 33771 36091 33813 36100
rect 33387 35972 33429 35981
rect 33387 35932 33388 35972
rect 33428 35932 33429 35972
rect 33387 35923 33429 35932
rect 33388 35477 33428 35923
rect 33387 35468 33429 35477
rect 33387 35428 33388 35468
rect 33428 35428 33429 35468
rect 33387 35419 33429 35428
rect 33388 35384 33428 35419
rect 33388 35333 33428 35344
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 33964 34637 34004 36688
rect 34444 36308 34484 37351
rect 35308 37241 35348 37360
rect 35692 37400 35732 37939
rect 37132 37460 37172 37948
rect 36556 37409 36596 37440
rect 37132 37420 37364 37460
rect 35692 37351 35732 37360
rect 36555 37400 36597 37409
rect 36555 37360 36556 37400
rect 36596 37360 36597 37400
rect 36555 37351 36597 37360
rect 36652 37400 36692 37409
rect 36940 37400 36980 37409
rect 36692 37360 36884 37400
rect 36652 37351 36692 37360
rect 36556 37316 36596 37351
rect 35307 37232 35349 37241
rect 35307 37192 35308 37232
rect 35348 37192 35349 37232
rect 36459 37232 36501 37241
rect 35307 37183 35349 37192
rect 36268 37190 36308 37199
rect 36459 37192 36460 37232
rect 36500 37192 36501 37232
rect 36459 37183 36501 37192
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 36076 36812 36116 36821
rect 36268 36812 36308 37150
rect 36116 36772 36308 36812
rect 36076 36763 36116 36772
rect 35308 36728 35348 36737
rect 35308 36644 35348 36688
rect 34828 36604 35348 36644
rect 35500 36728 35540 36737
rect 34444 36268 34580 36308
rect 34348 35720 34388 35729
rect 34540 35720 34580 36268
rect 33387 34628 33429 34637
rect 33387 34588 33388 34628
rect 33428 34588 33429 34628
rect 33387 34579 33429 34588
rect 33963 34628 34005 34637
rect 33963 34588 33964 34628
rect 34004 34588 34005 34628
rect 33963 34579 34005 34588
rect 33388 34376 33428 34579
rect 34348 34385 34388 35680
rect 34507 35680 34580 35720
rect 34828 35888 34868 36604
rect 35116 36476 35156 36485
rect 35308 36476 35348 36485
rect 35116 36233 35156 36436
rect 35212 36436 35308 36476
rect 35115 36224 35157 36233
rect 35115 36184 35116 36224
rect 35156 36184 35157 36224
rect 35115 36175 35157 36184
rect 35116 36056 35156 36065
rect 35020 36016 35116 36056
rect 34923 35972 34965 35981
rect 34923 35932 34924 35972
rect 34964 35932 34965 35972
rect 34923 35923 34965 35932
rect 34828 35720 34868 35848
rect 34924 35888 34964 35923
rect 34924 35837 34964 35848
rect 35020 35804 35060 36016
rect 35116 36007 35156 36016
rect 35116 35899 35156 35908
rect 35212 35888 35252 36436
rect 35308 36427 35348 36436
rect 35500 36065 35540 36688
rect 35691 36728 35733 36737
rect 35691 36688 35692 36728
rect 35732 36688 35733 36728
rect 35691 36679 35733 36688
rect 35884 36728 35924 36737
rect 36460 36728 36500 37183
rect 35692 36485 35732 36679
rect 35788 36644 35828 36653
rect 35691 36476 35733 36485
rect 35691 36436 35692 36476
rect 35732 36436 35733 36476
rect 35691 36427 35733 36436
rect 35788 36224 35828 36604
rect 35884 36308 35924 36688
rect 36364 36688 36460 36728
rect 35884 36268 36116 36308
rect 35788 36184 36020 36224
rect 35499 36056 35541 36065
rect 35499 36016 35500 36056
rect 35540 36016 35541 36056
rect 35499 36007 35541 36016
rect 35307 35972 35349 35981
rect 35307 35932 35308 35972
rect 35348 35932 35349 35972
rect 35307 35923 35349 35932
rect 35156 35859 35252 35888
rect 35116 35848 35252 35859
rect 35308 35838 35348 35923
rect 35404 35888 35444 35897
rect 35404 35804 35444 35848
rect 35596 35888 35636 35897
rect 35691 35888 35733 35897
rect 35636 35848 35692 35888
rect 35732 35848 35733 35888
rect 35596 35839 35636 35848
rect 35691 35839 35733 35848
rect 35788 35888 35828 35897
rect 35020 35764 35252 35804
rect 35404 35764 35446 35804
rect 34828 35680 35156 35720
rect 34507 35552 34547 35680
rect 34492 35512 34547 35552
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34492 35384 34532 35512
rect 34592 35503 34960 35512
rect 34492 35344 34580 35384
rect 34540 35225 34580 35344
rect 34539 35216 34581 35225
rect 34539 35176 34540 35216
rect 34580 35176 34581 35216
rect 34539 35167 34581 35176
rect 34540 35082 34580 35167
rect 35116 35057 35156 35680
rect 35212 35309 35252 35764
rect 35406 35645 35446 35764
rect 35403 35636 35446 35645
rect 35403 35596 35404 35636
rect 35444 35596 35446 35636
rect 35692 35720 35732 35729
rect 35403 35587 35445 35596
rect 35211 35300 35253 35309
rect 35211 35260 35212 35300
rect 35252 35260 35253 35300
rect 35211 35251 35253 35260
rect 35404 35216 35444 35225
rect 35404 35057 35444 35176
rect 35115 35048 35157 35057
rect 35115 35008 35116 35048
rect 35156 35008 35157 35048
rect 35115 34999 35157 35008
rect 35403 35048 35445 35057
rect 35403 35008 35404 35048
rect 35444 35008 35445 35048
rect 35403 34999 35445 35008
rect 35692 34889 35732 35680
rect 35788 35477 35828 35848
rect 35980 35888 36020 36184
rect 36076 35981 36116 36268
rect 36364 36065 36404 36688
rect 36460 36679 36500 36688
rect 36363 36056 36405 36065
rect 36363 36016 36364 36056
rect 36404 36016 36405 36056
rect 36363 36007 36405 36016
rect 36460 36056 36500 36065
rect 36075 35972 36117 35981
rect 36075 35932 36076 35972
rect 36116 35932 36117 35972
rect 36075 35923 36117 35932
rect 35980 35839 36020 35848
rect 36171 35888 36213 35897
rect 36171 35848 36172 35888
rect 36212 35848 36213 35888
rect 36171 35839 36213 35848
rect 36268 35888 36308 35897
rect 36172 35754 36212 35839
rect 36076 35720 36116 35729
rect 35787 35468 35829 35477
rect 35787 35428 35788 35468
rect 35828 35428 35829 35468
rect 35787 35419 35829 35428
rect 35787 35300 35829 35309
rect 35787 35260 35788 35300
rect 35828 35260 35829 35300
rect 35787 35251 35829 35260
rect 35980 35300 36020 35309
rect 36076 35300 36116 35680
rect 36171 35468 36213 35477
rect 36171 35428 36172 35468
rect 36212 35428 36213 35468
rect 36171 35419 36213 35428
rect 36020 35260 36116 35300
rect 35980 35251 36020 35260
rect 35788 35166 35828 35251
rect 36172 35141 36212 35419
rect 36171 35132 36213 35141
rect 36171 35092 36172 35132
rect 36212 35092 36213 35132
rect 36171 35083 36213 35092
rect 35691 34880 35733 34889
rect 35691 34840 35692 34880
rect 35732 34840 35733 34880
rect 35691 34831 35733 34840
rect 36268 34721 36308 35848
rect 36364 35216 36404 36007
rect 36364 35057 36404 35176
rect 36363 35048 36405 35057
rect 36363 35008 36364 35048
rect 36404 35008 36405 35048
rect 36363 34999 36405 35008
rect 36363 34796 36405 34805
rect 36363 34756 36364 34796
rect 36404 34756 36405 34796
rect 36363 34747 36405 34756
rect 36267 34712 36309 34721
rect 36267 34672 36268 34712
rect 36308 34672 36309 34712
rect 36267 34663 36309 34672
rect 35691 34544 35733 34553
rect 35691 34504 35692 34544
rect 35732 34504 35733 34544
rect 35691 34495 35733 34504
rect 33388 34327 33428 34336
rect 34347 34376 34389 34385
rect 34347 34336 34348 34376
rect 34388 34336 34389 34376
rect 34347 34327 34389 34336
rect 35692 34376 35732 34495
rect 35692 34327 35732 34336
rect 36268 34376 36308 34385
rect 36364 34376 36404 34747
rect 36308 34336 36404 34376
rect 36268 34327 36308 34336
rect 34540 34217 34580 34302
rect 34539 34208 34581 34217
rect 34539 34168 34540 34208
rect 34580 34168 34581 34208
rect 34539 34159 34581 34168
rect 35212 34208 35252 34217
rect 33195 34040 33237 34049
rect 33195 34000 33196 34040
rect 33236 34000 33237 34040
rect 33195 33991 33237 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 35212 32621 35252 34168
rect 35211 32612 35253 32621
rect 35211 32572 35212 32612
rect 35252 32572 35253 32612
rect 35211 32563 35253 32572
rect 36460 32537 36500 36016
rect 36556 35888 36596 37276
rect 36844 37241 36884 37360
rect 36843 37232 36885 37241
rect 36843 37192 36844 37232
rect 36884 37192 36885 37232
rect 36843 37183 36885 37192
rect 36748 35888 36788 35897
rect 36556 35848 36748 35888
rect 36748 35839 36788 35848
rect 36844 35888 36884 37183
rect 36940 36737 36980 37360
rect 37324 37400 37364 37420
rect 37420 37409 37460 38158
rect 37324 37351 37364 37360
rect 37419 37400 37461 37409
rect 37419 37360 37420 37400
rect 37460 37360 37461 37400
rect 37419 37351 37461 37360
rect 36939 36728 36981 36737
rect 37324 36728 37364 36737
rect 36939 36688 36940 36728
rect 36980 36688 36981 36728
rect 36939 36679 36981 36688
rect 37228 36688 37324 36728
rect 36844 35839 36884 35848
rect 36940 34805 36980 36679
rect 37131 35972 37173 35981
rect 37131 35932 37132 35972
rect 37172 35932 37173 35972
rect 37131 35923 37173 35932
rect 37132 35888 37172 35923
rect 37132 35837 37172 35848
rect 37228 35225 37268 36688
rect 37324 36679 37364 36688
rect 37516 35897 37556 38200
rect 37804 38240 37844 38249
rect 37708 37400 37748 37409
rect 37708 36065 37748 37360
rect 37804 36905 37844 38200
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 44043 37484 44085 37493
rect 44043 37444 44044 37484
rect 44084 37444 44085 37484
rect 44043 37435 44085 37444
rect 38379 37400 38421 37409
rect 38379 37360 38380 37400
rect 38420 37360 38421 37400
rect 38379 37351 38421 37360
rect 38571 37400 38613 37409
rect 38571 37360 38572 37400
rect 38612 37360 38613 37400
rect 38571 37351 38613 37360
rect 41068 37400 41108 37409
rect 37803 36896 37845 36905
rect 37803 36856 37804 36896
rect 37844 36856 37845 36896
rect 38380 36896 38420 37351
rect 38572 37266 38612 37351
rect 39724 37232 39764 37241
rect 38476 36896 38516 36905
rect 38380 36856 38476 36896
rect 37803 36847 37845 36856
rect 38476 36847 38516 36856
rect 37804 36401 37844 36847
rect 39627 36728 39669 36737
rect 39627 36688 39628 36728
rect 39668 36688 39669 36728
rect 39627 36679 39669 36688
rect 39628 36594 39668 36679
rect 37803 36392 37845 36401
rect 37803 36352 37804 36392
rect 37844 36352 37845 36392
rect 37803 36343 37845 36352
rect 39627 36392 39669 36401
rect 39627 36352 39628 36392
rect 39668 36352 39669 36392
rect 39627 36343 39669 36352
rect 37707 36056 37749 36065
rect 37707 36016 37708 36056
rect 37748 36016 37749 36056
rect 37707 36007 37749 36016
rect 39147 36056 39189 36065
rect 39147 36016 39148 36056
rect 39188 36016 39189 36056
rect 39147 36007 39189 36016
rect 37515 35888 37557 35897
rect 37515 35848 37516 35888
rect 37556 35848 37557 35888
rect 37515 35839 37557 35848
rect 38379 35636 38421 35645
rect 38379 35596 38380 35636
rect 38420 35596 38421 35636
rect 38379 35587 38421 35596
rect 38380 35384 38420 35587
rect 38380 35335 38420 35344
rect 37227 35216 37269 35225
rect 37227 35176 37228 35216
rect 37268 35176 37269 35216
rect 37227 35167 37269 35176
rect 37228 35082 37268 35167
rect 36939 34796 36981 34805
rect 36939 34756 36940 34796
rect 36980 34756 36981 34796
rect 36939 34747 36981 34756
rect 36940 34544 36980 34553
rect 36556 34376 36596 34385
rect 36556 34217 36596 34336
rect 36652 34292 36692 34301
rect 36555 34208 36597 34217
rect 36555 34168 36556 34208
rect 36596 34168 36597 34208
rect 36555 34159 36597 34168
rect 36652 34133 36692 34252
rect 36651 34124 36693 34133
rect 36651 34084 36652 34124
rect 36692 34084 36693 34124
rect 36651 34075 36693 34084
rect 36652 33881 36692 34075
rect 36940 33965 36980 34504
rect 38091 34544 38133 34553
rect 38091 34504 38092 34544
rect 38132 34504 38133 34544
rect 38091 34495 38133 34504
rect 38092 34376 38132 34495
rect 38092 34217 38132 34336
rect 39148 34376 39188 36007
rect 39628 35216 39668 36343
rect 39724 35897 39764 37192
rect 39915 37232 39957 37241
rect 39915 37192 39916 37232
rect 39956 37192 40052 37232
rect 39915 37183 39957 37192
rect 39916 37098 39956 37183
rect 40012 36812 40052 37192
rect 40012 36763 40052 36772
rect 41068 36737 41108 37360
rect 41932 37400 41972 37409
rect 39916 36728 39956 36737
rect 39916 36224 39956 36688
rect 40107 36728 40149 36737
rect 40107 36688 40108 36728
rect 40148 36688 40149 36728
rect 40107 36679 40149 36688
rect 41067 36728 41109 36737
rect 41067 36688 41068 36728
rect 41108 36688 41109 36728
rect 41067 36679 41109 36688
rect 41548 36728 41588 36737
rect 41932 36728 41972 37360
rect 41588 36688 41684 36728
rect 41548 36679 41588 36688
rect 39916 36184 40052 36224
rect 40012 35897 40052 36184
rect 39723 35888 39765 35897
rect 39916 35888 39956 35897
rect 39723 35848 39724 35888
rect 39764 35848 39916 35888
rect 39723 35839 39765 35848
rect 39916 35839 39956 35848
rect 40011 35888 40053 35897
rect 40011 35848 40012 35888
rect 40052 35848 40053 35888
rect 40011 35839 40053 35848
rect 40012 35216 40052 35225
rect 39628 35176 40012 35216
rect 40012 35167 40052 35176
rect 39148 34327 39188 34336
rect 40012 34376 40052 34385
rect 40108 34376 40148 36679
rect 40971 36644 41013 36653
rect 40971 36604 40972 36644
rect 41012 36604 41013 36644
rect 40971 36595 41013 36604
rect 40299 36560 40341 36569
rect 40299 36520 40300 36560
rect 40340 36520 40341 36560
rect 40299 36511 40341 36520
rect 40300 36426 40340 36511
rect 40588 36056 40628 36065
rect 40204 35888 40244 35899
rect 40204 35813 40244 35848
rect 40299 35888 40341 35897
rect 40299 35848 40300 35888
rect 40340 35848 40341 35888
rect 40299 35839 40341 35848
rect 40203 35804 40245 35813
rect 40203 35764 40204 35804
rect 40244 35764 40245 35804
rect 40203 35755 40245 35764
rect 40300 35754 40340 35839
rect 40395 35804 40437 35813
rect 40395 35764 40396 35804
rect 40436 35764 40437 35804
rect 40395 35755 40437 35764
rect 40396 35468 40436 35755
rect 40588 35561 40628 36016
rect 40972 35888 41012 36595
rect 41644 36140 41684 36688
rect 41932 36485 41972 36688
rect 42316 37316 42356 37325
rect 42316 36569 42356 37276
rect 42795 36728 42837 36737
rect 42795 36688 42796 36728
rect 42836 36688 42837 36728
rect 42795 36679 42837 36688
rect 42315 36560 42357 36569
rect 42315 36520 42316 36560
rect 42356 36520 42357 36560
rect 42315 36511 42357 36520
rect 41931 36476 41973 36485
rect 41931 36436 41932 36476
rect 41972 36436 41973 36476
rect 41931 36427 41973 36436
rect 41644 36091 41684 36100
rect 41163 36056 41205 36065
rect 41163 36016 41164 36056
rect 41204 36016 41205 36056
rect 41163 36007 41205 36016
rect 40972 35839 41012 35848
rect 40587 35552 40629 35561
rect 40587 35512 40588 35552
rect 40628 35512 40629 35552
rect 40587 35503 40629 35512
rect 40300 35428 40436 35468
rect 40300 35216 40340 35428
rect 40300 35167 40340 35176
rect 40396 35216 40436 35225
rect 40396 35048 40436 35176
rect 40876 35216 40916 35225
rect 41164 35216 41204 36007
rect 41260 35888 41300 35899
rect 41260 35813 41300 35848
rect 41355 35888 41397 35897
rect 41355 35848 41356 35888
rect 41396 35848 41397 35888
rect 41355 35839 41397 35848
rect 41259 35804 41301 35813
rect 41259 35764 41260 35804
rect 41300 35764 41301 35804
rect 41259 35755 41301 35764
rect 41356 35754 41396 35839
rect 41260 35216 41300 35225
rect 41164 35176 41260 35216
rect 40052 34336 40148 34376
rect 40300 35008 40436 35048
rect 40684 35048 40724 35057
rect 40876 35048 40916 35176
rect 41260 35167 41300 35176
rect 42124 35216 42164 35227
rect 42124 35141 42164 35176
rect 42796 35141 42836 36679
rect 43948 36476 43988 36485
rect 43852 36436 43948 36476
rect 43756 36056 43796 36065
rect 43084 35888 43124 35897
rect 42123 35132 42165 35141
rect 42123 35092 42124 35132
rect 42164 35092 42165 35132
rect 42123 35083 42165 35092
rect 42795 35132 42837 35141
rect 42795 35092 42796 35132
rect 42836 35092 42837 35132
rect 42795 35083 42837 35092
rect 40724 35008 40916 35048
rect 40012 34327 40052 34336
rect 38764 34292 38804 34301
rect 37612 34208 37652 34217
rect 36939 33956 36981 33965
rect 36939 33916 36940 33956
rect 36980 33916 36981 33956
rect 36939 33907 36981 33916
rect 36651 33872 36693 33881
rect 36651 33832 36652 33872
rect 36692 33832 36693 33872
rect 36651 33823 36693 33832
rect 36459 32528 36501 32537
rect 36459 32488 36460 32528
rect 36500 32488 36501 32528
rect 36459 32479 36501 32488
rect 37612 32453 37652 34168
rect 38091 34208 38133 34217
rect 38091 34168 38092 34208
rect 38132 34168 38133 34208
rect 38091 34159 38133 34168
rect 38764 33965 38804 34252
rect 40300 33965 40340 35008
rect 40684 34999 40724 35008
rect 43084 34973 43124 35848
rect 43372 35888 43412 35897
rect 43275 35804 43317 35813
rect 43275 35764 43276 35804
rect 43316 35764 43317 35804
rect 43275 35755 43317 35764
rect 43276 35384 43316 35755
rect 43276 35335 43316 35344
rect 43372 35216 43412 35848
rect 43276 35176 43412 35216
rect 43468 35804 43508 35813
rect 43083 34964 43125 34973
rect 43083 34924 43084 34964
rect 43124 34924 43125 34964
rect 43083 34915 43125 34924
rect 42220 34376 42260 34385
rect 42220 34217 42260 34336
rect 41164 34208 41204 34217
rect 38763 33956 38805 33965
rect 38763 33916 38764 33956
rect 38804 33916 38805 33956
rect 38763 33907 38805 33916
rect 40299 33956 40341 33965
rect 40299 33916 40300 33956
rect 40340 33916 40341 33956
rect 40299 33907 40341 33916
rect 41164 33881 41204 34168
rect 42219 34208 42261 34217
rect 42219 34168 42220 34208
rect 42260 34168 42261 34208
rect 42219 34159 42261 34168
rect 43276 33881 43316 35176
rect 43468 35132 43508 35764
rect 43659 35804 43701 35813
rect 43659 35764 43660 35804
rect 43700 35764 43701 35804
rect 43659 35755 43701 35764
rect 43372 35092 43508 35132
rect 43660 35132 43700 35755
rect 43372 34049 43412 35092
rect 43660 35083 43700 35092
rect 43467 34964 43509 34973
rect 43467 34924 43468 34964
rect 43508 34924 43509 34964
rect 43756 34964 43796 36016
rect 43852 35897 43892 36436
rect 43948 36427 43988 36436
rect 43948 35972 43988 35981
rect 44044 35972 44084 37435
rect 69291 37400 69333 37409
rect 69291 37360 69292 37400
rect 69332 37360 69333 37400
rect 69291 37351 69333 37360
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 46252 36056 46292 36065
rect 43988 35932 44084 35972
rect 44523 35972 44565 35981
rect 44523 35932 44524 35972
rect 44564 35932 44565 35972
rect 43948 35923 43988 35932
rect 44523 35923 44565 35932
rect 43851 35888 43893 35897
rect 43851 35848 43852 35888
rect 43892 35848 43893 35888
rect 43851 35839 43893 35848
rect 44524 35838 44564 35923
rect 45580 35888 45620 35897
rect 45580 35813 45620 35848
rect 45867 35888 45909 35897
rect 45867 35848 45868 35888
rect 45908 35848 45909 35888
rect 45867 35839 45909 35848
rect 44139 35804 44181 35813
rect 44139 35764 44140 35804
rect 44180 35764 44181 35804
rect 44139 35755 44181 35764
rect 45579 35804 45621 35813
rect 45579 35764 45580 35804
rect 45620 35764 45621 35804
rect 45579 35755 45621 35764
rect 43947 35720 43989 35729
rect 43947 35680 43948 35720
rect 43988 35680 43989 35720
rect 43947 35671 43989 35680
rect 44140 35720 44180 35755
rect 43948 35132 43988 35671
rect 44140 35669 44180 35680
rect 44715 35720 44757 35729
rect 44715 35680 44716 35720
rect 44756 35680 44757 35720
rect 44715 35671 44757 35680
rect 44716 35586 44756 35671
rect 44331 35468 44373 35477
rect 44331 35428 44332 35468
rect 44372 35428 44373 35468
rect 44331 35419 44373 35428
rect 44332 35384 44372 35419
rect 44332 35333 44372 35344
rect 44139 35216 44181 35225
rect 44139 35176 44140 35216
rect 44180 35176 44181 35216
rect 44139 35167 44181 35176
rect 45484 35216 45524 35227
rect 43948 35083 43988 35092
rect 44140 34964 44180 35167
rect 45484 35141 45524 35176
rect 45483 35132 45525 35141
rect 45483 35092 45484 35132
rect 45524 35092 45525 35132
rect 45483 35083 45525 35092
rect 43756 34924 43988 34964
rect 43467 34915 43509 34924
rect 43468 34830 43508 34915
rect 43660 34376 43700 34385
rect 43371 34040 43413 34049
rect 43371 34000 43372 34040
rect 43412 34000 43413 34040
rect 43371 33991 43413 34000
rect 41163 33872 41205 33881
rect 41163 33832 41164 33872
rect 41204 33832 41205 33872
rect 41163 33823 41205 33832
rect 43275 33872 43317 33881
rect 43275 33832 43276 33872
rect 43316 33832 43317 33872
rect 43275 33823 43317 33832
rect 43660 32453 43700 34336
rect 43948 34376 43988 34924
rect 44140 34376 44180 34924
rect 44332 34376 44372 34385
rect 44140 34336 44332 34376
rect 43948 34327 43988 34336
rect 44332 34327 44372 34336
rect 45195 34376 45237 34385
rect 45195 34336 45196 34376
rect 45236 34336 45237 34376
rect 45195 34327 45237 34336
rect 45196 34242 45236 34327
rect 45580 32705 45620 35755
rect 45868 35754 45908 35839
rect 45964 35804 46004 35813
rect 45964 35477 46004 35764
rect 46252 35636 46292 36016
rect 47979 36056 48021 36065
rect 47979 36016 47980 36056
rect 48020 36016 48021 36056
rect 47979 36007 48021 36016
rect 49612 36056 49652 36065
rect 47019 35888 47061 35897
rect 47019 35848 47020 35888
rect 47060 35848 47061 35888
rect 47019 35839 47061 35848
rect 47211 35888 47253 35897
rect 47211 35848 47212 35888
rect 47252 35848 47253 35888
rect 47211 35839 47253 35848
rect 46252 35596 46772 35636
rect 45963 35468 46005 35477
rect 45963 35428 45964 35468
rect 46004 35428 46005 35468
rect 45963 35419 46005 35428
rect 46732 35300 46772 35596
rect 46732 35251 46772 35260
rect 46347 35216 46389 35225
rect 46347 35176 46348 35216
rect 46388 35176 46389 35216
rect 46347 35167 46389 35176
rect 46924 35216 46964 35225
rect 46348 35082 46388 35167
rect 46540 34628 46580 34637
rect 46924 34628 46964 35176
rect 47020 34721 47060 35839
rect 47212 34973 47252 35839
rect 47307 35216 47349 35225
rect 47307 35176 47308 35216
rect 47348 35176 47349 35216
rect 47307 35167 47349 35176
rect 47308 35057 47348 35167
rect 47307 35048 47349 35057
rect 47307 35008 47308 35048
rect 47348 35008 47349 35048
rect 47307 34999 47349 35008
rect 47211 34964 47253 34973
rect 47211 34924 47212 34964
rect 47252 34924 47253 34964
rect 47211 34915 47253 34924
rect 47019 34712 47061 34721
rect 47019 34672 47020 34712
rect 47060 34672 47061 34712
rect 47019 34663 47061 34672
rect 46580 34588 46964 34628
rect 46540 34579 46580 34588
rect 47020 34544 47060 34663
rect 46828 34504 47060 34544
rect 46828 34376 46868 34504
rect 46828 34327 46868 34336
rect 46924 34376 46964 34385
rect 46348 34208 46388 34217
rect 46348 34049 46388 34168
rect 46347 34040 46389 34049
rect 46347 34000 46348 34040
rect 46388 34000 46389 34040
rect 46347 33991 46389 34000
rect 46924 33965 46964 34336
rect 47212 34376 47252 34915
rect 47980 34628 48020 36007
rect 48939 35888 48981 35897
rect 48939 35848 48940 35888
rect 48980 35848 48981 35888
rect 48939 35839 48981 35848
rect 49228 35888 49268 35897
rect 48940 35754 48980 35839
rect 48172 35216 48212 35225
rect 48172 35057 48212 35176
rect 48171 35048 48213 35057
rect 48171 35008 48172 35048
rect 48212 35008 48213 35048
rect 48171 34999 48213 35008
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 48075 34712 48117 34721
rect 48075 34672 48076 34712
rect 48116 34672 48117 34712
rect 48075 34663 48117 34672
rect 47980 34579 48020 34588
rect 47212 34327 47252 34336
rect 46923 33956 46965 33965
rect 46923 33916 46924 33956
rect 46964 33916 46965 33956
rect 46923 33907 46965 33916
rect 45579 32696 45621 32705
rect 45579 32656 45580 32696
rect 45620 32656 45621 32696
rect 45579 32647 45621 32656
rect 37611 32444 37653 32453
rect 37611 32404 37612 32444
rect 37652 32404 37653 32444
rect 37611 32395 37653 32404
rect 43659 32444 43701 32453
rect 43659 32404 43660 32444
rect 43700 32404 43701 32444
rect 43659 32395 43701 32404
rect 48076 31772 48116 34663
rect 49228 34049 49268 35848
rect 49324 35804 49364 35813
rect 49324 35645 49364 35764
rect 49323 35636 49365 35645
rect 49323 35596 49324 35636
rect 49364 35596 49365 35636
rect 49323 35587 49365 35596
rect 49516 35300 49556 35309
rect 49612 35300 49652 36016
rect 51340 36056 51380 36065
rect 50667 35888 50709 35897
rect 50667 35848 50668 35888
rect 50708 35848 50709 35888
rect 50667 35839 50709 35848
rect 50956 35888 50996 35899
rect 50668 35754 50708 35839
rect 50956 35813 50996 35848
rect 50955 35804 50997 35813
rect 50955 35764 50956 35804
rect 50996 35764 50997 35804
rect 50955 35755 50997 35764
rect 51052 35804 51092 35813
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 49556 35260 49652 35300
rect 49516 35251 49556 35260
rect 49900 35216 49940 35225
rect 49900 34973 49940 35176
rect 50764 35216 50804 35225
rect 50764 35057 50804 35176
rect 50763 35048 50805 35057
rect 50763 35008 50764 35048
rect 50804 35008 50805 35048
rect 50763 34999 50805 35008
rect 49324 34964 49364 34973
rect 49324 34721 49364 34924
rect 49899 34964 49941 34973
rect 49899 34924 49900 34964
rect 49940 34924 49941 34964
rect 49899 34915 49941 34924
rect 49900 34805 49940 34915
rect 49899 34796 49941 34805
rect 49899 34756 49900 34796
rect 49940 34756 49941 34796
rect 49899 34747 49941 34756
rect 49323 34712 49365 34721
rect 49323 34672 49324 34712
rect 49364 34672 49365 34712
rect 49323 34663 49365 34672
rect 49419 34544 49461 34553
rect 49419 34504 49420 34544
rect 49460 34504 49461 34544
rect 49419 34495 49461 34504
rect 49611 34544 49653 34553
rect 49611 34504 49612 34544
rect 49652 34504 49653 34544
rect 49611 34495 49653 34504
rect 48939 34040 48981 34049
rect 48939 34000 48940 34040
rect 48980 34000 48981 34040
rect 48939 33991 48981 34000
rect 49227 34040 49269 34049
rect 49227 34000 49228 34040
rect 49268 34000 49269 34040
rect 49227 33991 49269 34000
rect 32044 31732 32097 31772
rect 32812 31732 32865 31772
rect 33004 31732 33057 31772
rect 30175 31374 30215 31732
rect 31519 31374 31559 31732
rect 32057 31374 32097 31732
rect 32825 31374 32865 31732
rect 33017 31374 33057 31732
rect 47993 31732 48116 31772
rect 48940 31772 48980 33991
rect 49420 33881 49460 34495
rect 49612 34376 49652 34495
rect 49612 34327 49652 34336
rect 50860 34376 50900 34385
rect 50860 34217 50900 34336
rect 50380 34208 50420 34217
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 49419 33872 49461 33881
rect 49419 33832 49420 33872
rect 49460 33832 49461 33872
rect 49419 33823 49461 33832
rect 49131 33620 49173 33629
rect 49131 33580 49132 33620
rect 49172 33580 49173 33620
rect 49131 33571 49173 33580
rect 49132 31772 49172 33571
rect 50380 31781 50420 34168
rect 50859 34208 50901 34217
rect 50859 34168 50860 34208
rect 50900 34168 50901 34208
rect 50859 34159 50901 34168
rect 50860 34049 50900 34159
rect 50859 34040 50901 34049
rect 50859 34000 50860 34040
rect 50900 34000 50901 34040
rect 50859 33991 50901 34000
rect 51052 33629 51092 35764
rect 51340 33713 51380 36016
rect 52300 36056 52340 36065
rect 51627 35888 51669 35897
rect 51627 35848 51628 35888
rect 51668 35848 51669 35888
rect 51627 35839 51669 35848
rect 51916 35888 51956 35897
rect 51628 35754 51668 35839
rect 51916 35645 51956 35848
rect 52011 35804 52053 35813
rect 52011 35764 52012 35804
rect 52052 35764 52053 35804
rect 52011 35755 52053 35764
rect 51915 35636 51957 35645
rect 51915 35596 51916 35636
rect 51956 35596 51957 35636
rect 51915 35587 51957 35596
rect 51916 35384 51956 35587
rect 51916 35335 51956 35344
rect 51916 34964 51956 34975
rect 52012 34973 52052 35755
rect 52300 35636 52340 36016
rect 52108 35596 52340 35636
rect 52108 35300 52148 35596
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 52108 35251 52148 35260
rect 52492 35216 52532 35225
rect 51916 34889 51956 34924
rect 52011 34964 52053 34973
rect 52011 34924 52012 34964
rect 52052 34924 52053 34964
rect 52011 34915 52053 34924
rect 51915 34880 51957 34889
rect 51915 34840 51916 34880
rect 51956 34840 51957 34880
rect 51915 34831 51957 34840
rect 52492 34805 52532 35176
rect 53356 35216 53396 35225
rect 53356 35057 53396 35176
rect 64588 35216 64628 35225
rect 53355 35048 53397 35057
rect 53355 35008 53356 35048
rect 53396 35008 53397 35048
rect 53355 34999 53397 35008
rect 54027 35048 54069 35057
rect 54027 35008 54028 35048
rect 54068 35008 54069 35048
rect 54027 34999 54069 35008
rect 64395 35048 64437 35057
rect 64395 35008 64396 35048
rect 64436 35008 64437 35048
rect 64395 34999 64437 35008
rect 53835 34964 53877 34973
rect 53835 34924 53836 34964
rect 53876 34924 53877 34964
rect 53835 34915 53877 34924
rect 52971 34880 53013 34889
rect 52971 34840 52972 34880
rect 53012 34840 53013 34880
rect 52971 34831 53013 34840
rect 52491 34796 52533 34805
rect 52491 34756 52492 34796
rect 52532 34756 52533 34796
rect 52491 34747 52533 34756
rect 52492 34376 52532 34385
rect 52012 34208 52052 34217
rect 51339 33704 51381 33713
rect 51339 33664 51340 33704
rect 51380 33664 51381 33704
rect 51339 33655 51381 33664
rect 51051 33620 51093 33629
rect 51051 33580 51052 33620
rect 51092 33580 51093 33620
rect 51051 33571 51093 33580
rect 52012 32621 52052 34168
rect 52299 34208 52341 34217
rect 52299 34168 52300 34208
rect 52340 34168 52341 34208
rect 52299 34159 52341 34168
rect 52300 33881 52340 34159
rect 52492 34049 52532 34336
rect 52780 34292 52820 34301
rect 52491 34040 52533 34049
rect 52491 34000 52492 34040
rect 52532 34000 52533 34040
rect 52491 33991 52533 34000
rect 52299 33872 52341 33881
rect 52299 33832 52300 33872
rect 52340 33832 52341 33872
rect 52299 33823 52341 33832
rect 52780 33713 52820 34252
rect 52779 33704 52821 33713
rect 52779 33664 52780 33704
rect 52820 33664 52821 33704
rect 52779 33655 52821 33664
rect 52011 32612 52053 32621
rect 52011 32572 52012 32612
rect 52052 32572 52053 32612
rect 52011 32563 52053 32572
rect 50379 31772 50421 31781
rect 48940 31732 48993 31772
rect 49132 31732 49185 31772
rect 47993 31374 48033 31732
rect 48953 31374 48993 31732
rect 49145 31374 49185 31732
rect 50379 31732 50380 31772
rect 50420 31732 50421 31772
rect 52972 31772 53012 34831
rect 53163 34796 53205 34805
rect 53163 34756 53164 34796
rect 53204 34756 53205 34796
rect 53163 34747 53205 34756
rect 53164 34376 53204 34747
rect 53164 33797 53204 34336
rect 53163 33788 53205 33797
rect 53163 33748 53164 33788
rect 53204 33748 53205 33788
rect 53163 33739 53205 33748
rect 53836 31772 53876 34915
rect 54028 34376 54068 34999
rect 54507 34964 54549 34973
rect 54507 34924 54508 34964
rect 54548 34924 54549 34964
rect 54507 34915 54549 34924
rect 54508 34830 54548 34915
rect 64396 34914 64436 34999
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 64588 34385 64628 35176
rect 65451 35216 65493 35225
rect 65451 35176 65452 35216
rect 65492 35176 65493 35216
rect 65451 35167 65493 35176
rect 54028 33881 54068 34336
rect 61516 34376 61556 34385
rect 55180 34208 55220 34217
rect 54027 33872 54069 33881
rect 54027 33832 54028 33872
rect 54068 33832 54069 33872
rect 54027 33823 54069 33832
rect 55180 33629 55220 34168
rect 61516 34049 61556 34336
rect 62476 34376 62516 34385
rect 62476 34049 62516 34336
rect 62764 34376 62804 34385
rect 62764 34217 62804 34336
rect 64203 34376 64245 34385
rect 64587 34376 64629 34385
rect 64203 34336 64204 34376
rect 64244 34336 64245 34376
rect 64203 34327 64245 34336
rect 64396 34336 64588 34376
rect 64628 34336 64629 34376
rect 64204 34242 64244 34327
rect 62763 34208 62805 34217
rect 62763 34168 62764 34208
rect 62804 34168 62805 34208
rect 62763 34159 62805 34168
rect 61515 34040 61557 34049
rect 61515 34000 61516 34040
rect 61556 34000 61557 34040
rect 61515 33991 61557 34000
rect 62475 34040 62517 34049
rect 62475 34000 62476 34040
rect 62516 34000 62517 34040
rect 62475 33991 62517 34000
rect 61516 33713 61556 33991
rect 64396 33713 64436 34336
rect 64587 34327 64629 34336
rect 65452 34376 65492 35167
rect 68043 34544 68085 34553
rect 68043 34504 68044 34544
rect 68084 34504 68085 34544
rect 68043 34495 68085 34504
rect 65452 34327 65492 34336
rect 66315 34376 66357 34385
rect 66315 34336 66316 34376
rect 66356 34336 66357 34376
rect 66315 34327 66357 34336
rect 68044 34376 68084 34495
rect 68044 34327 68084 34336
rect 68907 34376 68949 34385
rect 68907 34336 68908 34376
rect 68948 34336 68949 34376
rect 68907 34327 68949 34336
rect 69292 34376 69332 37351
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 92427 36980 92469 36989
rect 92427 36940 92428 36980
rect 92468 36940 92469 36980
rect 92427 36931 92469 36940
rect 81579 36812 81621 36821
rect 81579 36772 81580 36812
rect 81620 36772 81621 36812
rect 81579 36763 81621 36772
rect 91024 36812 91066 36821
rect 91024 36772 91025 36812
rect 91065 36772 91066 36812
rect 91024 36763 91066 36772
rect 80427 36728 80469 36737
rect 80427 36688 80428 36728
rect 80468 36688 80469 36728
rect 80427 36679 80469 36688
rect 71979 36476 72021 36485
rect 71979 36436 71980 36476
rect 72020 36436 72021 36476
rect 71979 36427 72021 36436
rect 71980 36065 72020 36427
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 71403 36056 71445 36065
rect 71403 36016 71404 36056
rect 71444 36016 71445 36056
rect 71403 36007 71445 36016
rect 71979 36056 72021 36065
rect 71979 36016 71980 36056
rect 72020 36016 72021 36056
rect 71979 36007 72021 36016
rect 70156 35216 70196 35227
rect 70156 35141 70196 35176
rect 70155 35132 70197 35141
rect 70155 35092 70156 35132
rect 70196 35092 70197 35132
rect 70155 35083 70197 35092
rect 70923 35132 70965 35141
rect 70923 35092 70924 35132
rect 70964 35092 70965 35132
rect 70923 35083 70965 35092
rect 70924 34544 70964 35083
rect 70924 34495 70964 34504
rect 69292 34327 69332 34336
rect 70155 34376 70197 34385
rect 70155 34336 70156 34376
rect 70196 34336 70197 34376
rect 70155 34327 70197 34336
rect 70635 34376 70677 34385
rect 70635 34336 70636 34376
rect 70676 34336 70677 34376
rect 70635 34327 70677 34336
rect 66316 34242 66356 34327
rect 68908 34242 68948 34327
rect 70156 34242 70196 34327
rect 70636 34242 70676 34327
rect 64588 34208 64628 34217
rect 64588 33881 64628 34168
rect 68523 34208 68565 34217
rect 68523 34168 68524 34208
rect 68564 34168 68565 34208
rect 68523 34159 68565 34168
rect 68524 34074 68564 34159
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 64587 33872 64629 33881
rect 64587 33832 64588 33872
rect 64628 33832 64629 33872
rect 64587 33823 64629 33832
rect 61515 33704 61557 33713
rect 61515 33664 61516 33704
rect 61556 33664 61557 33704
rect 61515 33655 61557 33664
rect 64395 33704 64437 33713
rect 64395 33664 64396 33704
rect 64436 33664 64437 33704
rect 64395 33655 64437 33664
rect 55179 33620 55221 33629
rect 55179 33580 55180 33620
rect 55220 33580 55221 33620
rect 55179 33571 55221 33580
rect 52972 31732 53025 31772
rect 50379 31723 50421 31732
rect 52985 31374 53025 31732
rect 53791 31732 53876 31772
rect 53791 31374 53831 31732
rect 18617 7220 18657 7434
rect 20537 7220 20577 7434
rect 22841 7220 22881 7434
rect 23225 7220 23265 7434
rect 23417 7220 23457 7434
rect 18604 7180 18657 7220
rect 20524 7180 20577 7220
rect 22732 7180 22881 7220
rect 23212 7180 23265 7220
rect 23308 7180 23457 7220
rect 23644 7220 23684 7421
rect 23801 7220 23841 7434
rect 23993 7220 24033 7434
rect 25721 7220 25761 7434
rect 25913 7220 25953 7434
rect 26332 7253 26372 7421
rect 23644 7180 23732 7220
rect 17451 6824 17493 6833
rect 17451 6784 17452 6824
rect 17492 6784 17493 6824
rect 17451 6775 17493 6784
rect 17452 4892 17492 6775
rect 18604 5480 18644 7180
rect 18699 5648 18741 5657
rect 18699 5608 18700 5648
rect 18740 5608 18741 5648
rect 18699 5599 18741 5608
rect 17548 5440 18644 5480
rect 17548 5060 17588 5440
rect 17931 5312 17973 5321
rect 17931 5272 17932 5312
rect 17972 5272 17973 5312
rect 17931 5263 17973 5272
rect 17548 5011 17588 5020
rect 17644 4976 17684 4985
rect 17644 4892 17684 4936
rect 17932 4976 17972 5263
rect 18316 4976 18356 4985
rect 17972 4936 18316 4976
rect 17932 4927 17972 4936
rect 17452 4852 17684 4892
rect 18316 4733 18356 4936
rect 18604 4976 18644 5440
rect 18700 5405 18740 5599
rect 18699 5396 18741 5405
rect 18699 5356 18700 5396
rect 18740 5356 18741 5396
rect 18699 5347 18741 5356
rect 18700 5060 18740 5347
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 18700 5011 18740 5020
rect 18315 4724 18357 4733
rect 17260 4682 17300 4691
rect 18315 4684 18316 4724
rect 18356 4684 18357 4724
rect 18604 4724 18644 4936
rect 19180 4976 19220 4985
rect 18988 4808 19028 4817
rect 19180 4808 19220 4936
rect 19028 4768 19220 4808
rect 19564 4976 19604 4985
rect 18988 4759 19028 4768
rect 18604 4684 18740 4724
rect 18315 4675 18357 4684
rect 17260 4388 17300 4642
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 16876 4348 17300 4388
rect 16876 4136 16916 4348
rect 18700 4229 18740 4684
rect 18507 4220 18549 4229
rect 18507 4180 18508 4220
rect 18548 4180 18549 4220
rect 18507 4171 18549 4180
rect 18699 4220 18741 4229
rect 18699 4180 18700 4220
rect 18740 4180 18741 4220
rect 18699 4171 18741 4180
rect 19275 4220 19317 4229
rect 19275 4180 19276 4220
rect 19316 4180 19317 4220
rect 19275 4171 19317 4180
rect 18123 4136 18165 4145
rect 16876 4087 16916 4096
rect 17260 4123 17300 4132
rect 18123 4096 18124 4136
rect 18164 4096 18165 4136
rect 18123 4087 18165 4096
rect 17260 3977 17300 4083
rect 17355 4052 17397 4061
rect 17355 4012 17356 4052
rect 17396 4012 17397 4052
rect 17355 4003 17397 4012
rect 17259 3968 17301 3977
rect 17259 3928 17260 3968
rect 17300 3928 17301 3968
rect 17259 3919 17301 3928
rect 17356 3725 17396 4003
rect 18124 4002 18164 4087
rect 18508 3977 18548 4171
rect 19276 4086 19316 4171
rect 19564 4061 19604 4936
rect 20428 4976 20468 4985
rect 20428 4145 20468 4936
rect 20427 4136 20469 4145
rect 20427 4096 20428 4136
rect 20468 4096 20469 4136
rect 20427 4087 20469 4096
rect 19563 4052 19605 4061
rect 19563 4012 19564 4052
rect 19604 4012 19605 4052
rect 19563 4003 19605 4012
rect 18507 3968 18549 3977
rect 18507 3928 18508 3968
rect 18548 3928 18549 3968
rect 18507 3919 18549 3928
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 17355 3716 17397 3725
rect 17355 3676 17356 3716
rect 17396 3676 17397 3716
rect 17355 3667 17397 3676
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 8331 2876 8373 2885
rect 8331 2836 8332 2876
rect 8372 2836 8373 2876
rect 8331 2827 8373 2836
rect 20524 2717 20564 7180
rect 21579 5648 21621 5657
rect 21579 5608 21580 5648
rect 21620 5608 21621 5648
rect 21579 5599 21621 5608
rect 21580 5144 21620 5599
rect 21580 5095 21620 5104
rect 22444 4892 22484 4901
rect 21099 4724 21141 4733
rect 21099 4684 21100 4724
rect 21140 4684 21141 4724
rect 21099 4675 21141 4684
rect 21100 4304 21140 4675
rect 21140 4264 21236 4304
rect 21100 4255 21140 4264
rect 20907 4220 20949 4229
rect 20907 4180 20908 4220
rect 20948 4180 20949 4220
rect 20907 4171 20949 4180
rect 20715 4052 20757 4061
rect 20715 4012 20716 4052
rect 20756 4012 20757 4052
rect 20715 4003 20757 4012
rect 20619 2792 20661 2801
rect 20619 2752 20620 2792
rect 20660 2752 20661 2792
rect 20619 2743 20661 2752
rect 20523 2708 20565 2717
rect 20523 2668 20524 2708
rect 20564 2668 20565 2708
rect 20523 2659 20565 2668
rect 20332 2540 20372 2549
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 20332 1784 20372 2500
rect 20524 1868 20564 2659
rect 20620 2036 20660 2743
rect 20716 2624 20756 4003
rect 20908 3977 20948 4171
rect 20907 3968 20949 3977
rect 20907 3928 20908 3968
rect 20948 3928 20949 3968
rect 20907 3919 20949 3928
rect 21196 3464 21236 4264
rect 22444 4229 22484 4852
rect 22636 4724 22676 4735
rect 22636 4649 22676 4684
rect 22635 4640 22677 4649
rect 22635 4600 22636 4640
rect 22676 4600 22677 4640
rect 22635 4591 22677 4600
rect 22443 4220 22485 4229
rect 22443 4180 22444 4220
rect 22484 4180 22485 4220
rect 22443 4171 22485 4180
rect 21676 4136 21716 4147
rect 21676 4061 21716 4096
rect 21771 4136 21813 4145
rect 21771 4096 21772 4136
rect 21812 4096 21813 4136
rect 21771 4087 21813 4096
rect 20716 2575 20756 2584
rect 21004 3424 21196 3464
rect 20620 1987 20660 1996
rect 20716 1952 20756 1961
rect 20716 1868 20756 1912
rect 21004 1952 21044 3424
rect 21196 3415 21236 3424
rect 21292 4052 21332 4061
rect 21292 3305 21332 4012
rect 21675 4052 21717 4061
rect 21675 4012 21676 4052
rect 21716 4012 21717 4052
rect 21675 4003 21717 4012
rect 21579 3968 21621 3977
rect 21579 3928 21580 3968
rect 21620 3928 21621 3968
rect 21579 3919 21621 3928
rect 21580 3548 21620 3919
rect 21580 3499 21620 3508
rect 21484 3464 21524 3473
rect 21291 3296 21333 3305
rect 21291 3256 21292 3296
rect 21332 3256 21333 3296
rect 21291 3247 21333 3256
rect 21484 2801 21524 3424
rect 21483 2792 21525 2801
rect 21483 2752 21484 2792
rect 21524 2752 21525 2792
rect 21483 2743 21525 2752
rect 21580 2624 21620 2633
rect 21772 2624 21812 4087
rect 22444 3725 22484 4171
rect 22539 4136 22581 4145
rect 22539 4096 22540 4136
rect 22580 4096 22581 4136
rect 22539 4087 22581 4096
rect 22540 4002 22580 4087
rect 22443 3716 22485 3725
rect 22443 3676 22444 3716
rect 22484 3676 22485 3716
rect 22443 3667 22485 3676
rect 21867 3296 21909 3305
rect 21867 3256 21868 3296
rect 21908 3256 21909 3296
rect 21867 3247 21909 3256
rect 21868 3162 21908 3247
rect 22732 2876 22772 7180
rect 22924 4976 22964 4985
rect 22924 4649 22964 4936
rect 23212 4976 23252 7180
rect 23308 5237 23348 7180
rect 23692 5321 23732 7180
rect 23788 7180 23841 7220
rect 23980 7180 24033 7220
rect 25708 7180 25761 7220
rect 25900 7180 25953 7220
rect 26331 7244 26373 7253
rect 26331 7204 26332 7244
rect 26372 7204 26373 7244
rect 26331 7195 26373 7204
rect 31708 7220 31748 7421
rect 33785 7220 33825 7434
rect 31708 7180 31988 7220
rect 23788 7001 23828 7180
rect 23787 6992 23829 7001
rect 23787 6952 23788 6992
rect 23828 6952 23829 6992
rect 23787 6943 23829 6952
rect 23980 5657 24020 7180
rect 25611 7160 25653 7169
rect 25708 7160 25748 7180
rect 25611 7120 25612 7160
rect 25652 7120 25748 7160
rect 25611 7111 25653 7120
rect 23979 5648 24021 5657
rect 23979 5608 23980 5648
rect 24020 5608 24021 5648
rect 23979 5599 24021 5608
rect 23691 5312 23733 5321
rect 23691 5272 23692 5312
rect 23732 5272 23733 5312
rect 23691 5263 23733 5272
rect 24651 5312 24693 5321
rect 24651 5272 24652 5312
rect 24692 5272 24693 5312
rect 24651 5263 24693 5272
rect 23307 5228 23349 5237
rect 23307 5188 23308 5228
rect 23348 5188 23349 5228
rect 23307 5179 23349 5188
rect 23308 5060 23348 5179
rect 23308 5011 23348 5020
rect 24652 5060 24692 5263
rect 24747 5228 24789 5237
rect 25900 5228 25940 7180
rect 31755 6488 31797 6497
rect 31755 6448 31756 6488
rect 31796 6448 31797 6488
rect 31755 6439 31797 6448
rect 29259 5732 29301 5741
rect 29259 5692 29260 5732
rect 29300 5692 29301 5732
rect 29259 5683 29301 5692
rect 26283 5396 26325 5405
rect 26283 5356 26284 5396
rect 26324 5356 26325 5396
rect 26283 5347 26325 5356
rect 24747 5188 24748 5228
rect 24788 5188 24789 5228
rect 24747 5179 24789 5188
rect 25708 5188 25940 5228
rect 22923 4640 22965 4649
rect 22923 4600 22924 4640
rect 22964 4600 22965 4640
rect 22923 4591 22965 4600
rect 23212 3977 23252 4936
rect 23596 4724 23636 4733
rect 23308 4684 23596 4724
rect 23211 3968 23253 3977
rect 23211 3928 23212 3968
rect 23252 3928 23253 3968
rect 23211 3919 23253 3928
rect 23308 3548 23348 4684
rect 23596 4675 23636 4684
rect 24363 4724 24405 4733
rect 24363 4684 24364 4724
rect 24404 4684 24405 4724
rect 24363 4675 24405 4684
rect 24364 4590 24404 4675
rect 24652 4229 24692 5020
rect 24748 4976 24788 5179
rect 25708 5144 25748 5188
rect 25708 5095 25748 5104
rect 25036 4976 25076 4985
rect 24788 4936 24884 4976
rect 24748 4927 24788 4936
rect 24747 4724 24789 4733
rect 24747 4684 24748 4724
rect 24788 4684 24789 4724
rect 24747 4675 24789 4684
rect 24651 4220 24693 4229
rect 24651 4180 24652 4220
rect 24692 4180 24693 4220
rect 24651 4171 24693 4180
rect 24748 4136 24788 4675
rect 24844 4565 24884 4936
rect 25036 4649 25076 4936
rect 25900 4892 25940 4901
rect 25708 4724 25748 4733
rect 25612 4684 25708 4724
rect 25900 4724 25940 4852
rect 26284 4892 26324 5347
rect 26092 4724 26132 4733
rect 25900 4684 26092 4724
rect 25035 4640 25077 4649
rect 25035 4600 25036 4640
rect 25076 4600 25077 4640
rect 25035 4591 25077 4600
rect 24843 4556 24885 4565
rect 24843 4516 24844 4556
rect 24884 4516 24885 4556
rect 24843 4507 24885 4516
rect 24748 4087 24788 4096
rect 23691 3968 23733 3977
rect 23691 3928 23692 3968
rect 23732 3928 23733 3968
rect 23691 3919 23733 3928
rect 23692 3834 23732 3919
rect 23308 3499 23348 3508
rect 23691 3548 23733 3557
rect 23691 3508 23692 3548
rect 23732 3508 23733 3548
rect 23691 3499 23733 3508
rect 23692 3464 23732 3499
rect 23692 3413 23732 3424
rect 24555 3464 24597 3473
rect 24555 3424 24556 3464
rect 24596 3424 24692 3464
rect 24555 3415 24597 3424
rect 24556 3330 24596 3415
rect 22732 2801 22772 2836
rect 22731 2792 22773 2801
rect 22731 2752 22732 2792
rect 22772 2752 22773 2792
rect 22731 2743 22773 2752
rect 22732 2712 22772 2743
rect 23499 2708 23541 2717
rect 23499 2668 23500 2708
rect 23540 2668 23541 2708
rect 23499 2659 23541 2668
rect 24267 2708 24309 2717
rect 24267 2668 24268 2708
rect 24308 2668 24309 2708
rect 24267 2659 24309 2668
rect 21620 2584 21812 2624
rect 21580 2575 21620 2584
rect 23500 2574 23540 2659
rect 24268 2036 24308 2659
rect 24652 2624 24692 3424
rect 24652 2575 24692 2584
rect 25036 2045 25076 4591
rect 25612 4145 25652 4684
rect 25708 4675 25748 4684
rect 25707 4556 25749 4565
rect 25707 4516 25708 4556
rect 25748 4516 25749 4556
rect 25707 4507 25749 4516
rect 25131 4136 25173 4145
rect 25611 4136 25653 4145
rect 25131 4096 25132 4136
rect 25172 4096 25173 4136
rect 25131 4087 25173 4096
rect 25516 4096 25612 4136
rect 25652 4096 25653 4136
rect 25132 4002 25172 4087
rect 25516 3557 25556 4096
rect 25611 4087 25653 4096
rect 25708 3632 25748 4507
rect 25708 3583 25748 3592
rect 25996 4136 26036 4145
rect 25515 3548 25557 3557
rect 25515 3508 25516 3548
rect 25556 3508 25557 3548
rect 25515 3499 25557 3508
rect 25516 2624 25556 3499
rect 25996 2885 26036 4096
rect 25995 2876 26037 2885
rect 25995 2836 25996 2876
rect 26036 2836 26037 2876
rect 25995 2827 26037 2836
rect 25516 2575 25556 2584
rect 25900 2540 25940 2549
rect 24268 1987 24308 1996
rect 24651 2036 24693 2045
rect 24651 1996 24652 2036
rect 24692 1996 24693 2036
rect 24651 1987 24693 1996
rect 25035 2036 25077 2045
rect 25035 1996 25036 2036
rect 25076 1996 25077 2036
rect 25035 1987 25077 1996
rect 21004 1903 21044 1912
rect 24363 1952 24405 1961
rect 24363 1912 24364 1952
rect 24404 1912 24405 1952
rect 24363 1903 24405 1912
rect 24652 1952 24692 1987
rect 20524 1828 20756 1868
rect 24364 1818 24404 1903
rect 24652 1901 24692 1912
rect 25900 1793 25940 2500
rect 26092 1877 26132 4684
rect 26284 4649 26324 4852
rect 26283 4640 26325 4649
rect 26283 4600 26284 4640
rect 26324 4600 26325 4640
rect 26283 4591 26325 4600
rect 27147 4220 27189 4229
rect 27147 4180 27148 4220
rect 27188 4180 27189 4220
rect 27147 4171 27189 4180
rect 27435 4220 27477 4229
rect 27435 4180 27436 4220
rect 27476 4180 27477 4220
rect 27435 4171 27477 4180
rect 27148 4086 27188 4171
rect 27340 4052 27380 4061
rect 27244 4012 27340 4052
rect 27244 3716 27284 4012
rect 27340 3984 27380 4012
rect 27436 3884 27476 4171
rect 27723 4136 27765 4145
rect 27723 4096 27724 4136
rect 27764 4096 27765 4136
rect 27723 4087 27765 4096
rect 28588 4136 28628 4145
rect 26956 3676 27284 3716
rect 27340 3844 27476 3884
rect 26956 3296 26996 3676
rect 27243 3548 27285 3557
rect 27243 3508 27244 3548
rect 27284 3508 27285 3548
rect 27243 3499 27285 3508
rect 27244 3414 27284 3499
rect 27340 3491 27380 3844
rect 27340 3442 27380 3451
rect 27628 3464 27668 3473
rect 26956 3247 26996 3256
rect 27243 2960 27285 2969
rect 27243 2920 27244 2960
rect 27284 2920 27285 2960
rect 27243 2911 27285 2920
rect 27147 2624 27189 2633
rect 27147 2584 27148 2624
rect 27188 2584 27189 2624
rect 27147 2575 27189 2584
rect 27148 2045 27188 2575
rect 27147 2036 27189 2045
rect 27147 1996 27148 2036
rect 27188 1996 27189 2036
rect 27147 1987 27189 1996
rect 26860 1952 26900 1961
rect 26091 1868 26133 1877
rect 26091 1828 26092 1868
rect 26132 1828 26133 1868
rect 26091 1819 26133 1828
rect 20332 1735 20372 1744
rect 23979 1784 24021 1793
rect 23979 1744 23980 1784
rect 24020 1744 24021 1784
rect 23979 1735 24021 1744
rect 25899 1784 25941 1793
rect 25899 1744 25900 1784
rect 25940 1744 25941 1784
rect 25899 1735 25941 1744
rect 23980 1650 24020 1735
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 26668 1364 26708 1373
rect 26860 1364 26900 1912
rect 26955 1952 26997 1961
rect 26955 1912 26956 1952
rect 26996 1912 26997 1952
rect 26955 1903 26997 1912
rect 26956 1709 26996 1903
rect 26955 1700 26997 1709
rect 26955 1660 26956 1700
rect 26996 1660 26997 1700
rect 26955 1651 26997 1660
rect 26708 1324 26900 1364
rect 26668 1315 26708 1324
rect 26956 1112 26996 1651
rect 27148 1448 27188 1987
rect 27244 1952 27284 2911
rect 27628 2633 27668 3424
rect 27724 2969 27764 4087
rect 28588 3473 28628 4096
rect 28587 3464 28629 3473
rect 28587 3424 28588 3464
rect 28628 3424 28629 3464
rect 28587 3415 28629 3424
rect 27723 2960 27765 2969
rect 27723 2920 27724 2960
rect 27764 2920 27765 2960
rect 27723 2911 27765 2920
rect 28107 2876 28149 2885
rect 28107 2836 28108 2876
rect 28148 2836 28149 2876
rect 28107 2827 28149 2836
rect 27627 2624 27669 2633
rect 27627 2584 27628 2624
rect 27668 2584 27669 2624
rect 27627 2575 27669 2584
rect 28011 2624 28053 2633
rect 28011 2584 28012 2624
rect 28052 2584 28053 2624
rect 28011 2575 28053 2584
rect 28012 2490 28052 2575
rect 28108 2045 28148 2827
rect 28300 2624 28340 2633
rect 28107 2036 28149 2045
rect 28107 1996 28108 2036
rect 28148 1996 28149 2036
rect 28107 1987 28149 1996
rect 27244 1903 27284 1912
rect 28108 1952 28148 1987
rect 28108 1901 28148 1912
rect 28300 1709 28340 2584
rect 28396 2540 28436 2549
rect 28299 1700 28341 1709
rect 28299 1660 28300 1700
rect 28340 1660 28341 1700
rect 28299 1651 28341 1660
rect 27148 1408 27380 1448
rect 27340 1129 27380 1408
rect 28396 1373 28436 2500
rect 28588 1961 28628 3415
rect 28779 2960 28821 2969
rect 28779 2920 28780 2960
rect 28820 2920 28821 2960
rect 28779 2911 28821 2920
rect 28684 2792 28724 2801
rect 28587 1952 28629 1961
rect 28587 1912 28588 1952
rect 28628 1912 28629 1952
rect 28587 1903 28629 1912
rect 28395 1364 28437 1373
rect 26956 1063 26996 1072
rect 27052 1112 27092 1121
rect 27340 1080 27380 1089
rect 28300 1324 28396 1364
rect 28436 1324 28437 1364
rect 27052 953 27092 1072
rect 28300 953 28340 1324
rect 28395 1315 28437 1324
rect 28396 1112 28436 1121
rect 28684 1112 28724 2752
rect 28436 1072 28724 1112
rect 28780 1112 28820 2911
rect 29260 2120 29300 5683
rect 31756 5060 31796 6439
rect 31756 5011 31796 5020
rect 31660 4976 31700 4985
rect 31660 4397 31700 4936
rect 31852 4976 31892 4985
rect 31659 4388 31701 4397
rect 31659 4348 31660 4388
rect 31700 4348 31701 4388
rect 31659 4339 31701 4348
rect 31852 4304 31892 4936
rect 31852 4255 31892 4264
rect 31756 4220 31796 4229
rect 29932 4136 29972 4147
rect 29932 4061 29972 4096
rect 31180 4136 31220 4145
rect 29931 4052 29973 4061
rect 29931 4012 29932 4052
rect 29972 4012 29973 4052
rect 29931 4003 29973 4012
rect 29740 3968 29780 3979
rect 29740 3893 29780 3928
rect 29739 3884 29781 3893
rect 29739 3844 29740 3884
rect 29780 3844 29781 3884
rect 29739 3835 29781 3844
rect 29740 3557 29780 3835
rect 29739 3548 29781 3557
rect 29739 3508 29740 3548
rect 29780 3508 29781 3548
rect 29739 3499 29781 3508
rect 31180 3221 31220 4096
rect 31660 4136 31700 4145
rect 31372 4052 31412 4061
rect 31660 4052 31700 4096
rect 31412 4012 31700 4052
rect 31276 3464 31316 3473
rect 31372 3464 31412 4012
rect 31756 3977 31796 4180
rect 31948 4220 31988 7180
rect 33772 7180 33825 7220
rect 34012 7220 34052 7421
rect 34361 7220 34401 7434
rect 34012 7180 34100 7220
rect 33772 7085 33812 7180
rect 33771 7076 33813 7085
rect 33771 7036 33772 7076
rect 33812 7036 33813 7076
rect 33771 7027 33813 7036
rect 33387 6824 33429 6833
rect 33387 6784 33388 6824
rect 33428 6784 33429 6824
rect 33387 6775 33429 6784
rect 32715 5396 32757 5405
rect 32715 5356 32716 5396
rect 32756 5356 32757 5396
rect 32715 5347 32757 5356
rect 32716 4976 32756 5347
rect 32716 4927 32756 4936
rect 32908 4976 32948 4985
rect 32908 4817 32948 4936
rect 33100 4976 33140 4985
rect 32715 4808 32757 4817
rect 32812 4808 32852 4817
rect 32715 4768 32716 4808
rect 32756 4768 32812 4808
rect 32715 4759 32757 4768
rect 32812 4759 32852 4768
rect 32907 4808 32949 4817
rect 32907 4768 32908 4808
rect 32948 4768 32949 4808
rect 32907 4759 32949 4768
rect 32043 4724 32085 4733
rect 32043 4684 32044 4724
rect 32084 4684 32085 4724
rect 32043 4675 32085 4684
rect 32427 4724 32469 4733
rect 32427 4684 32428 4724
rect 32468 4684 32469 4724
rect 32427 4675 32469 4684
rect 31948 4171 31988 4180
rect 32044 4136 32084 4675
rect 32139 4388 32181 4397
rect 32139 4348 32140 4388
rect 32180 4348 32181 4388
rect 32139 4339 32181 4348
rect 32044 4087 32084 4096
rect 31755 3968 31797 3977
rect 31755 3928 31756 3968
rect 31796 3928 31797 3968
rect 31755 3919 31797 3928
rect 32140 3473 32180 4339
rect 32428 4304 32468 4675
rect 32428 4255 32468 4264
rect 33100 4145 33140 4936
rect 33196 4892 33236 4901
rect 32619 4136 32661 4145
rect 32619 4096 32620 4136
rect 32660 4096 32661 4136
rect 32619 4087 32661 4096
rect 33099 4136 33141 4145
rect 33099 4096 33100 4136
rect 33140 4096 33141 4136
rect 33099 4087 33141 4096
rect 32620 4002 32660 4087
rect 32716 3968 32756 3977
rect 32716 3800 32756 3928
rect 32620 3760 32756 3800
rect 32235 3716 32277 3725
rect 32235 3676 32236 3716
rect 32276 3676 32277 3716
rect 32235 3667 32277 3676
rect 31316 3424 31412 3464
rect 32139 3464 32181 3473
rect 32139 3424 32140 3464
rect 32180 3424 32181 3464
rect 31276 3415 31316 3424
rect 32139 3415 32181 3424
rect 30411 3212 30453 3221
rect 30411 3172 30412 3212
rect 30452 3172 30453 3212
rect 30411 3163 30453 3172
rect 31179 3212 31221 3221
rect 31179 3172 31180 3212
rect 31220 3172 31221 3212
rect 31179 3163 31221 3172
rect 30028 2792 30068 2801
rect 29260 1793 29300 2080
rect 29644 2752 30028 2792
rect 29644 2036 29684 2752
rect 30028 2743 30068 2752
rect 30412 2624 30452 3163
rect 32236 2708 32276 3667
rect 32236 2659 32276 2668
rect 32524 3464 32564 3473
rect 30412 2575 30452 2584
rect 30699 2624 30741 2633
rect 30699 2584 30700 2624
rect 30740 2584 30741 2624
rect 30699 2575 30741 2584
rect 30316 2540 30356 2549
rect 30316 2129 30356 2500
rect 30700 2490 30740 2575
rect 32428 2456 32468 2465
rect 30315 2120 30357 2129
rect 30315 2080 30316 2120
rect 30356 2080 30357 2120
rect 30315 2071 30357 2080
rect 32043 2120 32085 2129
rect 32043 2080 32044 2120
rect 32084 2080 32085 2120
rect 32043 2071 32085 2080
rect 29644 1987 29684 1996
rect 29739 2036 29781 2045
rect 29739 1996 29740 2036
rect 29780 1996 29781 2036
rect 29739 1987 29781 1996
rect 30891 2036 30933 2045
rect 30891 1996 30892 2036
rect 30932 1996 30933 2036
rect 30891 1987 30933 1996
rect 29259 1784 29301 1793
rect 29259 1744 29260 1784
rect 29300 1744 29301 1784
rect 29259 1735 29301 1744
rect 28396 1063 28436 1072
rect 28780 1063 28820 1072
rect 29644 1112 29684 1121
rect 29740 1112 29780 1987
rect 30028 1952 30068 1963
rect 30028 1877 30068 1912
rect 30892 1952 30932 1987
rect 32044 1986 32084 2071
rect 30892 1901 30932 1912
rect 32236 1952 32276 1961
rect 30027 1868 30069 1877
rect 30027 1828 30028 1868
rect 30068 1828 30069 1868
rect 30027 1819 30069 1828
rect 30795 1364 30837 1373
rect 30795 1324 30796 1364
rect 30836 1324 30837 1364
rect 30795 1315 30837 1324
rect 32044 1364 32084 1373
rect 32236 1364 32276 1912
rect 32428 1868 32468 2416
rect 32524 2129 32564 3424
rect 32620 3389 32660 3760
rect 33100 3641 33140 4087
rect 33196 3977 33236 4852
rect 33292 4817 33332 4902
rect 33388 4892 33428 6775
rect 33388 4843 33428 4852
rect 33484 4976 33524 4985
rect 33484 4817 33524 4936
rect 33291 4808 33333 4817
rect 33291 4768 33292 4808
rect 33332 4768 33333 4808
rect 33291 4759 33333 4768
rect 33483 4808 33525 4817
rect 33483 4768 33484 4808
rect 33524 4768 33525 4808
rect 33483 4759 33525 4768
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 33195 3968 33237 3977
rect 33195 3928 33196 3968
rect 33236 3928 33237 3968
rect 33195 3919 33237 3928
rect 32715 3632 32757 3641
rect 32715 3592 32716 3632
rect 32756 3592 32757 3632
rect 32715 3583 32757 3592
rect 33099 3632 33141 3641
rect 33099 3592 33100 3632
rect 33140 3592 33141 3632
rect 33099 3583 33141 3592
rect 32716 3498 32756 3583
rect 33484 3464 33524 3473
rect 33196 3424 33484 3464
rect 32619 3380 32661 3389
rect 32619 3340 32620 3380
rect 32660 3340 32661 3380
rect 32619 3331 32661 3340
rect 32619 2960 32661 2969
rect 32619 2920 32620 2960
rect 32660 2920 32661 2960
rect 32619 2911 32661 2920
rect 32523 2120 32565 2129
rect 32523 2080 32524 2120
rect 32564 2080 32565 2120
rect 32523 2071 32565 2080
rect 32620 1952 32660 2911
rect 33196 2633 33236 3424
rect 33484 3415 33524 3424
rect 33772 3464 33812 7027
rect 34060 3641 34100 7180
rect 34348 7180 34401 7220
rect 34588 7220 34628 7421
rect 34745 7220 34785 7434
rect 34937 7220 34977 7434
rect 34588 7180 34676 7220
rect 34059 3632 34101 3641
rect 34059 3592 34060 3632
rect 34100 3592 34101 3632
rect 34059 3583 34101 3592
rect 34348 3557 34388 7180
rect 34636 5657 34676 7180
rect 34732 7180 34785 7220
rect 34924 7180 34977 7220
rect 35164 7220 35204 7421
rect 35356 7220 35396 7421
rect 35513 7220 35553 7434
rect 36665 7220 36705 7434
rect 35164 7180 35252 7220
rect 35356 7180 35444 7220
rect 34635 5648 34677 5657
rect 34635 5608 34636 5648
rect 34676 5608 34677 5648
rect 34635 5599 34677 5608
rect 34732 5480 34772 7180
rect 34924 5741 34964 7180
rect 34923 5732 34965 5741
rect 34923 5692 34924 5732
rect 34964 5692 34965 5732
rect 34923 5683 34965 5692
rect 35019 5648 35061 5657
rect 35019 5608 35020 5648
rect 35060 5608 35061 5648
rect 35019 5599 35061 5608
rect 34444 5440 34772 5480
rect 34444 5144 34484 5440
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 35020 5144 35060 5599
rect 35115 5564 35157 5573
rect 35115 5524 35116 5564
rect 35156 5524 35157 5564
rect 35115 5515 35157 5524
rect 34444 5104 34580 5144
rect 34443 4808 34485 4817
rect 34443 4768 34444 4808
rect 34484 4768 34485 4808
rect 34443 4759 34485 4768
rect 34444 4397 34484 4759
rect 34443 4388 34485 4397
rect 34443 4348 34444 4388
rect 34484 4348 34485 4388
rect 34443 4339 34485 4348
rect 34444 4052 34484 4339
rect 34540 4229 34580 5104
rect 34924 5104 35060 5144
rect 34635 4472 34677 4481
rect 34635 4432 34636 4472
rect 34676 4432 34677 4472
rect 34924 4472 34964 5104
rect 35020 4976 35060 4985
rect 35020 4817 35060 4936
rect 35116 4976 35156 5515
rect 35212 5321 35252 7180
rect 35404 5825 35444 7180
rect 35500 7180 35553 7220
rect 36652 7180 36705 7220
rect 37468 7220 37508 7421
rect 37625 7220 37665 7434
rect 39545 7220 39585 7434
rect 39737 7220 39777 7434
rect 39929 7220 39969 7434
rect 40121 7220 40161 7434
rect 37468 7180 37556 7220
rect 35403 5816 35445 5825
rect 35403 5776 35404 5816
rect 35444 5776 35445 5816
rect 35403 5767 35445 5776
rect 35500 5648 35540 7180
rect 36171 6572 36213 6581
rect 36171 6532 36172 6572
rect 36212 6532 36213 6572
rect 36171 6523 36213 6532
rect 35308 5608 35540 5648
rect 35211 5312 35253 5321
rect 35211 5272 35212 5312
rect 35252 5272 35253 5312
rect 35211 5263 35253 5272
rect 35116 4927 35156 4936
rect 35212 4976 35252 4985
rect 35019 4808 35061 4817
rect 35019 4768 35020 4808
rect 35060 4768 35061 4808
rect 35019 4759 35061 4768
rect 35212 4733 35252 4936
rect 35211 4724 35253 4733
rect 35211 4684 35212 4724
rect 35252 4684 35253 4724
rect 35211 4675 35253 4684
rect 34924 4432 35060 4472
rect 34635 4423 34677 4432
rect 34539 4220 34581 4229
rect 34539 4180 34540 4220
rect 34580 4180 34581 4220
rect 34539 4171 34581 4180
rect 34636 4136 34676 4423
rect 34923 4304 34965 4313
rect 34923 4264 34924 4304
rect 34964 4264 34965 4304
rect 34923 4255 34965 4264
rect 34636 4087 34676 4096
rect 34732 4136 34772 4145
rect 34444 4012 34580 4052
rect 34540 3968 34580 4012
rect 34732 3968 34772 4096
rect 34827 4136 34869 4145
rect 34827 4096 34828 4136
rect 34868 4096 34869 4136
rect 34827 4087 34869 4096
rect 34924 4136 34964 4255
rect 34924 4087 34964 4096
rect 34828 4002 34868 4087
rect 34540 3928 34772 3968
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 33867 3548 33909 3557
rect 33867 3508 33868 3548
rect 33908 3508 33909 3548
rect 33867 3499 33909 3508
rect 34347 3548 34389 3557
rect 34347 3508 34348 3548
rect 34388 3508 34389 3548
rect 34347 3499 34389 3508
rect 33772 3415 33812 3424
rect 33868 3414 33908 3499
rect 34156 3212 34196 3221
rect 33772 3172 34156 3212
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 33195 2624 33237 2633
rect 33195 2584 33196 2624
rect 33236 2584 33237 2624
rect 33195 2575 33237 2584
rect 33483 2624 33525 2633
rect 33483 2584 33484 2624
rect 33524 2584 33525 2624
rect 33483 2575 33525 2584
rect 33580 2624 33620 2633
rect 33772 2624 33812 3172
rect 34156 3163 34196 3172
rect 33620 2584 33812 2624
rect 33964 2624 34004 2633
rect 33580 2575 33620 2584
rect 33484 1961 33524 2575
rect 32620 1903 32660 1912
rect 33483 1952 33525 1961
rect 33483 1912 33484 1952
rect 33524 1912 33525 1952
rect 33483 1903 33525 1912
rect 32428 1828 32564 1868
rect 32331 1700 32373 1709
rect 32331 1660 32332 1700
rect 32372 1660 32373 1700
rect 32331 1651 32373 1660
rect 32084 1324 32276 1364
rect 32044 1315 32084 1324
rect 30796 1230 30836 1315
rect 29684 1072 29780 1112
rect 32332 1112 32372 1651
rect 29644 1063 29684 1072
rect 32332 1063 32372 1072
rect 32427 1112 32469 1121
rect 32427 1072 32428 1112
rect 32468 1072 32469 1112
rect 32427 1063 32469 1072
rect 32428 978 32468 1063
rect 32524 1037 32564 1828
rect 33484 1818 33524 1903
rect 33964 1877 34004 2584
rect 34827 2624 34869 2633
rect 34827 2584 34828 2624
rect 34868 2584 34869 2624
rect 34827 2575 34869 2584
rect 34828 2490 34868 2575
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 34635 2120 34677 2129
rect 34635 2080 34636 2120
rect 34676 2080 34677 2120
rect 34635 2071 34677 2080
rect 34924 2120 34964 2129
rect 35020 2120 35060 4432
rect 35115 4136 35157 4145
rect 35115 4096 35116 4136
rect 35156 4096 35157 4136
rect 35115 4087 35157 4096
rect 34964 2080 35060 2120
rect 34924 2071 34964 2080
rect 34636 1986 34676 2071
rect 33963 1868 34005 1877
rect 33963 1828 33964 1868
rect 34004 1828 34005 1868
rect 33963 1819 34005 1828
rect 34635 1700 34677 1709
rect 34635 1660 34636 1700
rect 34676 1660 34677 1700
rect 34635 1651 34677 1660
rect 34636 1566 34676 1651
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 34924 1112 34964 1123
rect 35020 1121 35060 2080
rect 35116 1373 35156 4087
rect 35308 2204 35348 5608
rect 35403 5480 35445 5489
rect 35403 5440 35404 5480
rect 35444 5440 35445 5480
rect 35403 5431 35445 5440
rect 35404 4976 35444 5431
rect 35787 5228 35829 5237
rect 35787 5188 35788 5228
rect 35828 5188 35924 5228
rect 35787 5179 35829 5188
rect 35884 5144 35924 5188
rect 35884 5095 35924 5104
rect 35979 5144 36021 5153
rect 35979 5104 35980 5144
rect 36020 5104 36021 5144
rect 35979 5095 36021 5104
rect 35404 4927 35444 4936
rect 35500 4976 35540 4985
rect 35500 4817 35540 4936
rect 35596 4976 35636 4985
rect 35499 4808 35541 4817
rect 35499 4768 35500 4808
rect 35540 4768 35541 4808
rect 35499 4759 35541 4768
rect 35596 4481 35636 4936
rect 35692 4976 35732 4985
rect 35980 4976 36020 5095
rect 35732 4936 36020 4976
rect 36076 4976 36116 4985
rect 35692 4927 35732 4936
rect 35595 4472 35637 4481
rect 35595 4432 35596 4472
rect 35636 4432 35637 4472
rect 35595 4423 35637 4432
rect 36076 4397 36116 4936
rect 36172 4976 36212 6523
rect 36212 4936 36308 4976
rect 36172 4927 36212 4936
rect 36075 4388 36117 4397
rect 36075 4348 36076 4388
rect 36116 4348 36117 4388
rect 36075 4339 36117 4348
rect 35595 4304 35637 4313
rect 35595 4264 35596 4304
rect 35636 4264 35637 4304
rect 35595 4255 35637 4264
rect 35788 4304 35828 4313
rect 36171 4304 36213 4313
rect 35828 4264 36020 4304
rect 35788 4255 35828 4264
rect 35403 4136 35445 4145
rect 35403 4096 35404 4136
rect 35444 4096 35445 4136
rect 35403 4087 35445 4096
rect 35596 4136 35636 4255
rect 35596 4087 35636 4096
rect 35788 4136 35828 4145
rect 35212 2164 35348 2204
rect 35212 1793 35252 2164
rect 35404 2129 35444 4087
rect 35788 3725 35828 4096
rect 35980 4136 36020 4264
rect 36171 4264 36172 4304
rect 36212 4264 36213 4304
rect 36171 4255 36213 4264
rect 35980 4087 36020 4096
rect 36172 4136 36212 4255
rect 36172 4087 36212 4096
rect 36268 4136 36308 4936
rect 36268 4087 36308 4096
rect 36075 4052 36117 4061
rect 36075 4012 36076 4052
rect 36116 4012 36117 4052
rect 36075 4003 36117 4012
rect 36076 3918 36116 4003
rect 36652 3884 36692 7180
rect 37516 7085 37556 7180
rect 37612 7180 37665 7220
rect 39532 7180 39585 7220
rect 39724 7180 39777 7220
rect 39916 7180 39969 7220
rect 40012 7180 40161 7220
rect 40348 7220 40388 7421
rect 40505 7220 40545 7434
rect 40348 7180 40436 7220
rect 37515 7076 37557 7085
rect 37515 7036 37516 7076
rect 37556 7036 37557 7076
rect 37515 7027 37557 7036
rect 37612 6833 37652 7180
rect 37899 7076 37941 7085
rect 37899 7036 37900 7076
rect 37940 7036 37941 7076
rect 37899 7027 37941 7036
rect 37611 6824 37653 6833
rect 37611 6784 37612 6824
rect 37652 6784 37653 6824
rect 37611 6775 37653 6784
rect 37611 6656 37653 6665
rect 37611 6616 37612 6656
rect 37652 6616 37653 6656
rect 37611 6607 37653 6616
rect 37612 4976 37652 6607
rect 37612 4927 37652 4936
rect 37708 4892 37748 4901
rect 36939 4808 36981 4817
rect 36939 4768 36940 4808
rect 36980 4768 36981 4808
rect 36939 4759 36981 4768
rect 36940 4304 36980 4759
rect 37708 4472 37748 4852
rect 37900 4892 37940 7027
rect 39435 5144 39477 5153
rect 39435 5104 39436 5144
rect 39476 5104 39477 5144
rect 39435 5095 39477 5104
rect 39436 5010 39476 5095
rect 37900 4843 37940 4852
rect 37996 4976 38036 4985
rect 37803 4808 37845 4817
rect 37803 4768 37804 4808
rect 37844 4768 37845 4808
rect 37803 4759 37845 4768
rect 37804 4674 37844 4759
rect 36940 4255 36980 4264
rect 37612 4432 37748 4472
rect 36844 4220 36884 4229
rect 36747 4136 36789 4145
rect 36747 4096 36748 4136
rect 36788 4096 36789 4136
rect 36747 4087 36789 4096
rect 36748 4002 36788 4087
rect 36844 4061 36884 4180
rect 37035 4220 37077 4229
rect 37035 4180 37036 4220
rect 37076 4180 37077 4220
rect 37035 4171 37077 4180
rect 37612 4220 37652 4432
rect 37036 4086 37076 4171
rect 37132 4136 37172 4145
rect 36843 4052 36885 4061
rect 36843 4012 36844 4052
rect 36884 4012 36885 4052
rect 36843 4003 36885 4012
rect 36652 3844 36788 3884
rect 35787 3716 35829 3725
rect 35787 3676 35788 3716
rect 35828 3676 35829 3716
rect 35787 3667 35829 3676
rect 35691 3632 35733 3641
rect 35691 3592 35692 3632
rect 35732 3592 35733 3632
rect 35691 3583 35733 3592
rect 35883 3632 35925 3641
rect 35883 3592 35884 3632
rect 35924 3592 35925 3632
rect 35883 3583 35925 3592
rect 35500 3464 35540 3473
rect 35403 2120 35445 2129
rect 35403 2080 35404 2120
rect 35444 2080 35445 2120
rect 35403 2071 35445 2080
rect 35211 1784 35253 1793
rect 35211 1744 35212 1784
rect 35252 1744 35253 1784
rect 35211 1735 35253 1744
rect 35115 1364 35157 1373
rect 35115 1324 35116 1364
rect 35156 1324 35157 1364
rect 35115 1315 35157 1324
rect 32734 1097 32774 1106
rect 32734 1037 32774 1057
rect 34924 1037 34964 1072
rect 35019 1112 35061 1121
rect 35019 1072 35020 1112
rect 35060 1072 35061 1112
rect 35019 1063 35061 1072
rect 35212 1112 35252 1735
rect 35212 1063 35252 1072
rect 35307 1112 35349 1121
rect 35307 1072 35308 1112
rect 35348 1072 35349 1112
rect 35307 1063 35349 1072
rect 32523 1028 32565 1037
rect 32523 988 32524 1028
rect 32564 988 32565 1028
rect 32523 979 32565 988
rect 32715 1028 32774 1037
rect 32715 988 32716 1028
rect 32756 988 32774 1028
rect 34923 1028 34965 1037
rect 34923 988 34924 1028
rect 34964 988 34965 1028
rect 32715 979 32757 988
rect 34923 979 34965 988
rect 35308 978 35348 1063
rect 35500 1037 35540 3424
rect 35692 3053 35732 3583
rect 35787 3548 35829 3557
rect 35787 3508 35788 3548
rect 35828 3508 35829 3548
rect 35787 3499 35829 3508
rect 35884 3548 35924 3583
rect 35788 3464 35828 3499
rect 35884 3497 35924 3508
rect 35788 3296 35828 3424
rect 35788 3256 36020 3296
rect 35691 3044 35733 3053
rect 35691 3004 35692 3044
rect 35732 3004 35733 3044
rect 35691 2995 35733 3004
rect 35980 2876 36020 3256
rect 36172 3212 36212 3221
rect 36212 3172 36692 3212
rect 36172 3163 36212 3172
rect 35980 2827 36020 2836
rect 36075 2624 36117 2633
rect 36075 2584 36076 2624
rect 36116 2584 36117 2624
rect 36075 2575 36117 2584
rect 36652 2624 36692 3172
rect 36652 2575 36692 2584
rect 36076 1952 36116 2575
rect 36076 1903 36116 1912
rect 36748 1457 36788 3844
rect 37132 3809 37172 4096
rect 37515 4136 37557 4145
rect 37515 4096 37516 4136
rect 37556 4096 37557 4136
rect 37515 4087 37557 4096
rect 37516 4002 37556 4087
rect 37612 4061 37652 4180
rect 37708 4136 37748 4145
rect 37611 4052 37653 4061
rect 37611 4012 37612 4052
rect 37652 4012 37653 4052
rect 37611 4003 37653 4012
rect 37708 3977 37748 4096
rect 37707 3968 37749 3977
rect 37707 3928 37708 3968
rect 37748 3928 37749 3968
rect 37707 3919 37749 3928
rect 37131 3800 37173 3809
rect 37131 3760 37132 3800
rect 37172 3760 37173 3800
rect 37131 3751 37173 3760
rect 37708 3389 37748 3919
rect 37996 3809 38036 4936
rect 39243 4808 39285 4817
rect 39243 4768 39244 4808
rect 39284 4768 39285 4808
rect 39243 4759 39285 4768
rect 39244 4674 39284 4759
rect 38859 4136 38901 4145
rect 38859 4096 38860 4136
rect 38900 4096 38901 4136
rect 38859 4087 38901 4096
rect 39148 4136 39188 4145
rect 38860 4002 38900 4087
rect 39148 3977 39188 4096
rect 39532 4052 39572 7180
rect 39436 4012 39572 4052
rect 39628 4962 39668 4971
rect 39052 3968 39092 3977
rect 39052 3809 39092 3928
rect 39147 3968 39189 3977
rect 39147 3928 39148 3968
rect 39188 3928 39189 3968
rect 39147 3919 39189 3928
rect 37995 3800 38037 3809
rect 37995 3760 37996 3800
rect 38036 3760 38037 3800
rect 37995 3751 38037 3760
rect 39051 3800 39093 3809
rect 39051 3760 39052 3800
rect 39092 3760 39093 3800
rect 39051 3751 39093 3760
rect 39052 3464 39092 3751
rect 39052 3415 39092 3424
rect 39147 3464 39189 3473
rect 39147 3424 39148 3464
rect 39188 3424 39189 3464
rect 39147 3415 39189 3424
rect 39244 3464 39284 3473
rect 37707 3380 37749 3389
rect 37707 3340 37708 3380
rect 37748 3340 37749 3380
rect 37707 3331 37749 3340
rect 39148 3330 39188 3415
rect 39051 3044 39093 3053
rect 39051 3004 39052 3044
rect 39092 3004 39093 3044
rect 39051 2995 39093 3004
rect 39052 2876 39092 2995
rect 39052 2827 39092 2836
rect 37036 2624 37076 2633
rect 36940 2584 37036 2624
rect 36940 1961 36980 2584
rect 37036 2575 37076 2584
rect 37899 2624 37941 2633
rect 37899 2584 37900 2624
rect 37940 2584 37941 2624
rect 37899 2575 37941 2584
rect 38859 2624 38901 2633
rect 38859 2584 38860 2624
rect 38900 2584 38901 2624
rect 38859 2575 38901 2584
rect 37900 2045 37940 2575
rect 38187 2540 38229 2549
rect 38187 2500 38188 2540
rect 38228 2500 38229 2540
rect 38187 2491 38229 2500
rect 37899 2036 37941 2045
rect 37899 1996 37900 2036
rect 37940 1996 37941 2036
rect 37899 1987 37941 1996
rect 36939 1957 36981 1961
rect 36939 1912 36940 1957
rect 36980 1912 36981 1957
rect 36939 1903 36981 1912
rect 37324 1952 37364 1961
rect 36747 1448 36789 1457
rect 36747 1408 36748 1448
rect 36788 1408 36789 1448
rect 36747 1399 36789 1408
rect 37324 1373 37364 1912
rect 37707 1700 37749 1709
rect 37707 1660 37708 1700
rect 37748 1660 37749 1700
rect 37707 1651 37749 1660
rect 37708 1566 37748 1651
rect 35595 1364 35637 1373
rect 35595 1324 35596 1364
rect 35636 1324 35637 1364
rect 35595 1315 35637 1324
rect 37323 1364 37365 1373
rect 37323 1324 37324 1364
rect 37364 1324 37365 1364
rect 37323 1315 37365 1324
rect 35596 1230 35636 1315
rect 38188 1112 38228 2491
rect 38860 1952 38900 2575
rect 38860 1903 38900 1912
rect 38571 1700 38613 1709
rect 38571 1660 38572 1700
rect 38612 1660 38613 1700
rect 38571 1651 38613 1660
rect 38188 1037 38228 1072
rect 38475 1112 38517 1121
rect 38475 1072 38476 1112
rect 38516 1072 38517 1112
rect 38475 1063 38517 1072
rect 38572 1112 38612 1651
rect 39244 1625 39284 3424
rect 39436 2717 39476 4012
rect 39628 3977 39668 4922
rect 39627 3968 39669 3977
rect 39627 3928 39628 3968
rect 39668 3928 39669 3968
rect 39627 3919 39669 3928
rect 39531 3884 39573 3893
rect 39531 3844 39532 3884
rect 39572 3844 39573 3884
rect 39531 3835 39573 3844
rect 39532 3473 39572 3835
rect 39531 3464 39573 3473
rect 39531 3424 39532 3464
rect 39572 3424 39573 3464
rect 39531 3415 39573 3424
rect 39628 3464 39668 3473
rect 39435 2708 39477 2717
rect 39435 2668 39436 2708
rect 39476 2668 39477 2708
rect 39435 2659 39477 2668
rect 39628 2549 39668 3424
rect 39724 2633 39764 7180
rect 39916 3632 39956 7180
rect 40012 4061 40052 7180
rect 40108 4976 40148 4985
rect 40011 4052 40053 4061
rect 40011 4012 40012 4052
rect 40052 4012 40053 4052
rect 40011 4003 40053 4012
rect 39820 3592 39956 3632
rect 39820 2960 39860 3592
rect 40012 3548 40052 4003
rect 40108 3725 40148 4936
rect 40107 3716 40149 3725
rect 40107 3676 40108 3716
rect 40148 3676 40149 3716
rect 40107 3667 40149 3676
rect 40396 3632 40436 7180
rect 40492 7180 40545 7220
rect 40732 7220 40772 7421
rect 40889 7337 40929 7434
rect 40888 7328 40930 7337
rect 40888 7288 40889 7328
rect 40929 7288 41012 7328
rect 40888 7279 40930 7288
rect 40732 7180 40820 7220
rect 40492 4229 40532 7180
rect 40780 6329 40820 7180
rect 40779 6320 40821 6329
rect 40779 6280 40780 6320
rect 40820 6280 40821 6320
rect 40779 6271 40821 6280
rect 40587 5480 40629 5489
rect 40587 5440 40588 5480
rect 40628 5440 40629 5480
rect 40587 5431 40629 5440
rect 40588 4976 40628 5431
rect 40588 4927 40628 4936
rect 40684 4892 40724 4901
rect 40684 4817 40724 4852
rect 40683 4808 40725 4817
rect 40683 4768 40684 4808
rect 40724 4768 40725 4808
rect 40683 4759 40725 4768
rect 40491 4220 40533 4229
rect 40491 4180 40492 4220
rect 40532 4180 40533 4220
rect 40491 4171 40533 4180
rect 40396 3592 40628 3632
rect 40012 3499 40052 3508
rect 39915 3464 39957 3473
rect 39915 3424 39916 3464
rect 39956 3424 39957 3464
rect 39915 3415 39957 3424
rect 40492 3464 40532 3473
rect 39916 3330 39956 3415
rect 40300 3296 40340 3305
rect 40492 3296 40532 3424
rect 40340 3256 40532 3296
rect 40300 3247 40340 3256
rect 39820 2920 40244 2960
rect 39723 2624 39765 2633
rect 39723 2584 39724 2624
rect 39764 2584 39765 2624
rect 39723 2575 39765 2584
rect 39820 2624 39860 2635
rect 39820 2549 39860 2584
rect 40107 2624 40149 2633
rect 40107 2584 40108 2624
rect 40148 2584 40149 2624
rect 40107 2575 40149 2584
rect 40204 2624 40244 2920
rect 39627 2540 39669 2549
rect 39627 2500 39628 2540
rect 39668 2500 39669 2540
rect 39627 2491 39669 2500
rect 39819 2540 39861 2549
rect 39819 2500 39820 2540
rect 39860 2500 39861 2540
rect 39819 2491 39861 2500
rect 40108 2490 40148 2575
rect 39724 1952 39764 1963
rect 39724 1877 39764 1912
rect 40108 1952 40148 1961
rect 39723 1868 39765 1877
rect 39723 1828 39724 1868
rect 39764 1828 39765 1868
rect 39723 1819 39765 1828
rect 39243 1616 39285 1625
rect 39243 1576 39244 1616
rect 39284 1576 39285 1616
rect 39243 1567 39285 1576
rect 40108 1373 40148 1912
rect 38859 1364 38901 1373
rect 38859 1324 38860 1364
rect 38900 1324 38901 1364
rect 38859 1315 38901 1324
rect 40107 1364 40149 1373
rect 40107 1324 40108 1364
rect 40148 1324 40149 1364
rect 40107 1315 40149 1324
rect 40204 1364 40244 2584
rect 38860 1230 38900 1315
rect 40204 1121 40244 1324
rect 40492 2792 40532 2801
rect 40492 1121 40532 2752
rect 40588 1961 40628 3592
rect 40587 1952 40629 1961
rect 40587 1912 40588 1952
rect 40628 1912 40629 1952
rect 40587 1903 40629 1912
rect 40684 1205 40724 4759
rect 40875 4640 40917 4649
rect 40875 4600 40876 4640
rect 40916 4600 40917 4640
rect 40875 4591 40917 4600
rect 40876 3977 40916 4591
rect 40875 3968 40917 3977
rect 40875 3928 40876 3968
rect 40916 3928 40917 3968
rect 40875 3919 40917 3928
rect 40876 3464 40916 3919
rect 40972 3557 41012 7288
rect 43036 7220 43076 7421
rect 46876 7220 46916 7421
rect 47068 7220 47108 7421
rect 47260 7220 47300 7421
rect 47417 7220 47457 7434
rect 47609 7220 47649 7434
rect 43036 7180 43124 7220
rect 46876 7180 46964 7220
rect 47068 7180 47156 7220
rect 47260 7180 47348 7220
rect 41067 6320 41109 6329
rect 41067 6280 41068 6320
rect 41108 6280 41109 6320
rect 41067 6271 41109 6280
rect 41068 4976 41108 6271
rect 41068 4927 41108 4936
rect 41164 4976 41204 4985
rect 41164 4145 41204 4936
rect 42891 4976 42933 4985
rect 42891 4936 42892 4976
rect 42932 4936 42933 4976
rect 42891 4927 42933 4936
rect 42412 4892 42452 4901
rect 41931 4724 41973 4733
rect 41931 4684 41932 4724
rect 41972 4684 41973 4724
rect 41931 4675 41973 4684
rect 42219 4724 42261 4733
rect 42219 4684 42220 4724
rect 42260 4684 42261 4724
rect 42219 4675 42261 4684
rect 41163 4136 41205 4145
rect 41163 4096 41164 4136
rect 41204 4096 41205 4136
rect 41163 4087 41205 4096
rect 41739 4136 41781 4145
rect 41739 4096 41740 4136
rect 41780 4096 41781 4136
rect 41739 4087 41781 4096
rect 41932 4136 41972 4675
rect 42220 4590 42260 4675
rect 42412 4481 42452 4852
rect 42892 4842 42932 4927
rect 42411 4472 42453 4481
rect 42411 4432 42412 4472
rect 42452 4432 42453 4472
rect 42411 4423 42453 4432
rect 42604 4304 42644 4313
rect 42644 4264 42836 4304
rect 42604 4255 42644 4264
rect 42315 4220 42357 4229
rect 42315 4180 42316 4220
rect 42356 4180 42357 4220
rect 42315 4171 42357 4180
rect 41932 4087 41972 4096
rect 42220 4136 42260 4147
rect 40971 3548 41013 3557
rect 40971 3508 40972 3548
rect 41012 3508 41013 3548
rect 40971 3499 41013 3508
rect 41740 3464 41780 4087
rect 42220 4061 42260 4096
rect 42316 4136 42356 4171
rect 42316 4085 42356 4096
rect 42796 4136 42836 4264
rect 42796 4087 42836 4096
rect 42219 4052 42261 4061
rect 42219 4012 42220 4052
rect 42260 4012 42261 4052
rect 42219 4003 42261 4012
rect 42891 4052 42933 4061
rect 42891 4012 42892 4052
rect 42932 4012 42933 4052
rect 42891 4003 42933 4012
rect 42892 3632 42932 4003
rect 42892 3583 42932 3592
rect 43084 3473 43124 7180
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44524 5144 44564 6439
rect 44524 5095 44564 5104
rect 46347 5060 46389 5069
rect 46347 5020 46348 5060
rect 46388 5020 46389 5060
rect 46347 5011 46389 5020
rect 43851 4976 43893 4985
rect 43851 4936 43852 4976
rect 43892 4936 43893 4976
rect 43851 4927 43893 4936
rect 43852 4733 43892 4927
rect 46348 4926 46388 5011
rect 46444 4976 46484 4985
rect 45195 4892 45237 4901
rect 45195 4852 45196 4892
rect 45236 4852 45237 4892
rect 45195 4843 45237 4852
rect 45196 4758 45236 4843
rect 43851 4724 43893 4733
rect 43851 4684 43852 4724
rect 43892 4684 43893 4724
rect 43851 4675 43893 4684
rect 45388 4724 45428 4733
rect 43180 4136 43220 4145
rect 43180 3977 43220 4096
rect 43179 3968 43221 3977
rect 43179 3928 43180 3968
rect 43220 3928 43221 3968
rect 43179 3919 43221 3928
rect 40876 3415 40916 3424
rect 41452 3424 41740 3464
rect 41355 2624 41397 2633
rect 41355 2584 41356 2624
rect 41396 2584 41397 2624
rect 41355 2575 41397 2584
rect 40971 2540 41013 2549
rect 40971 2500 40972 2540
rect 41012 2500 41013 2540
rect 40971 2491 41013 2500
rect 40972 1952 41012 2491
rect 41356 2129 41396 2575
rect 41355 2120 41397 2129
rect 41355 2080 41356 2120
rect 41396 2080 41397 2120
rect 41355 2071 41397 2080
rect 41356 2036 41396 2071
rect 41356 1986 41396 1996
rect 40972 1903 41012 1912
rect 41259 1952 41301 1961
rect 41259 1912 41260 1952
rect 41300 1912 41301 1952
rect 41259 1903 41301 1912
rect 41260 1818 41300 1903
rect 40683 1196 40725 1205
rect 40683 1156 40684 1196
rect 40724 1156 40725 1196
rect 40683 1147 40725 1156
rect 38572 1063 38612 1072
rect 40203 1112 40245 1121
rect 40203 1072 40204 1112
rect 40244 1072 40245 1112
rect 40203 1063 40245 1072
rect 40491 1112 40533 1121
rect 40491 1072 40492 1112
rect 40532 1072 40533 1112
rect 40491 1063 40533 1072
rect 41356 1112 41396 1121
rect 41452 1112 41492 3424
rect 41740 3415 41780 3424
rect 43083 3464 43125 3473
rect 43852 3464 43892 4675
rect 45388 4229 45428 4684
rect 46060 4724 46100 4733
rect 44139 4220 44181 4229
rect 44139 4180 44140 4220
rect 44180 4180 44181 4220
rect 44139 4171 44181 4180
rect 45195 4220 45237 4229
rect 45195 4180 45196 4220
rect 45236 4180 45237 4220
rect 45195 4171 45237 4180
rect 45387 4220 45429 4229
rect 45387 4180 45388 4220
rect 45428 4180 45429 4220
rect 45387 4171 45429 4180
rect 44043 4136 44085 4145
rect 44043 4096 44044 4136
rect 44084 4096 44085 4136
rect 44043 4087 44085 4096
rect 44044 4002 44084 4087
rect 44140 3464 44180 4171
rect 45196 4086 45236 4171
rect 45964 4136 46004 4145
rect 46060 4136 46100 4684
rect 46347 4220 46389 4229
rect 46347 4180 46348 4220
rect 46388 4180 46389 4220
rect 46347 4171 46389 4180
rect 46004 4096 46100 4136
rect 46348 4136 46388 4171
rect 45964 4087 46004 4096
rect 46348 4085 46388 4096
rect 44716 3632 44756 3643
rect 44716 3557 44756 3592
rect 44235 3548 44277 3557
rect 44235 3508 44236 3548
rect 44276 3508 44277 3548
rect 44235 3499 44277 3508
rect 44715 3548 44757 3557
rect 44715 3508 44716 3548
rect 44756 3508 44757 3548
rect 44715 3499 44757 3508
rect 43083 3424 43084 3464
rect 43124 3424 43125 3464
rect 43083 3415 43125 3424
rect 43564 3424 43852 3464
rect 43892 3424 44084 3464
rect 43564 2624 43604 3424
rect 43852 3415 43892 3424
rect 44044 3128 44084 3424
rect 44140 3415 44180 3424
rect 44236 3414 44276 3499
rect 44523 3464 44565 3473
rect 44523 3424 44524 3464
rect 44564 3424 44565 3464
rect 44523 3415 44565 3424
rect 45868 3464 45908 3473
rect 44524 3296 44564 3415
rect 44524 3247 44564 3256
rect 44044 3088 44564 3128
rect 44236 2792 44276 2801
rect 44276 2752 44372 2792
rect 44236 2743 44276 2752
rect 43851 2708 43893 2717
rect 43851 2668 43852 2708
rect 43892 2668 43893 2708
rect 43851 2659 43893 2668
rect 43564 2575 43604 2584
rect 43852 2624 43892 2659
rect 43852 2573 43892 2584
rect 43948 2540 43988 2549
rect 43948 2045 43988 2500
rect 44235 2120 44277 2129
rect 44235 2080 44236 2120
rect 44276 2080 44277 2120
rect 44235 2071 44277 2080
rect 43947 2036 43989 2045
rect 43947 1996 43948 2036
rect 43988 1996 43989 2036
rect 43947 1987 43989 1996
rect 44139 2036 44181 2045
rect 44139 1996 44140 2036
rect 44180 1996 44181 2036
rect 44139 1987 44181 1996
rect 41836 1952 41876 1961
rect 41644 1784 41684 1793
rect 41836 1784 41876 1912
rect 42220 1952 42260 1963
rect 42220 1877 42260 1912
rect 43083 1952 43125 1961
rect 43083 1912 43084 1952
rect 43124 1912 43125 1952
rect 43083 1903 43125 1912
rect 42219 1868 42261 1877
rect 42219 1828 42220 1868
rect 42260 1828 42261 1868
rect 42219 1819 42261 1828
rect 41684 1744 41876 1784
rect 41644 1735 41684 1744
rect 41396 1072 41492 1112
rect 42220 1112 42260 1819
rect 43084 1818 43124 1903
rect 44140 1364 44180 1987
rect 44236 1986 44276 2071
rect 44140 1315 44180 1324
rect 44332 1121 44372 2752
rect 44524 2624 44564 3088
rect 45196 2792 45236 2801
rect 44908 2717 44948 2761
rect 44907 2708 44949 2717
rect 44907 2668 44908 2708
rect 44948 2668 44949 2708
rect 44907 2666 44949 2668
rect 44907 2659 44908 2666
rect 44524 2575 44564 2584
rect 44812 2624 44852 2633
rect 44948 2659 44949 2666
rect 45099 2708 45141 2717
rect 45099 2668 45100 2708
rect 45140 2668 45141 2708
rect 45099 2659 45141 2668
rect 44908 2617 44948 2626
rect 44812 1457 44852 2584
rect 45100 2120 45140 2659
rect 45100 2071 45140 2080
rect 45196 2045 45236 2752
rect 45195 2036 45237 2045
rect 45195 1996 45196 2036
rect 45236 1996 45237 2036
rect 45195 1987 45237 1996
rect 45868 1961 45908 3424
rect 46444 3053 46484 4936
rect 46731 4976 46773 4985
rect 46731 4936 46732 4976
rect 46772 4936 46773 4976
rect 46731 4927 46773 4936
rect 46732 4842 46772 4927
rect 46827 4472 46869 4481
rect 46827 4432 46828 4472
rect 46868 4432 46869 4472
rect 46827 4423 46869 4432
rect 46731 4220 46773 4229
rect 46731 4180 46732 4220
rect 46772 4180 46773 4220
rect 46731 4171 46773 4180
rect 46732 4061 46772 4171
rect 46731 4052 46773 4061
rect 46731 4012 46732 4052
rect 46772 4012 46773 4052
rect 46731 4003 46773 4012
rect 46732 3464 46772 4003
rect 46443 3044 46485 3053
rect 46443 3004 46444 3044
rect 46484 3004 46485 3044
rect 46443 2995 46485 3004
rect 46732 2969 46772 3424
rect 46155 2960 46197 2969
rect 46155 2920 46156 2960
rect 46196 2920 46197 2960
rect 46155 2911 46197 2920
rect 46731 2960 46773 2969
rect 46731 2920 46732 2960
rect 46772 2920 46773 2960
rect 46731 2911 46773 2920
rect 45291 1952 45333 1961
rect 45291 1912 45292 1952
rect 45332 1912 45333 1952
rect 45291 1903 45333 1912
rect 45867 1952 45909 1961
rect 45867 1912 45868 1952
rect 45908 1912 45909 1952
rect 45867 1903 45909 1912
rect 44811 1448 44853 1457
rect 44811 1408 44812 1448
rect 44852 1408 44853 1448
rect 44811 1399 44853 1408
rect 41356 1063 41396 1072
rect 42220 1063 42260 1072
rect 42603 1112 42645 1121
rect 42603 1072 42604 1112
rect 42644 1072 42645 1112
rect 42603 1063 42645 1072
rect 44331 1112 44373 1121
rect 44331 1072 44332 1112
rect 44372 1072 44373 1112
rect 44331 1063 44373 1072
rect 45292 1112 45332 1903
rect 45292 1063 45332 1072
rect 46156 1112 46196 2911
rect 46251 2204 46293 2213
rect 46251 2164 46252 2204
rect 46292 2164 46293 2204
rect 46251 2155 46293 2164
rect 46252 1961 46292 2155
rect 46251 1952 46293 1961
rect 46251 1912 46252 1952
rect 46292 1912 46293 1952
rect 46251 1903 46293 1912
rect 46252 1818 46292 1903
rect 46156 1063 46196 1072
rect 46539 1112 46581 1121
rect 46539 1072 46540 1112
rect 46580 1072 46581 1112
rect 46828 1112 46868 4423
rect 46924 3725 46964 7180
rect 47116 4397 47156 7180
rect 47115 4388 47157 4397
rect 47115 4348 47116 4388
rect 47156 4348 47157 4388
rect 47115 4339 47157 4348
rect 47212 4136 47252 4145
rect 46923 3716 46965 3725
rect 46923 3676 46924 3716
rect 46964 3676 46965 3716
rect 46923 3667 46965 3676
rect 47115 3464 47157 3473
rect 47115 3424 47116 3464
rect 47156 3424 47157 3464
rect 47115 3415 47157 3424
rect 47116 3330 47156 3415
rect 47115 2960 47157 2969
rect 47115 2920 47116 2960
rect 47156 2920 47157 2960
rect 47115 2911 47157 2920
rect 47116 1952 47156 2911
rect 47212 2213 47252 4096
rect 47308 3557 47348 7180
rect 47404 7180 47457 7220
rect 47596 7180 47649 7220
rect 47307 3548 47349 3557
rect 47307 3508 47308 3548
rect 47348 3508 47349 3548
rect 47307 3499 47349 3508
rect 47404 2633 47444 7180
rect 47596 5069 47636 7180
rect 71404 7169 71444 36007
rect 79179 35720 79221 35729
rect 79179 35680 79180 35720
rect 79220 35680 79221 35720
rect 79179 35671 79221 35680
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 74187 33872 74229 33881
rect 74187 33832 74188 33872
rect 74228 33832 74229 33872
rect 74187 33823 74229 33832
rect 72651 32612 72693 32621
rect 72651 32572 72652 32612
rect 72692 32572 72693 32612
rect 72651 32563 72693 32572
rect 71403 7160 71445 7169
rect 71403 7120 71404 7160
rect 71444 7120 71445 7160
rect 71403 7111 71445 7120
rect 49035 6740 49077 6749
rect 49035 6700 49036 6740
rect 49076 6700 49077 6740
rect 49035 6691 49077 6700
rect 47595 5060 47637 5069
rect 47595 5020 47596 5060
rect 47636 5020 47637 5060
rect 47595 5011 47637 5020
rect 48363 5060 48405 5069
rect 48363 5020 48364 5060
rect 48404 5020 48405 5060
rect 48363 5011 48405 5020
rect 47979 4976 48021 4985
rect 47979 4936 47980 4976
rect 48020 4936 48021 4976
rect 47979 4927 48021 4936
rect 47980 3548 48020 4927
rect 48075 4892 48117 4901
rect 48075 4852 48076 4892
rect 48116 4852 48117 4892
rect 48075 4843 48117 4852
rect 48076 4397 48116 4843
rect 48075 4388 48117 4397
rect 48075 4348 48076 4388
rect 48116 4348 48117 4388
rect 48075 4339 48117 4348
rect 47788 3508 48020 3548
rect 47788 3389 47828 3508
rect 47980 3464 48020 3508
rect 47980 3415 48020 3424
rect 47787 3380 47829 3389
rect 47787 3340 47788 3380
rect 47828 3340 47829 3380
rect 47787 3331 47829 3340
rect 47403 2624 47445 2633
rect 47308 2584 47404 2624
rect 47444 2584 47445 2624
rect 47211 2204 47253 2213
rect 47211 2164 47212 2204
rect 47252 2164 47253 2204
rect 47211 2155 47253 2164
rect 47308 2036 47348 2584
rect 47403 2575 47445 2584
rect 47788 2624 47828 3331
rect 47788 2575 47828 2584
rect 48076 2624 48116 4339
rect 48364 4304 48404 5011
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 48268 4264 48364 4304
rect 48268 3464 48308 4264
rect 48364 4255 48404 4264
rect 48940 4136 48980 4147
rect 48940 4061 48980 4096
rect 48556 4052 48596 4061
rect 48939 4052 48981 4061
rect 48596 4012 48692 4052
rect 48556 4003 48596 4012
rect 48268 3415 48308 3424
rect 48363 3464 48405 3473
rect 48363 3424 48364 3464
rect 48404 3424 48405 3464
rect 48363 3415 48405 3424
rect 48364 3330 48404 3415
rect 48652 3296 48692 4012
rect 48939 4012 48940 4052
rect 48980 4012 48981 4052
rect 48939 4003 48981 4012
rect 49036 3632 49076 6691
rect 49611 6236 49653 6245
rect 49611 6196 49612 6236
rect 49652 6196 49653 6236
rect 49611 6187 49653 6196
rect 49419 5396 49461 5405
rect 49419 5356 49420 5396
rect 49460 5356 49461 5396
rect 49419 5347 49461 5356
rect 49420 5060 49460 5347
rect 49420 5011 49460 5020
rect 49324 4976 49364 4985
rect 49228 4936 49324 4976
rect 49228 4313 49268 4936
rect 49324 4927 49364 4936
rect 49515 4976 49557 4985
rect 49515 4936 49516 4976
rect 49556 4936 49557 4976
rect 49515 4927 49557 4936
rect 49516 4842 49556 4927
rect 49612 4724 49652 6187
rect 72652 5489 72692 32563
rect 74188 28328 74228 33823
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 78507 32696 78549 32705
rect 78507 32656 78508 32696
rect 78548 32656 78549 32696
rect 78507 32647 78549 32656
rect 74188 28279 74228 28288
rect 75820 28160 75860 28169
rect 75820 18005 75860 28120
rect 75819 17996 75861 18005
rect 75819 17956 75820 17996
rect 75860 17956 75861 17996
rect 75819 17947 75861 17956
rect 78220 17072 78260 17081
rect 78124 17032 78220 17072
rect 78124 16484 78164 17032
rect 78220 17023 78260 17032
rect 78411 16820 78453 16829
rect 78411 16780 78412 16820
rect 78452 16780 78453 16820
rect 78411 16771 78453 16780
rect 78124 16435 78164 16444
rect 78412 16232 78452 16771
rect 78508 16736 78548 32647
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 79180 31697 79220 35671
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 80140 32948 80180 32957
rect 80140 32705 80180 32908
rect 80428 32780 80468 36679
rect 81483 35048 81525 35057
rect 81483 35008 81484 35048
rect 81524 35008 81525 35048
rect 81483 34999 81525 35008
rect 80907 33872 80949 33881
rect 80907 33832 80908 33872
rect 80948 33832 80949 33872
rect 80907 33823 80949 33832
rect 80812 33704 80852 33713
rect 80812 33368 80852 33664
rect 80620 33328 80852 33368
rect 80524 33116 80564 33125
rect 80620 33116 80660 33328
rect 80811 33200 80853 33209
rect 80908 33200 80948 33823
rect 81196 33704 81236 33713
rect 80811 33160 80812 33200
rect 80852 33160 80948 33200
rect 81100 33664 81196 33704
rect 80811 33151 80853 33160
rect 80564 33076 80660 33116
rect 80524 33067 80564 33076
rect 80812 32864 80852 33151
rect 80812 32815 80852 32824
rect 80908 32864 80948 32873
rect 80428 32740 80660 32780
rect 80139 32696 80181 32705
rect 80139 32656 80140 32696
rect 80180 32656 80181 32696
rect 80139 32647 80181 32656
rect 80332 32696 80372 32705
rect 80372 32656 80468 32696
rect 80332 32647 80372 32656
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 79179 31688 79221 31697
rect 79179 31648 79180 31688
rect 79220 31648 79221 31688
rect 79179 31639 79221 31648
rect 79180 30605 79220 31639
rect 80331 31436 80373 31445
rect 80428 31436 80468 32656
rect 80331 31396 80332 31436
rect 80372 31396 80468 31436
rect 80331 31387 80373 31396
rect 80332 31302 80372 31387
rect 80140 31184 80180 31193
rect 79660 31144 80140 31184
rect 79660 30680 79700 31144
rect 79660 30631 79700 30640
rect 78603 30596 78645 30605
rect 78603 30556 78604 30596
rect 78644 30556 78645 30596
rect 78603 30547 78645 30556
rect 79179 30596 79221 30605
rect 79179 30556 79180 30596
rect 79220 30556 79221 30596
rect 79179 30547 79221 30556
rect 78604 17072 78644 30547
rect 79180 30462 79220 30547
rect 79372 30428 79412 30437
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 79180 29840 79220 29849
rect 79372 29840 79412 30388
rect 79659 30176 79701 30185
rect 79659 30136 79660 30176
rect 79700 30136 79701 30176
rect 79659 30127 79701 30136
rect 79220 29800 79412 29840
rect 78796 29756 78836 29765
rect 78796 29009 78836 29716
rect 78795 29000 78837 29009
rect 78795 28960 78796 29000
rect 78836 28960 78837 29000
rect 78795 28951 78837 28960
rect 79180 28925 79220 29800
rect 79660 29252 79700 30127
rect 79660 29203 79700 29212
rect 79756 29168 79796 29177
rect 79852 29168 79892 31144
rect 80140 31135 80180 31144
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 80043 30848 80085 30857
rect 80043 30808 80044 30848
rect 80084 30808 80085 30848
rect 80043 30799 80085 30808
rect 80044 30764 80084 30799
rect 80044 30713 80084 30724
rect 79948 30680 79988 30689
rect 79948 30185 79988 30640
rect 80524 30680 80564 30689
rect 80332 30512 80372 30521
rect 80524 30512 80564 30640
rect 80372 30472 80564 30512
rect 80332 30463 80372 30472
rect 80043 30260 80085 30269
rect 80043 30220 80044 30260
rect 80084 30220 80085 30260
rect 80043 30211 80085 30220
rect 79947 30176 79989 30185
rect 79947 30136 79948 30176
rect 79988 30136 79989 30176
rect 79947 30127 79989 30136
rect 80044 29840 80084 30211
rect 80620 30185 80660 32740
rect 80812 32192 80852 32201
rect 80716 32152 80812 32192
rect 80716 31604 80756 32152
rect 80812 32143 80852 32152
rect 80716 31555 80756 31564
rect 80908 31268 80948 32824
rect 81100 32696 81140 33664
rect 81196 33655 81236 33664
rect 81196 32864 81236 32873
rect 81236 32824 81332 32864
rect 81196 32815 81236 32824
rect 81195 32696 81237 32705
rect 81100 32656 81196 32696
rect 81236 32656 81237 32696
rect 81195 32647 81237 32656
rect 81196 32192 81236 32647
rect 81099 31352 81141 31361
rect 81099 31312 81100 31352
rect 81140 31312 81141 31352
rect 81099 31303 81141 31312
rect 81004 31268 81044 31277
rect 80908 31228 81004 31268
rect 81004 31109 81044 31228
rect 81100 31218 81140 31303
rect 81003 31100 81045 31109
rect 81003 31060 81004 31100
rect 81044 31060 81045 31100
rect 81003 31051 81045 31060
rect 80715 30848 80757 30857
rect 80715 30808 80716 30848
rect 80756 30808 80757 30848
rect 80715 30799 80757 30808
rect 80619 30176 80661 30185
rect 80619 30136 80620 30176
rect 80660 30136 80661 30176
rect 80619 30127 80661 30136
rect 80044 29791 80084 29800
rect 80620 29681 80660 30127
rect 80619 29672 80661 29681
rect 80619 29632 80620 29672
rect 80660 29632 80661 29672
rect 80619 29623 80661 29632
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 80044 29168 80084 29177
rect 79852 29128 80044 29168
rect 79371 29000 79413 29009
rect 79371 28960 79372 29000
rect 79412 28960 79413 29000
rect 79371 28951 79413 28960
rect 79179 28916 79221 28925
rect 79179 28876 79180 28916
rect 79220 28876 79221 28916
rect 79179 28867 79221 28876
rect 79372 28866 79412 28951
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 79756 27749 79796 29128
rect 79948 28328 79988 29128
rect 80044 29119 80084 29128
rect 80331 28748 80373 28757
rect 80331 28708 80332 28748
rect 80372 28708 80373 28748
rect 80331 28699 80373 28708
rect 79852 28288 79948 28328
rect 79755 27740 79797 27749
rect 79755 27700 79756 27740
rect 79796 27700 79797 27740
rect 79755 27691 79797 27700
rect 79852 27656 79892 28288
rect 79948 28279 79988 28288
rect 80235 28328 80277 28337
rect 80235 28288 80236 28328
rect 80276 28288 80277 28328
rect 80235 28279 80277 28288
rect 80332 28328 80372 28699
rect 80716 28580 80756 30799
rect 80908 30680 80948 30689
rect 81196 30680 81236 32152
rect 81292 31436 81332 32824
rect 81388 31445 81428 31476
rect 81387 31436 81429 31445
rect 81292 31396 81388 31436
rect 81428 31396 81429 31436
rect 81387 31387 81429 31396
rect 80948 30640 81236 30680
rect 81388 31352 81428 31387
rect 80811 29252 80853 29261
rect 80811 29212 80812 29252
rect 80852 29212 80853 29252
rect 80811 29203 80853 29212
rect 80812 29118 80852 29203
rect 80908 29168 80948 30640
rect 81388 30521 81428 31312
rect 81387 30512 81429 30521
rect 81387 30472 81388 30512
rect 81428 30472 81429 30512
rect 81387 30463 81429 30472
rect 81388 30008 81428 30017
rect 81195 29672 81237 29681
rect 81195 29632 81196 29672
rect 81236 29632 81237 29672
rect 81195 29623 81237 29632
rect 81196 29538 81236 29623
rect 81388 29261 81428 29968
rect 81387 29252 81429 29261
rect 81387 29212 81388 29252
rect 81428 29212 81429 29252
rect 81387 29203 81429 29212
rect 81196 29168 81236 29177
rect 80908 29128 81196 29168
rect 81196 29119 81236 29128
rect 81195 28916 81237 28925
rect 81195 28876 81196 28916
rect 81236 28876 81237 28916
rect 81195 28867 81237 28876
rect 80716 28540 80948 28580
rect 80620 28496 80660 28505
rect 80660 28456 80852 28496
rect 80620 28447 80660 28456
rect 80812 28328 80852 28456
rect 80372 28288 80468 28328
rect 80332 28279 80372 28288
rect 80236 28194 80276 28279
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 80428 27824 80468 28288
rect 80812 28279 80852 28288
rect 80908 28232 80948 28540
rect 80236 27784 80468 27824
rect 80716 28192 80948 28232
rect 81196 28328 81236 28867
rect 80140 27656 80180 27665
rect 79852 27616 80140 27656
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 79852 26984 79892 26993
rect 79852 26312 79892 26944
rect 80140 26909 80180 27616
rect 80139 26900 80181 26909
rect 80139 26860 80140 26900
rect 80180 26860 80181 26900
rect 80139 26851 80181 26860
rect 80236 26816 80276 27784
rect 80523 27740 80565 27749
rect 80523 27700 80524 27740
rect 80564 27700 80565 27740
rect 80523 27691 80565 27700
rect 80236 26767 80276 26776
rect 80428 27656 80468 27665
rect 80428 26741 80468 27616
rect 80524 27606 80564 27691
rect 80524 26909 80564 26940
rect 80523 26900 80565 26909
rect 80523 26860 80524 26900
rect 80564 26860 80565 26900
rect 80523 26851 80565 26860
rect 80524 26816 80564 26851
rect 80139 26732 80181 26741
rect 80139 26692 80140 26732
rect 80180 26692 80181 26732
rect 80139 26683 80181 26692
rect 80427 26732 80469 26741
rect 80427 26692 80428 26732
rect 80468 26692 80469 26732
rect 80427 26683 80469 26692
rect 80140 26598 80180 26683
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 79852 26272 80276 26312
rect 80236 26228 80276 26272
rect 80236 26179 80276 26188
rect 80524 25976 80564 26776
rect 80620 26153 80660 26238
rect 80619 26144 80661 26153
rect 80619 26104 80620 26144
rect 80660 26104 80661 26144
rect 80619 26095 80661 26104
rect 80524 25936 80660 25976
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 80620 25481 80660 25936
rect 80236 25472 80276 25481
rect 80619 25472 80661 25481
rect 80276 25432 80468 25472
rect 80236 25423 80276 25432
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 80236 24716 80276 24725
rect 80428 24716 80468 25432
rect 80619 25432 80620 25472
rect 80660 25432 80661 25472
rect 80619 25423 80661 25432
rect 80620 25304 80660 25313
rect 80716 25304 80756 28192
rect 80812 27404 80852 27413
rect 80812 26816 80852 27364
rect 80812 26767 80852 26776
rect 81196 26816 81236 28288
rect 81196 26153 81236 26776
rect 81195 26144 81237 26153
rect 81484 26144 81524 34999
rect 81580 28337 81620 36763
rect 83307 36644 83349 36653
rect 83307 36604 83308 36644
rect 83348 36604 83349 36644
rect 83307 36595 83349 36604
rect 82059 34292 82101 34301
rect 82059 34252 82060 34292
rect 82100 34252 82101 34292
rect 82059 34243 82101 34252
rect 82060 33704 82100 34243
rect 82251 34124 82293 34133
rect 82251 34084 82252 34124
rect 82292 34084 82293 34124
rect 82251 34075 82293 34084
rect 82100 33664 82196 33704
rect 82060 33655 82100 33664
rect 82060 32948 82100 32957
rect 81964 32908 82060 32948
rect 81867 32696 81909 32705
rect 81867 32656 81868 32696
rect 81908 32656 81909 32696
rect 81867 32647 81909 32656
rect 81868 32562 81908 32647
rect 81964 31697 82004 32908
rect 82060 32899 82100 32908
rect 82060 32192 82100 32201
rect 82156 32192 82196 33664
rect 82100 32152 82196 32192
rect 81963 31688 82005 31697
rect 81963 31648 81964 31688
rect 82004 31648 82005 31688
rect 81963 31639 82005 31648
rect 81675 31352 81717 31361
rect 81675 31312 81676 31352
rect 81716 31312 81717 31352
rect 81675 31303 81717 31312
rect 81676 29849 81716 31303
rect 81772 30680 81812 30689
rect 82060 30680 82100 32152
rect 81812 30640 82196 30680
rect 81772 30269 81812 30640
rect 82059 30512 82101 30521
rect 82059 30472 82060 30512
rect 82100 30472 82101 30512
rect 82059 30463 82101 30472
rect 81771 30260 81813 30269
rect 81771 30220 81772 30260
rect 81812 30220 81813 30260
rect 81771 30211 81813 30220
rect 81675 29840 81717 29849
rect 81675 29800 81676 29840
rect 81716 29800 81717 29840
rect 81675 29791 81717 29800
rect 81772 29840 81812 29849
rect 81676 29706 81716 29791
rect 81579 28328 81621 28337
rect 81579 28288 81580 28328
rect 81620 28288 81621 28328
rect 81579 28279 81621 28288
rect 81580 27380 81620 28279
rect 81580 27340 81716 27380
rect 81195 26104 81196 26144
rect 81236 26104 81237 26144
rect 81195 26095 81237 26104
rect 81388 26104 81484 26144
rect 81291 25640 81333 25649
rect 81291 25600 81292 25640
rect 81332 25600 81333 25640
rect 81291 25591 81333 25600
rect 81196 25472 81236 25481
rect 80660 25264 80756 25304
rect 80812 25432 81196 25472
rect 80620 25255 80660 25264
rect 80523 25220 80565 25229
rect 80523 25180 80524 25220
rect 80564 25180 80565 25220
rect 80523 25171 80565 25180
rect 80524 25086 80564 25171
rect 80619 25136 80661 25145
rect 80619 25096 80620 25136
rect 80660 25096 80661 25136
rect 80619 25087 80661 25096
rect 80276 24676 80468 24716
rect 80236 24667 80276 24676
rect 80620 24632 80660 25087
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 80620 23717 80660 24592
rect 80812 23792 80852 25432
rect 81196 25423 81236 25432
rect 80907 25304 80949 25313
rect 80907 25264 80908 25304
rect 80948 25264 80949 25304
rect 80907 25255 80949 25264
rect 80812 23743 80852 23752
rect 80619 23708 80661 23717
rect 80619 23668 80620 23708
rect 80660 23668 80661 23708
rect 80619 23659 80661 23668
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 79467 20768 79509 20777
rect 79467 20728 79468 20768
rect 79508 20728 79509 20768
rect 80908 20768 80948 25255
rect 81196 23792 81236 23803
rect 81196 23717 81236 23752
rect 81195 23708 81237 23717
rect 81195 23668 81196 23708
rect 81236 23668 81237 23708
rect 81195 23659 81237 23668
rect 81292 22868 81332 25591
rect 81388 24632 81428 26104
rect 81484 26095 81524 26104
rect 81676 25649 81716 27340
rect 81675 25640 81717 25649
rect 81675 25600 81676 25640
rect 81716 25600 81717 25640
rect 81675 25591 81717 25600
rect 81772 25472 81812 29800
rect 82060 29840 82100 30463
rect 82060 29791 82100 29800
rect 82060 29168 82100 29177
rect 82156 29168 82196 30640
rect 82100 29128 82196 29168
rect 82060 29119 82100 29128
rect 82060 28328 82100 28337
rect 82252 28328 82292 34075
rect 83212 33452 83252 33461
rect 83116 33412 83212 33452
rect 83116 33209 83156 33412
rect 83212 33403 83252 33412
rect 83115 33200 83157 33209
rect 83115 33160 83116 33200
rect 83156 33160 83157 33200
rect 83115 33151 83157 33160
rect 83116 30941 83156 33151
rect 83212 31940 83252 31949
rect 83212 31109 83252 31900
rect 83211 31100 83253 31109
rect 83211 31060 83212 31100
rect 83252 31060 83253 31100
rect 83211 31051 83253 31060
rect 83115 30932 83157 30941
rect 83115 30892 83116 30932
rect 83156 30892 83157 30932
rect 83115 30883 83157 30892
rect 82923 30848 82965 30857
rect 82923 30808 82924 30848
rect 82964 30808 82965 30848
rect 82923 30799 82965 30808
rect 82924 30714 82964 30799
rect 83308 29849 83348 36595
rect 91025 36540 91065 36763
rect 92176 36728 92218 36737
rect 92176 36688 92177 36728
rect 92217 36688 92218 36728
rect 92176 36679 92218 36688
rect 92177 36540 92217 36679
rect 92428 36560 92468 36931
rect 92752 36896 92794 36905
rect 92752 36856 92753 36896
rect 92793 36856 92794 36896
rect 92752 36847 92794 36856
rect 92753 36540 92793 36847
rect 83307 29840 83349 29849
rect 83307 29800 83308 29840
rect 83348 29800 83349 29840
rect 83307 29791 83349 29800
rect 83212 29336 83252 29345
rect 83308 29336 83348 29791
rect 83252 29296 83348 29336
rect 83212 29287 83252 29296
rect 83211 28748 83253 28757
rect 83211 28708 83212 28748
rect 83252 28708 83253 28748
rect 83211 28699 83253 28708
rect 83212 28580 83252 28699
rect 83212 28531 83252 28540
rect 82100 28288 82292 28328
rect 82060 26816 82100 28288
rect 83307 28244 83349 28253
rect 83307 28204 83308 28244
rect 83348 28204 83349 28244
rect 83307 28195 83349 28204
rect 83308 27749 83348 28195
rect 83307 27740 83349 27749
rect 83307 27700 83308 27740
rect 83348 27700 83349 27740
rect 83307 27691 83349 27700
rect 83212 27068 83252 27077
rect 83308 27068 83348 27691
rect 83252 27028 83348 27068
rect 83212 27019 83252 27028
rect 82060 26767 82100 26776
rect 82635 26732 82677 26741
rect 82635 26692 82636 26732
rect 82676 26692 82677 26732
rect 82635 26683 82677 26692
rect 82636 25976 82676 26683
rect 82676 25936 82772 25976
rect 82636 25927 82676 25936
rect 81484 25432 81812 25472
rect 81484 25304 81524 25432
rect 81484 25255 81524 25264
rect 81580 25304 81620 25313
rect 81580 25229 81620 25264
rect 81579 25220 81621 25229
rect 81579 25180 81580 25220
rect 81620 25180 81621 25220
rect 81579 25171 81621 25180
rect 81484 24632 81524 24641
rect 81388 24592 81484 24632
rect 81484 23801 81524 24592
rect 81580 24557 81620 25171
rect 81579 24548 81621 24557
rect 81579 24508 81580 24548
rect 81620 24508 81621 24548
rect 81579 24499 81621 24508
rect 81676 24053 81716 25432
rect 81867 25304 81909 25313
rect 81867 25264 81868 25304
rect 81908 25264 81909 25304
rect 81867 25255 81909 25264
rect 81868 25170 81908 25255
rect 82636 24548 82676 24559
rect 82636 24473 82676 24508
rect 82635 24464 82677 24473
rect 82635 24424 82636 24464
rect 82676 24424 82677 24464
rect 82635 24415 82677 24424
rect 82732 24389 82772 25936
rect 85420 24634 85861 24674
rect 82731 24380 82773 24389
rect 82731 24340 82732 24380
rect 82772 24340 82773 24380
rect 82731 24331 82773 24340
rect 81675 24044 81717 24053
rect 81675 24004 81676 24044
rect 81716 24004 81717 24044
rect 81675 23995 81717 24004
rect 83211 24044 83253 24053
rect 83211 24004 83212 24044
rect 83252 24004 83253 24044
rect 83211 23995 83253 24004
rect 83212 23910 83252 23995
rect 81483 23792 81525 23801
rect 81483 23752 81484 23792
rect 81524 23752 81525 23792
rect 81483 23743 81525 23752
rect 82059 23792 82101 23801
rect 82059 23752 82060 23792
rect 82100 23752 82101 23792
rect 82059 23743 82101 23752
rect 81292 22828 81524 22868
rect 81484 21029 81524 22828
rect 81483 21020 81525 21029
rect 81483 20980 81484 21020
rect 81524 20980 81525 21020
rect 81483 20971 81525 20980
rect 81100 20768 81140 20777
rect 80908 20728 81100 20768
rect 79467 20719 79509 20728
rect 81100 20719 81140 20728
rect 81388 20768 81428 20777
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 78604 17023 78644 17032
rect 79468 17072 79508 20719
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 78508 16696 78644 16736
rect 78412 16183 78452 16192
rect 78507 16232 78549 16241
rect 78507 16192 78508 16232
rect 78548 16192 78549 16232
rect 78604 16232 78644 16696
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 78796 16232 78836 16241
rect 78604 16192 78796 16232
rect 78507 16183 78549 16192
rect 78796 16183 78836 16192
rect 78508 16098 78548 16183
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 78507 6488 78549 6497
rect 78507 6448 78508 6488
rect 78548 6448 78549 6488
rect 78507 6439 78549 6448
rect 78508 6354 78548 6439
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 72651 5480 72693 5489
rect 72651 5440 72652 5480
rect 72692 5440 72693 5480
rect 72651 5431 72693 5440
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 52203 5228 52245 5237
rect 52203 5188 52204 5228
rect 52244 5188 52245 5228
rect 52203 5179 52245 5188
rect 49995 5144 50037 5153
rect 49995 5104 49996 5144
rect 50036 5104 50037 5144
rect 49995 5095 50037 5104
rect 49996 5010 50036 5095
rect 49900 4976 49940 4985
rect 49516 4684 49652 4724
rect 49707 4724 49749 4733
rect 49707 4684 49708 4724
rect 49748 4684 49749 4724
rect 49227 4304 49269 4313
rect 49227 4264 49228 4304
rect 49268 4264 49269 4304
rect 49227 4255 49269 4264
rect 49228 3809 49268 4255
rect 49227 3800 49269 3809
rect 49227 3760 49228 3800
rect 49268 3760 49269 3800
rect 49227 3751 49269 3760
rect 49036 3583 49076 3592
rect 49228 3557 49268 3751
rect 49323 3632 49365 3641
rect 49323 3592 49324 3632
rect 49364 3592 49365 3632
rect 49323 3583 49365 3592
rect 49516 3632 49556 4684
rect 49707 4675 49749 4684
rect 49708 4590 49748 4675
rect 49900 4313 49940 4936
rect 52204 4976 52244 5179
rect 79468 5069 79508 17032
rect 81388 16829 81428 20728
rect 81484 20768 81524 20971
rect 81484 20719 81524 20728
rect 81772 20936 81812 20945
rect 81772 20684 81812 20896
rect 82060 20861 82100 23743
rect 85420 23717 85460 24634
rect 87953 24296 87993 24640
rect 90460 24389 90500 24621
rect 92572 24473 92612 24621
rect 92571 24464 92613 24473
rect 92571 24424 92572 24464
rect 92612 24424 92613 24464
rect 92571 24415 92613 24424
rect 90459 24380 90501 24389
rect 90459 24340 90460 24380
rect 90500 24340 90501 24380
rect 90459 24331 90501 24340
rect 87916 24256 87993 24296
rect 87916 24053 87956 24256
rect 87915 24044 87957 24053
rect 87915 24004 87916 24044
rect 87956 24004 87957 24044
rect 87915 23995 87957 24004
rect 82443 23708 82485 23717
rect 82443 23668 82444 23708
rect 82484 23668 82485 23708
rect 82443 23659 82485 23668
rect 85419 23708 85461 23717
rect 85419 23668 85420 23708
rect 85460 23668 85461 23708
rect 85419 23659 85461 23668
rect 82059 20852 82101 20861
rect 82059 20812 82060 20852
rect 82100 20812 82101 20852
rect 82059 20803 82101 20812
rect 82444 20768 82484 23659
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 84459 21020 84501 21029
rect 84459 20980 84460 21020
rect 84500 20980 84501 21020
rect 84459 20971 84501 20980
rect 84460 20886 84500 20971
rect 82444 20719 82484 20728
rect 83307 20768 83349 20777
rect 83307 20728 83308 20768
rect 83348 20728 83349 20768
rect 83307 20719 83349 20728
rect 82060 20684 82100 20693
rect 81772 20644 82060 20684
rect 82060 20635 82100 20644
rect 83308 20634 83348 20719
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 82731 20096 82773 20105
rect 82731 20056 82732 20096
rect 82772 20056 82773 20096
rect 82731 20047 82773 20056
rect 96747 20096 96789 20105
rect 96747 20056 96748 20096
rect 96788 20056 96789 20096
rect 96747 20047 96789 20056
rect 80619 16820 80661 16829
rect 80619 16780 80620 16820
rect 80660 16780 80661 16820
rect 80619 16771 80661 16780
rect 81387 16820 81429 16829
rect 81387 16780 81388 16820
rect 81428 16780 81429 16820
rect 81387 16771 81429 16780
rect 80620 16686 80660 16771
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 81388 9269 81428 16771
rect 81387 9260 81429 9269
rect 81387 9220 81388 9260
rect 81428 9220 81429 9260
rect 81387 9211 81429 9220
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 82732 7085 82772 20047
rect 96748 19962 96788 20047
rect 98571 19928 98613 19937
rect 98571 19888 98572 19928
rect 98612 19888 98613 19928
rect 98571 19879 98613 19888
rect 98572 19794 98612 19879
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 98859 17996 98901 18005
rect 98859 17956 98860 17996
rect 98900 17956 98901 17996
rect 98859 17947 98901 17956
rect 98860 9428 98900 17947
rect 98859 9419 98901 9428
rect 98859 9379 98860 9419
rect 98900 9379 98901 9419
rect 98859 9370 98901 9379
rect 82731 7076 82773 7085
rect 82731 7036 82732 7076
rect 82772 7036 82773 7076
rect 82731 7027 82773 7036
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 80523 6656 80565 6665
rect 80523 6616 80524 6656
rect 80564 6616 80565 6656
rect 80523 6607 80565 6616
rect 80524 6522 80564 6607
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 53931 5060 53973 5069
rect 53931 5020 53932 5060
rect 53972 5020 53973 5060
rect 53931 5011 53973 5020
rect 79467 5060 79509 5069
rect 79467 5020 79468 5060
rect 79508 5020 79509 5060
rect 79467 5011 79509 5020
rect 50379 4808 50421 4817
rect 50379 4768 50380 4808
rect 50420 4768 50421 4808
rect 50379 4759 50421 4768
rect 49899 4304 49941 4313
rect 49899 4264 49900 4304
rect 49940 4264 49941 4304
rect 49899 4255 49941 4264
rect 49611 4136 49653 4145
rect 49611 4096 49612 4136
rect 49652 4096 49653 4136
rect 49611 4087 49653 4096
rect 49803 4136 49845 4145
rect 49803 4096 49804 4136
rect 49844 4096 49845 4136
rect 49803 4087 49845 4096
rect 49516 3583 49556 3592
rect 49227 3548 49269 3557
rect 49227 3508 49228 3548
rect 49268 3508 49269 3548
rect 49227 3499 49269 3508
rect 49228 3464 49268 3499
rect 49324 3498 49364 3583
rect 49228 3414 49268 3424
rect 48652 3247 48692 3256
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 48460 2792 48500 2801
rect 48076 2575 48116 2584
rect 48171 2624 48213 2633
rect 48171 2584 48172 2624
rect 48212 2584 48213 2624
rect 48171 2575 48213 2584
rect 48363 2624 48405 2633
rect 48363 2584 48364 2624
rect 48404 2584 48405 2624
rect 48363 2575 48405 2584
rect 48172 2490 48212 2575
rect 47116 1903 47156 1912
rect 47212 1996 47348 2036
rect 47499 2036 47541 2045
rect 47499 1996 47500 2036
rect 47540 1996 47541 2036
rect 46924 1112 46964 1121
rect 46828 1072 46924 1112
rect 46539 1063 46581 1072
rect 46924 1063 46964 1072
rect 47212 1112 47252 1996
rect 47499 1987 47541 1996
rect 47500 1902 47540 1987
rect 48364 1868 48404 2575
rect 48460 2045 48500 2752
rect 48939 2204 48981 2213
rect 48939 2164 48940 2204
rect 48980 2164 48981 2204
rect 48939 2155 48981 2164
rect 48459 2036 48501 2045
rect 48459 1996 48460 2036
rect 48500 1996 48501 2036
rect 48459 1987 48501 1996
rect 48460 1868 48500 1877
rect 48364 1828 48460 1868
rect 48460 1819 48500 1828
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 47307 1448 47349 1457
rect 47307 1408 47308 1448
rect 47348 1408 47349 1448
rect 47307 1399 47349 1408
rect 47787 1448 47829 1457
rect 47787 1408 47788 1448
rect 47828 1408 47829 1448
rect 47787 1399 47829 1408
rect 47212 1063 47252 1072
rect 47308 1112 47348 1399
rect 47788 1364 47828 1399
rect 47788 1313 47828 1324
rect 47596 1280 47636 1289
rect 47596 1121 47636 1240
rect 47308 1063 47348 1072
rect 47595 1112 47637 1121
rect 47595 1072 47596 1112
rect 47636 1072 47637 1112
rect 47595 1063 47637 1072
rect 48940 1112 48980 2155
rect 49612 1952 49652 4087
rect 49804 4002 49844 4087
rect 50187 4052 50229 4061
rect 50187 4012 50188 4052
rect 50228 4012 50229 4052
rect 50187 4003 50229 4012
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 49804 3632 49844 3641
rect 49707 3548 49749 3557
rect 49707 3508 49708 3548
rect 49748 3508 49749 3548
rect 49804 3548 49844 3592
rect 49899 3548 49941 3557
rect 49804 3508 49900 3548
rect 49940 3508 49941 3548
rect 49707 3499 49749 3508
rect 49899 3499 49941 3508
rect 49708 3464 49748 3499
rect 49708 3413 49748 3424
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 50188 2120 50228 4003
rect 49612 1903 49652 1912
rect 49804 2080 50228 2120
rect 48940 1063 48980 1072
rect 49804 1112 49844 2080
rect 50380 1952 50420 4759
rect 52204 4481 52244 4936
rect 52492 4976 52532 4985
rect 52203 4472 52245 4481
rect 52203 4432 52204 4472
rect 52244 4432 52245 4472
rect 52203 4423 52245 4432
rect 51532 4136 51572 4147
rect 51532 4061 51572 4096
rect 52395 4136 52437 4145
rect 52395 4096 52396 4136
rect 52436 4096 52437 4136
rect 52395 4087 52437 4096
rect 51148 4052 51188 4061
rect 50956 3968 50996 3977
rect 50764 3928 50956 3968
rect 50476 3464 50516 3475
rect 50764 3473 50804 3928
rect 50956 3919 50996 3928
rect 50859 3716 50901 3725
rect 50859 3676 50860 3716
rect 50900 3676 50901 3716
rect 50859 3667 50901 3676
rect 50860 3548 50900 3667
rect 50860 3499 50900 3508
rect 50476 3389 50516 3424
rect 50763 3464 50805 3473
rect 50763 3424 50764 3464
rect 50804 3424 50805 3464
rect 50763 3415 50805 3424
rect 50475 3380 50517 3389
rect 50475 3340 50476 3380
rect 50516 3340 50517 3380
rect 50475 3331 50517 3340
rect 50764 3330 50804 3415
rect 51148 3296 51188 4012
rect 51531 4052 51573 4061
rect 51531 4012 51532 4052
rect 51572 4012 51573 4052
rect 51531 4003 51573 4012
rect 52396 4002 52436 4087
rect 52492 3725 52532 4936
rect 52588 4976 52628 4987
rect 52588 4901 52628 4936
rect 52587 4892 52629 4901
rect 52587 4852 52588 4892
rect 52628 4852 52629 4892
rect 52587 4843 52629 4852
rect 52876 4724 52916 4733
rect 52684 4684 52876 4724
rect 52491 3716 52533 3725
rect 52491 3676 52492 3716
rect 52532 3676 52533 3716
rect 52491 3667 52533 3676
rect 52684 3548 52724 4684
rect 52876 4675 52916 4684
rect 53067 4052 53109 4061
rect 53067 4012 53068 4052
rect 53108 4012 53109 4052
rect 53067 4003 53109 4012
rect 52684 3499 52724 3508
rect 53068 3464 53108 4003
rect 53548 3968 53588 3977
rect 53548 3725 53588 3928
rect 53547 3716 53589 3725
rect 53547 3676 53548 3716
rect 53588 3676 53589 3716
rect 53547 3667 53589 3676
rect 53068 3415 53108 3424
rect 53932 3464 53972 5011
rect 55083 4892 55125 4901
rect 55083 4852 55084 4892
rect 55124 4852 55125 4892
rect 55083 4843 55125 4852
rect 55084 3632 55124 4843
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 55084 3583 55124 3592
rect 80715 3632 80757 3641
rect 80715 3592 80716 3632
rect 80756 3592 80757 3632
rect 80715 3583 80757 3592
rect 53932 3415 53972 3424
rect 51148 3247 51188 3256
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 50859 2036 50901 2045
rect 50859 1996 50860 2036
rect 50900 1996 50901 2036
rect 50859 1987 50901 1996
rect 50476 1952 50516 1961
rect 50380 1912 50476 1952
rect 50476 1903 50516 1912
rect 50860 1902 50900 1987
rect 80716 1541 80756 3583
rect 80907 3548 80949 3557
rect 80907 3508 80908 3548
rect 80948 3508 80949 3548
rect 80907 3499 80949 3508
rect 80908 1877 80948 3499
rect 80907 1868 80949 1877
rect 80907 1828 80908 1868
rect 80948 1828 80949 1868
rect 80907 1819 80949 1828
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 80715 1532 80757 1541
rect 80715 1492 80716 1532
rect 80756 1492 80757 1532
rect 80715 1483 80757 1492
rect 90920 1479 90978 1480
rect 90536 1460 90578 1469
rect 90536 1420 90537 1460
rect 90577 1420 90578 1460
rect 90920 1439 90929 1479
rect 90969 1439 90978 1479
rect 90920 1438 90978 1439
rect 91112 1479 91170 1480
rect 91112 1439 91121 1479
rect 91161 1439 91170 1479
rect 91112 1438 91170 1439
rect 91304 1479 91362 1480
rect 91304 1439 91313 1479
rect 91353 1439 91362 1479
rect 91304 1438 91362 1439
rect 90536 1411 90578 1420
rect 90729 1205 90769 1421
rect 90728 1196 90770 1205
rect 90728 1156 90729 1196
rect 90769 1156 90770 1196
rect 90728 1147 90770 1156
rect 49804 1063 49844 1072
rect 50187 1112 50229 1121
rect 50187 1072 50188 1112
rect 50228 1072 50229 1112
rect 50187 1063 50229 1072
rect 35499 1028 35541 1037
rect 35499 988 35500 1028
rect 35540 988 35541 1028
rect 35499 979 35541 988
rect 38187 1028 38229 1037
rect 38187 988 38188 1028
rect 38228 988 38229 1028
rect 38187 979 38229 988
rect 38476 978 38516 1063
rect 42604 978 42644 1063
rect 46540 978 46580 1063
rect 50188 978 50228 1063
rect 27051 944 27093 953
rect 27051 904 27052 944
rect 27092 904 27093 944
rect 27051 895 27093 904
rect 28299 944 28341 953
rect 28299 904 28300 944
rect 28340 904 28341 944
rect 28299 895 28341 904
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 844 37948 884 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 652 37528 692 37568
rect 19756 37444 19796 37484
rect 20428 37444 20468 37484
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 13900 36772 13940 36812
rect 7084 36688 7124 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7084 36016 7124 36056
rect 2380 35848 2420 35888
rect 940 35428 980 35468
rect 652 24928 692 24968
rect 652 24088 692 24128
rect 652 23248 692 23288
rect 652 22408 692 22448
rect 652 21568 692 21608
rect 652 20728 692 20768
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 652 15688 692 15728
rect 652 14008 692 14048
rect 652 13168 692 13208
rect 652 11488 692 11528
rect 652 10732 692 10772
rect 652 9808 692 9848
rect 652 8968 692 9008
rect 556 8128 596 8168
rect 652 7288 692 7328
rect 652 6448 692 6488
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 652 3928 692 3968
rect 844 24760 884 24800
rect 844 24004 884 24044
rect 2284 18628 2324 18668
rect 2188 18544 2228 18584
rect 2092 17284 2132 17324
rect 1324 17200 1364 17240
rect 1804 16444 1844 16484
rect 1228 15436 1268 15476
rect 844 15352 884 15392
rect 1036 14848 1076 14888
rect 2284 17200 2324 17240
rect 1516 15352 1556 15392
rect 1612 14848 1652 14888
rect 1900 14848 1940 14888
rect 1228 13168 1268 13208
rect 1420 13168 1460 13208
rect 844 12580 884 12620
rect 1036 12328 1076 12368
rect 844 10900 884 10940
rect 844 10228 884 10268
rect 844 9388 884 9428
rect 940 5440 980 5480
rect 1420 12580 1460 12620
rect 2092 14680 2132 14720
rect 1996 13000 2036 13040
rect 1804 12496 1844 12536
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4972 34504 5012 34544
rect 4876 34168 4916 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 4588 32320 4628 32360
rect 2956 32068 2996 32108
rect 4396 32068 4436 32108
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 3820 31312 3860 31352
rect 4588 31312 4628 31352
rect 5740 34336 5780 34376
rect 5164 34000 5204 34040
rect 4972 32320 5012 32360
rect 5548 32908 5588 32948
rect 5260 32572 5300 32612
rect 3436 30472 3476 30512
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 4492 30724 4532 30764
rect 4588 30640 4628 30680
rect 4204 30472 4244 30512
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 4492 29044 4532 29084
rect 3820 28960 3860 29000
rect 3436 28876 3476 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3436 26104 3476 26144
rect 4492 28120 4532 28160
rect 4876 29044 4916 29084
rect 4876 28876 4916 28916
rect 4780 28288 4820 28328
rect 4876 28204 4916 28244
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3628 25936 3668 25976
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 3436 23668 3476 23708
rect 3532 23080 3572 23120
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 3340 22408 3380 22448
rect 4204 26104 4244 26144
rect 4876 27952 4916 27992
rect 4492 25852 4532 25892
rect 4588 25264 4628 25304
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3628 22408 3668 22448
rect 4204 23668 4244 23708
rect 3916 23332 3956 23372
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3340 21652 3380 21692
rect 3436 21568 3476 21608
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4876 23500 4916 23540
rect 4588 23248 4628 23288
rect 4492 23164 4532 23204
rect 4588 23080 4628 23120
rect 4780 23080 4820 23120
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 3916 19972 3956 20012
rect 2956 19048 2996 19088
rect 2572 18544 2612 18584
rect 4204 20728 4244 20768
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 4012 19888 4052 19928
rect 4012 19048 4052 19088
rect 3244 18628 3284 18668
rect 2572 17872 2612 17912
rect 2860 17872 2900 17912
rect 2476 17788 2516 17828
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 3916 18544 3956 18584
rect 3820 17788 3860 17828
rect 3052 17200 3092 17240
rect 3916 17284 3956 17324
rect 3916 16864 3956 16904
rect 2572 16444 2612 16484
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 3244 16444 3284 16484
rect 3916 16444 3956 16484
rect 3436 15436 3476 15476
rect 2956 15352 2996 15392
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 3244 14848 3284 14888
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 3820 14512 3860 14552
rect 3724 13168 3764 13208
rect 2572 13000 2612 13040
rect 1708 12244 1748 12284
rect 1804 10900 1844 10940
rect 1900 10228 1940 10268
rect 1804 6700 1844 6740
rect 2476 12496 2516 12536
rect 2764 12748 2804 12788
rect 2956 12328 2996 12368
rect 3244 12244 3284 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3916 12664 3956 12704
rect 3916 12328 3956 12368
rect 3724 11488 3764 11528
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 2668 10144 2708 10184
rect 2956 10144 2996 10184
rect 4300 19888 4340 19928
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 4204 18544 4244 18584
rect 4684 18544 4724 18584
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4659 17260 4699 17300
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4204 15436 4244 15476
rect 4108 15352 4148 15392
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 3436 7960 3476 8000
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 2188 7120 2228 7160
rect 1900 6616 1940 6656
rect 1420 6448 1460 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 1132 5524 1172 5564
rect 1036 4768 1076 4808
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4492 15604 4532 15644
rect 4588 15520 4628 15560
rect 4684 14680 4724 14720
rect 4588 14512 4628 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 4204 14176 4244 14216
rect 4684 13168 4724 13208
rect 4204 13000 4244 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 4300 11656 4340 11696
rect 4684 11488 4724 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 4588 10144 4628 10184
rect 4204 10060 4244 10100
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 5068 30640 5108 30680
rect 5164 29128 5204 29168
rect 5068 25264 5108 25304
rect 5164 24004 5204 24044
rect 5164 23332 5204 23372
rect 6412 32404 6452 32444
rect 5356 32068 5396 32108
rect 5836 31564 5876 31604
rect 5932 31480 5972 31520
rect 5836 30724 5876 30764
rect 5836 29128 5876 29168
rect 5452 28960 5492 29000
rect 5356 28204 5396 28244
rect 5260 23164 5300 23204
rect 5836 25852 5876 25892
rect 5836 24004 5876 24044
rect 5740 23332 5780 23372
rect 5068 21904 5108 21944
rect 4972 20728 5012 20768
rect 5068 19972 5108 20012
rect 4972 18628 5012 18668
rect 5068 17872 5108 17912
rect 4876 14680 4916 14720
rect 5068 14176 5108 14216
rect 4876 13168 4916 13208
rect 4972 12496 5012 12536
rect 4876 11488 4916 11528
rect 4972 10144 5012 10184
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 4588 8128 4628 8168
rect 4300 7960 4340 8000
rect 4684 7960 4724 8000
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 4780 5356 4820 5396
rect 5356 21652 5396 21692
rect 5836 23248 5876 23288
rect 5740 20896 5780 20936
rect 5836 19972 5876 20012
rect 5836 19048 5876 19088
rect 5932 18880 5972 18920
rect 5836 16696 5876 16736
rect 5932 16528 5972 16568
rect 5836 15604 5876 15644
rect 5932 15520 5972 15560
rect 6412 14680 6452 14720
rect 5740 12748 5780 12788
rect 5260 11992 5300 12032
rect 5260 11656 5300 11696
rect 5164 10144 5204 10184
rect 5836 12664 5876 12704
rect 5836 12328 5876 12368
rect 5836 10060 5876 10100
rect 5740 8128 5780 8168
rect 5164 7960 5204 8000
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 5068 5272 5108 5312
rect 5932 6952 5972 6992
rect 18700 36688 18740 36728
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 13804 35680 13844 35720
rect 8140 35596 8180 35636
rect 7276 34504 7316 34544
rect 7564 34504 7604 34544
rect 7852 34336 7892 34376
rect 7372 34168 7412 34208
rect 7276 34084 7316 34124
rect 7948 33664 7988 33704
rect 7948 7036 7988 7076
rect 7084 4936 7124 4976
rect 10636 35092 10676 35132
rect 10252 34168 10292 34208
rect 9964 34000 10004 34040
rect 8332 33916 8372 33956
rect 8236 33832 8276 33872
rect 8140 4264 8180 4304
rect 5164 4096 5204 4136
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 4108 3676 4148 3716
rect 8236 3424 8276 3464
rect 748 3340 788 3380
rect 652 3088 692 3128
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 10636 34840 10676 34880
rect 12076 34504 12116 34544
rect 12940 34504 12980 34544
rect 13420 34504 13460 34544
rect 11212 34084 11252 34124
rect 13324 34168 13364 34208
rect 13612 35176 13652 35216
rect 10444 34000 10484 34040
rect 13228 34000 13268 34040
rect 13516 34000 13556 34040
rect 10348 33748 10388 33788
rect 13228 33748 13268 33788
rect 14188 35848 14228 35888
rect 16204 35848 16244 35888
rect 14092 35680 14132 35720
rect 15340 35680 15380 35720
rect 14092 35176 14132 35216
rect 14668 35176 14708 35216
rect 14476 35008 14516 35048
rect 16204 35176 16244 35216
rect 15340 34924 15380 34964
rect 14380 34168 14420 34208
rect 15820 34168 15860 34208
rect 16012 34000 16052 34040
rect 15820 33748 15860 33788
rect 16012 33664 16052 33704
rect 13900 32068 13940 32108
rect 15161 31564 15201 31604
rect 16588 34588 16628 34628
rect 18508 35848 18548 35888
rect 17548 35764 17588 35804
rect 18892 35764 18932 35804
rect 18796 35680 18836 35720
rect 18124 35176 18164 35216
rect 18700 35176 18740 35216
rect 17452 35092 17492 35132
rect 17260 35008 17300 35048
rect 17356 34756 17396 34796
rect 18028 34756 18068 34796
rect 19084 35848 19124 35888
rect 18988 35092 19028 35132
rect 19660 35848 19700 35888
rect 19948 35848 19988 35888
rect 19276 35512 19316 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 19084 35008 19124 35048
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 20044 35680 20084 35720
rect 19564 35092 19604 35132
rect 20140 35176 20180 35216
rect 20524 36688 20564 36728
rect 21004 37360 21044 37400
rect 20620 35848 20660 35888
rect 21388 36520 21428 36560
rect 20908 35848 20948 35888
rect 20908 35344 20948 35384
rect 21100 35344 21140 35384
rect 20524 35176 20564 35216
rect 20140 35008 20180 35048
rect 20044 34924 20084 34964
rect 20332 34840 20372 34880
rect 19276 34588 19316 34628
rect 19564 34420 19604 34460
rect 21100 35092 21140 35132
rect 21772 37360 21812 37400
rect 21868 36688 21908 36728
rect 21676 36520 21716 36560
rect 21772 36184 21812 36224
rect 22252 37360 22292 37400
rect 22348 37192 22388 37232
rect 22540 37276 22580 37316
rect 22444 36604 22484 36644
rect 22540 36520 22580 36560
rect 22444 36184 22484 36224
rect 21580 35344 21620 35384
rect 21964 35176 22004 35216
rect 21388 35008 21428 35048
rect 22636 35764 22676 35804
rect 23404 37192 23444 37232
rect 23116 37024 23156 37064
rect 23020 36688 23060 36728
rect 23884 37948 23924 37988
rect 24652 37948 24692 37988
rect 24460 37528 24500 37568
rect 24556 37360 24596 37400
rect 24844 37360 24884 37400
rect 24172 37192 24212 37232
rect 23788 37108 23828 37148
rect 24076 37108 24116 37148
rect 23692 36772 23732 36812
rect 23308 36436 23348 36476
rect 22732 35008 22772 35048
rect 21292 34420 21332 34460
rect 22540 34420 22580 34460
rect 22252 34336 22292 34376
rect 23980 37024 24020 37064
rect 24460 36940 24500 36980
rect 24172 36856 24212 36896
rect 23884 36604 23924 36644
rect 25612 37024 25652 37064
rect 24844 36856 24884 36896
rect 25132 36856 25172 36896
rect 25516 36856 25556 36896
rect 25996 37024 26036 37064
rect 24652 36772 24692 36812
rect 25324 36772 25364 36812
rect 24940 36688 24980 36728
rect 25708 36688 25748 36728
rect 25612 36604 25652 36644
rect 24652 36436 24692 36476
rect 26668 37780 26708 37820
rect 26092 36940 26132 36980
rect 25996 36604 26036 36644
rect 23116 34924 23156 34964
rect 23788 34924 23828 34964
rect 21004 34252 21044 34292
rect 18796 34168 18836 34208
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 25036 35848 25076 35888
rect 26380 36772 26420 36812
rect 26668 37108 26708 37148
rect 27532 37276 27572 37316
rect 27724 37780 27764 37820
rect 27628 37192 27668 37232
rect 27436 37108 27476 37148
rect 26860 37024 26900 37064
rect 27244 37024 27284 37064
rect 26476 36268 26516 36308
rect 25036 34588 25076 34628
rect 24364 34336 24404 34376
rect 25516 34336 25556 34376
rect 25228 33916 25268 33956
rect 27340 36940 27380 36980
rect 27244 36772 27284 36812
rect 27148 36604 27188 36644
rect 27532 36604 27572 36644
rect 27436 36520 27476 36560
rect 26860 36268 26900 36308
rect 26764 36184 26804 36224
rect 27100 35848 27140 35888
rect 27820 36940 27860 36980
rect 27820 36520 27860 36560
rect 27724 36184 27764 36224
rect 29260 38200 29300 38240
rect 29260 37780 29300 37820
rect 28108 37360 28148 37400
rect 28972 37360 29012 37400
rect 28012 37108 28052 37148
rect 28204 37024 28244 37064
rect 28012 36688 28052 36728
rect 28012 36436 28052 36476
rect 28108 36184 28148 36224
rect 29740 38200 29780 38240
rect 30412 37528 30452 37568
rect 32908 37528 32948 37568
rect 29932 37360 29972 37400
rect 29740 37192 29780 37232
rect 30028 37024 30068 37064
rect 29260 36688 29300 36728
rect 30028 36688 30068 36728
rect 28972 36436 29012 36476
rect 28492 36184 28532 36224
rect 26284 34840 26324 34880
rect 26476 34672 26516 34712
rect 26764 34672 26804 34712
rect 27340 34588 27380 34628
rect 27052 34336 27092 34376
rect 28876 34588 28916 34628
rect 30892 37360 30932 37400
rect 31468 37360 31508 37400
rect 30604 36688 30644 36728
rect 32044 37276 32084 37316
rect 32620 37192 32660 37232
rect 31564 36436 31604 36476
rect 31948 36184 31988 36224
rect 30892 34672 30932 34712
rect 29548 34336 29588 34376
rect 30508 34336 30548 34376
rect 27148 34252 27188 34292
rect 26188 33832 26228 33872
rect 23980 33748 24020 33788
rect 29740 34252 29780 34292
rect 30028 34252 30068 34292
rect 31276 34588 31316 34628
rect 32332 36436 32372 36476
rect 33100 37192 33140 37232
rect 33292 38200 33332 38240
rect 33868 38200 33908 38240
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 32908 36520 32948 36560
rect 32524 36016 32564 36056
rect 31852 35092 31892 35132
rect 31564 34336 31604 34376
rect 32044 34336 32084 34376
rect 32524 34840 32564 34880
rect 32428 34336 32468 34376
rect 32812 35092 32852 35132
rect 32716 34672 32756 34712
rect 30604 34252 30644 34292
rect 31660 34168 31700 34208
rect 30220 34084 30260 34124
rect 17548 31648 17588 31688
rect 16313 31480 16353 31520
rect 16492 31480 16532 31520
rect 18233 31648 18273 31688
rect 33004 36184 33044 36224
rect 32908 34840 32948 34880
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 33964 37948 34004 37988
rect 35692 37948 35732 37988
rect 34444 37360 34484 37400
rect 33964 37276 34004 37316
rect 33868 36436 33908 36476
rect 33772 36100 33812 36140
rect 33388 35932 33428 35972
rect 33388 35428 33428 35468
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 36556 37360 36596 37400
rect 35308 37192 35348 37232
rect 36460 37192 36500 37232
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 33388 34588 33428 34628
rect 33964 34588 34004 34628
rect 35116 36184 35156 36224
rect 34924 35932 34964 35972
rect 35692 36688 35732 36728
rect 35692 36436 35732 36476
rect 35500 36016 35540 36056
rect 35308 35932 35348 35972
rect 35692 35848 35732 35888
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 34540 35176 34580 35216
rect 35404 35596 35444 35636
rect 35212 35260 35252 35300
rect 35116 35008 35156 35048
rect 35404 35008 35444 35048
rect 36364 36016 36404 36056
rect 36076 35932 36116 35972
rect 36172 35848 36212 35888
rect 35788 35428 35828 35468
rect 35788 35260 35828 35300
rect 36172 35428 36212 35468
rect 36172 35092 36212 35132
rect 35692 34840 35732 34880
rect 36364 35008 36404 35048
rect 36364 34756 36404 34796
rect 36268 34672 36308 34712
rect 35692 34504 35732 34544
rect 34348 34336 34388 34376
rect 34540 34168 34580 34208
rect 33196 34000 33236 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 35212 32572 35252 32612
rect 36844 37192 36884 37232
rect 37420 37360 37460 37400
rect 36940 36688 36980 36728
rect 37132 35932 37172 35972
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 44044 37444 44084 37484
rect 38380 37360 38420 37400
rect 38572 37360 38612 37400
rect 37804 36856 37844 36896
rect 39628 36688 39668 36728
rect 37804 36352 37844 36392
rect 39628 36352 39668 36392
rect 37708 36016 37748 36056
rect 39148 36016 39188 36056
rect 37516 35848 37556 35888
rect 38380 35596 38420 35636
rect 37228 35176 37268 35216
rect 36940 34756 36980 34796
rect 36556 34168 36596 34208
rect 36652 34084 36692 34124
rect 38092 34504 38132 34544
rect 39916 37192 39956 37232
rect 40108 36688 40148 36728
rect 41068 36688 41108 36728
rect 39724 35848 39764 35888
rect 40012 35848 40052 35888
rect 40972 36604 41012 36644
rect 40300 36520 40340 36560
rect 40300 35848 40340 35888
rect 40204 35764 40244 35804
rect 40396 35764 40436 35804
rect 42796 36688 42836 36728
rect 42316 36520 42356 36560
rect 41932 36436 41972 36476
rect 41164 36016 41204 36056
rect 40588 35512 40628 35552
rect 41356 35848 41396 35888
rect 41260 35764 41300 35804
rect 42124 35092 42164 35132
rect 42796 35092 42836 35132
rect 36940 33916 36980 33956
rect 36652 33832 36692 33872
rect 36460 32488 36500 32528
rect 38092 34168 38132 34208
rect 43276 35764 43316 35804
rect 43084 34924 43124 34964
rect 38764 33916 38804 33956
rect 40300 33916 40340 33956
rect 42220 34168 42260 34208
rect 43660 35764 43700 35804
rect 43468 34924 43508 34964
rect 69292 37360 69332 37400
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 44524 35932 44564 35972
rect 43852 35848 43892 35888
rect 45868 35848 45908 35888
rect 44140 35764 44180 35804
rect 45580 35764 45620 35804
rect 43948 35680 43988 35720
rect 44716 35680 44756 35720
rect 44332 35428 44372 35468
rect 44140 35176 44180 35216
rect 45484 35092 45524 35132
rect 43372 34000 43412 34040
rect 41164 33832 41204 33872
rect 43276 33832 43316 33872
rect 45196 34336 45236 34376
rect 47980 36016 48020 36056
rect 47020 35848 47060 35888
rect 47212 35848 47252 35888
rect 45964 35428 46004 35468
rect 46348 35176 46388 35216
rect 47308 35176 47348 35216
rect 47308 35008 47348 35048
rect 47212 34924 47252 34964
rect 47020 34672 47060 34712
rect 46348 34000 46388 34040
rect 48940 35848 48980 35888
rect 48172 35008 48212 35048
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 48076 34672 48116 34712
rect 46924 33916 46964 33956
rect 45580 32656 45620 32696
rect 37612 32404 37652 32444
rect 43660 32404 43700 32444
rect 49324 35596 49364 35636
rect 50668 35848 50708 35888
rect 50956 35764 50996 35804
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 50764 35008 50804 35048
rect 49900 34924 49940 34964
rect 49900 34756 49940 34796
rect 49324 34672 49364 34712
rect 49420 34504 49460 34544
rect 49612 34504 49652 34544
rect 48940 34000 48980 34040
rect 49228 34000 49268 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 49420 33832 49460 33872
rect 49132 33580 49172 33620
rect 50860 34168 50900 34208
rect 50860 34000 50900 34040
rect 51628 35848 51668 35888
rect 52012 35764 52052 35804
rect 51916 35596 51956 35636
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 52012 34924 52052 34964
rect 51916 34840 51956 34880
rect 53356 35008 53396 35048
rect 54028 35008 54068 35048
rect 64396 35008 64436 35048
rect 53836 34924 53876 34964
rect 52972 34840 53012 34880
rect 52492 34756 52532 34796
rect 51340 33664 51380 33704
rect 51052 33580 51092 33620
rect 52300 34168 52340 34208
rect 52492 34000 52532 34040
rect 52300 33832 52340 33872
rect 52780 33664 52820 33704
rect 52012 32572 52052 32612
rect 50380 31732 50420 31772
rect 53164 34756 53204 34796
rect 53164 33748 53204 33788
rect 54508 34924 54548 34964
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 65452 35176 65492 35216
rect 54028 33832 54068 33872
rect 64204 34336 64244 34376
rect 64588 34336 64628 34376
rect 62764 34168 62804 34208
rect 61516 34000 61556 34040
rect 62476 34000 62516 34040
rect 68044 34504 68084 34544
rect 66316 34336 66356 34376
rect 68908 34336 68948 34376
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 92428 36940 92468 36980
rect 81580 36772 81620 36812
rect 91025 36772 91065 36812
rect 80428 36688 80468 36728
rect 71980 36436 72020 36476
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 71404 36016 71444 36056
rect 71980 36016 72020 36056
rect 70156 35092 70196 35132
rect 70924 35092 70964 35132
rect 70156 34336 70196 34376
rect 70636 34336 70676 34376
rect 68524 34168 68564 34208
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 64588 33832 64628 33872
rect 61516 33664 61556 33704
rect 64396 33664 64436 33704
rect 55180 33580 55220 33620
rect 17452 6784 17492 6824
rect 18700 5608 18740 5648
rect 17932 5272 17972 5312
rect 18700 5356 18740 5396
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 18316 4684 18356 4724
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 18508 4180 18548 4220
rect 18700 4180 18740 4220
rect 19276 4180 19316 4220
rect 18124 4096 18164 4136
rect 17356 4012 17396 4052
rect 17260 3928 17300 3968
rect 20428 4096 20468 4136
rect 19564 4012 19604 4052
rect 18508 3928 18548 3968
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 17356 3676 17396 3716
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 8332 2836 8372 2876
rect 21580 5608 21620 5648
rect 21100 4684 21140 4724
rect 20908 4180 20948 4220
rect 20716 4012 20756 4052
rect 20620 2752 20660 2792
rect 20524 2668 20564 2708
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 20908 3928 20948 3968
rect 22636 4600 22676 4640
rect 22444 4180 22484 4220
rect 21772 4096 21812 4136
rect 21676 4012 21716 4052
rect 21580 3928 21620 3968
rect 21292 3256 21332 3296
rect 21484 2752 21524 2792
rect 22540 4096 22580 4136
rect 22444 3676 22484 3716
rect 21868 3256 21908 3296
rect 26332 7204 26372 7244
rect 23788 6952 23828 6992
rect 25612 7120 25652 7160
rect 23980 5608 24020 5648
rect 23692 5272 23732 5312
rect 24652 5272 24692 5312
rect 23308 5188 23348 5228
rect 31756 6448 31796 6488
rect 29260 5692 29300 5732
rect 26284 5356 26324 5396
rect 24748 5188 24788 5228
rect 22924 4600 22964 4640
rect 23212 3928 23252 3968
rect 24364 4684 24404 4724
rect 24748 4684 24788 4724
rect 24652 4180 24692 4220
rect 25036 4600 25076 4640
rect 24844 4516 24884 4556
rect 23692 3928 23732 3968
rect 23692 3508 23732 3548
rect 24556 3424 24596 3464
rect 22732 2752 22772 2792
rect 23500 2668 23540 2708
rect 24268 2668 24308 2708
rect 25708 4516 25748 4556
rect 25132 4096 25172 4136
rect 25612 4096 25652 4136
rect 25516 3508 25556 3548
rect 25996 2836 26036 2876
rect 24652 1996 24692 2036
rect 25036 1996 25076 2036
rect 24364 1912 24404 1952
rect 26284 4600 26324 4640
rect 27148 4180 27188 4220
rect 27436 4180 27476 4220
rect 27724 4096 27764 4136
rect 27244 3508 27284 3548
rect 27244 2920 27284 2960
rect 27148 2584 27188 2624
rect 27148 1996 27188 2036
rect 26092 1828 26132 1868
rect 23980 1744 24020 1784
rect 25900 1744 25940 1784
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 26956 1912 26996 1952
rect 26956 1660 26996 1700
rect 28588 3424 28628 3464
rect 27724 2920 27764 2960
rect 28108 2836 28148 2876
rect 27628 2584 27668 2624
rect 28012 2584 28052 2624
rect 28108 1996 28148 2036
rect 28300 1660 28340 1700
rect 28780 2920 28820 2960
rect 28588 1912 28628 1952
rect 28396 1324 28436 1364
rect 31660 4348 31700 4388
rect 29932 4012 29972 4052
rect 29740 3844 29780 3884
rect 29740 3508 29780 3548
rect 33772 7036 33812 7076
rect 33388 6784 33428 6824
rect 32716 5356 32756 5396
rect 32716 4768 32756 4808
rect 32908 4768 32948 4808
rect 32044 4684 32084 4724
rect 32428 4684 32468 4724
rect 32140 4348 32180 4388
rect 31756 3928 31796 3968
rect 32620 4096 32660 4136
rect 33100 4096 33140 4136
rect 32236 3676 32276 3716
rect 32140 3424 32180 3464
rect 30412 3172 30452 3212
rect 31180 3172 31220 3212
rect 30700 2584 30740 2624
rect 30316 2080 30356 2120
rect 32044 2080 32084 2120
rect 29740 1996 29780 2036
rect 30892 1996 30932 2036
rect 29260 1744 29300 1784
rect 30028 1828 30068 1868
rect 30796 1324 30836 1364
rect 33292 4768 33332 4808
rect 33484 4768 33524 4808
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 33196 3928 33236 3968
rect 32716 3592 32756 3632
rect 33100 3592 33140 3632
rect 32620 3340 32660 3380
rect 32620 2920 32660 2960
rect 32524 2080 32564 2120
rect 34060 3592 34100 3632
rect 34636 5608 34676 5648
rect 34924 5692 34964 5732
rect 35020 5608 35060 5648
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 35116 5524 35156 5564
rect 34444 4768 34484 4808
rect 34444 4348 34484 4388
rect 34636 4432 34676 4472
rect 35404 5776 35444 5816
rect 36172 6532 36212 6572
rect 35212 5272 35252 5312
rect 35020 4768 35060 4808
rect 35212 4684 35252 4724
rect 34540 4180 34580 4220
rect 34924 4264 34964 4304
rect 34828 4096 34868 4136
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 33868 3508 33908 3548
rect 34348 3508 34388 3548
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 33196 2584 33236 2624
rect 33484 2584 33524 2624
rect 33484 1912 33524 1952
rect 32332 1660 32372 1700
rect 32428 1072 32468 1112
rect 34828 2584 34868 2624
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 34636 2080 34676 2120
rect 35116 4096 35156 4136
rect 33964 1828 34004 1868
rect 34636 1660 34676 1700
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 35404 5440 35444 5480
rect 35788 5188 35828 5228
rect 35980 5104 36020 5144
rect 35500 4768 35540 4808
rect 35596 4432 35636 4472
rect 36076 4348 36116 4388
rect 35596 4264 35636 4304
rect 35404 4096 35444 4136
rect 36172 4264 36212 4304
rect 36076 4012 36116 4052
rect 37516 7036 37556 7076
rect 37900 7036 37940 7076
rect 37612 6784 37652 6824
rect 37612 6616 37652 6656
rect 36940 4768 36980 4808
rect 39436 5104 39476 5144
rect 37804 4768 37844 4808
rect 36748 4096 36788 4136
rect 37036 4180 37076 4220
rect 36844 4012 36884 4052
rect 35788 3676 35828 3716
rect 35692 3592 35732 3632
rect 35884 3592 35924 3632
rect 35404 2080 35444 2120
rect 35212 1744 35252 1784
rect 35116 1324 35156 1364
rect 35020 1072 35060 1112
rect 35308 1072 35348 1112
rect 32524 988 32564 1028
rect 32716 988 32756 1028
rect 34924 988 34964 1028
rect 35788 3508 35828 3548
rect 35692 3004 35732 3044
rect 36076 2584 36116 2624
rect 37516 4096 37556 4136
rect 37612 4012 37652 4052
rect 37708 3928 37748 3968
rect 37132 3760 37172 3800
rect 39244 4768 39284 4808
rect 38860 4096 38900 4136
rect 39148 3928 39188 3968
rect 37996 3760 38036 3800
rect 39052 3760 39092 3800
rect 39148 3424 39188 3464
rect 37708 3340 37748 3380
rect 39052 3004 39092 3044
rect 37900 2584 37940 2624
rect 38860 2584 38900 2624
rect 38188 2500 38228 2540
rect 37900 1996 37940 2036
rect 36940 1917 36980 1952
rect 36940 1912 36980 1917
rect 36748 1408 36788 1448
rect 37708 1660 37748 1700
rect 35596 1324 35636 1364
rect 37324 1324 37364 1364
rect 38572 1660 38612 1700
rect 38476 1072 38516 1112
rect 39628 3928 39668 3968
rect 39532 3844 39572 3884
rect 39532 3424 39572 3464
rect 39436 2668 39476 2708
rect 40012 4012 40052 4052
rect 40108 3676 40148 3716
rect 40889 7288 40929 7328
rect 40780 6280 40820 6320
rect 40588 5440 40628 5480
rect 40684 4768 40724 4808
rect 40492 4180 40532 4220
rect 39916 3424 39956 3464
rect 39724 2584 39764 2624
rect 40108 2584 40148 2624
rect 39628 2500 39668 2540
rect 39820 2500 39860 2540
rect 39724 1828 39764 1868
rect 39244 1576 39284 1616
rect 38860 1324 38900 1364
rect 40108 1324 40148 1364
rect 40588 1912 40628 1952
rect 40876 4600 40916 4640
rect 40876 3928 40916 3968
rect 41068 6280 41108 6320
rect 42892 4936 42932 4976
rect 41932 4684 41972 4724
rect 42220 4684 42260 4724
rect 41164 4096 41204 4136
rect 41740 4096 41780 4136
rect 42412 4432 42452 4472
rect 42316 4180 42356 4220
rect 40972 3508 41012 3548
rect 42220 4012 42260 4052
rect 42892 4012 42932 4052
rect 44524 6448 44564 6488
rect 46348 5020 46388 5060
rect 43852 4936 43892 4976
rect 45196 4852 45236 4892
rect 43852 4684 43892 4724
rect 43180 3928 43220 3968
rect 41356 2584 41396 2624
rect 40972 2500 41012 2540
rect 41356 2080 41396 2120
rect 41260 1912 41300 1952
rect 40684 1156 40724 1196
rect 40204 1072 40244 1112
rect 40492 1072 40532 1112
rect 44140 4180 44180 4220
rect 45196 4180 45236 4220
rect 45388 4180 45428 4220
rect 44044 4096 44084 4136
rect 46348 4180 46388 4220
rect 44236 3508 44276 3548
rect 44716 3508 44756 3548
rect 43084 3424 43124 3464
rect 44524 3424 44564 3464
rect 43852 2668 43892 2708
rect 44236 2080 44276 2120
rect 43948 1996 43988 2036
rect 44140 1996 44180 2036
rect 43084 1912 43124 1952
rect 42220 1828 42260 1868
rect 44908 2668 44948 2708
rect 45100 2668 45140 2708
rect 45196 1996 45236 2036
rect 46732 4936 46772 4976
rect 46828 4432 46868 4472
rect 46732 4180 46772 4220
rect 46732 4012 46772 4052
rect 46444 3004 46484 3044
rect 46156 2920 46196 2960
rect 46732 2920 46772 2960
rect 45292 1912 45332 1952
rect 45868 1912 45908 1952
rect 44812 1408 44852 1448
rect 42604 1072 42644 1112
rect 44332 1072 44372 1112
rect 46252 2164 46292 2204
rect 46252 1912 46292 1952
rect 46540 1072 46580 1112
rect 47116 4348 47156 4388
rect 46924 3676 46964 3716
rect 47116 3424 47156 3464
rect 47116 2920 47156 2960
rect 47308 3508 47348 3548
rect 79180 35680 79220 35720
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 74188 33832 74228 33872
rect 72652 32572 72692 32612
rect 71404 7120 71444 7160
rect 49036 6700 49076 6740
rect 47596 5020 47636 5060
rect 48364 5020 48404 5060
rect 47980 4936 48020 4976
rect 48076 4852 48116 4892
rect 48076 4348 48116 4388
rect 47788 3340 47828 3380
rect 47404 2584 47444 2624
rect 47212 2164 47252 2204
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 48364 3424 48404 3464
rect 48940 4012 48980 4052
rect 49612 6196 49652 6236
rect 49420 5356 49460 5396
rect 49516 4936 49556 4976
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 78508 32656 78548 32696
rect 75820 17956 75860 17996
rect 78412 16780 78452 16820
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 81484 35008 81524 35048
rect 80908 33832 80948 33872
rect 80812 33160 80852 33200
rect 80140 32656 80180 32696
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 79180 31648 79220 31688
rect 80332 31396 80372 31436
rect 78604 30556 78644 30596
rect 79180 30556 79220 30596
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 79660 30136 79700 30176
rect 78796 28960 78836 29000
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 80044 30808 80084 30848
rect 80044 30220 80084 30260
rect 79948 30136 79988 30176
rect 81196 32656 81236 32696
rect 81100 31312 81140 31352
rect 81004 31060 81044 31100
rect 80716 30808 80756 30848
rect 80620 30136 80660 30176
rect 80620 29632 80660 29672
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 79372 28960 79412 29000
rect 79180 28876 79220 28916
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 80332 28708 80372 28748
rect 79756 27700 79796 27740
rect 80236 28288 80276 28328
rect 81388 31396 81428 31436
rect 80812 29212 80852 29252
rect 81388 30472 81428 30512
rect 81196 29632 81236 29672
rect 81388 29212 81428 29252
rect 81196 28876 81236 28916
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 80140 26860 80180 26900
rect 80524 27700 80564 27740
rect 80524 26860 80564 26900
rect 80140 26692 80180 26732
rect 80428 26692 80468 26732
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 80620 26104 80660 26144
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 80620 25432 80660 25472
rect 83308 36604 83348 36644
rect 82060 34252 82100 34292
rect 82252 34084 82292 34124
rect 81868 32656 81908 32696
rect 81964 31648 82004 31688
rect 81676 31312 81716 31352
rect 82060 30472 82100 30512
rect 81772 30220 81812 30260
rect 81676 29800 81716 29840
rect 81580 28288 81620 28328
rect 81196 26104 81236 26144
rect 81292 25600 81332 25640
rect 80524 25180 80564 25220
rect 80620 25096 80660 25136
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 80908 25264 80948 25304
rect 80620 23668 80660 23708
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 79468 20728 79508 20768
rect 81196 23668 81236 23708
rect 81676 25600 81716 25640
rect 83116 33160 83156 33200
rect 83212 31060 83252 31100
rect 83116 30892 83156 30932
rect 82924 30808 82964 30848
rect 92177 36688 92217 36728
rect 92753 36856 92793 36896
rect 83308 29800 83348 29840
rect 83212 28708 83252 28748
rect 83308 28204 83348 28244
rect 83308 27700 83348 27740
rect 82636 26692 82676 26732
rect 81580 25180 81620 25220
rect 81580 24508 81620 24548
rect 81868 25264 81908 25304
rect 82636 24424 82676 24464
rect 82732 24340 82772 24380
rect 81676 24004 81716 24044
rect 83212 24004 83252 24044
rect 81484 23752 81524 23792
rect 82060 23752 82100 23792
rect 81484 20980 81524 21020
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 78508 16192 78548 16232
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 78508 6448 78548 6488
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 72652 5440 72692 5480
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 52204 5188 52244 5228
rect 49996 5104 50036 5144
rect 49708 4684 49748 4724
rect 49228 4264 49268 4304
rect 49228 3760 49268 3800
rect 49324 3592 49364 3632
rect 92572 24424 92612 24464
rect 90460 24340 90500 24380
rect 87916 24004 87956 24044
rect 82444 23668 82484 23708
rect 85420 23668 85460 23708
rect 82060 20812 82100 20852
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 84460 20980 84500 21020
rect 83308 20728 83348 20768
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 82732 20056 82772 20096
rect 96748 20056 96788 20096
rect 80620 16780 80660 16820
rect 81388 16780 81428 16820
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 81388 9220 81428 9260
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 98572 19888 98612 19928
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 98860 17956 98900 17996
rect 98860 9379 98900 9419
rect 82732 7036 82772 7076
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 80524 6616 80564 6656
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 53932 5020 53972 5060
rect 79468 5020 79508 5060
rect 50380 4768 50420 4808
rect 49900 4264 49940 4304
rect 49612 4096 49652 4136
rect 49804 4096 49844 4136
rect 49228 3508 49268 3548
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 48172 2584 48212 2624
rect 48364 2584 48404 2624
rect 47500 1996 47540 2036
rect 48940 2164 48980 2204
rect 48460 1996 48500 2036
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 47308 1408 47348 1448
rect 47788 1408 47828 1448
rect 47596 1072 47636 1112
rect 50188 4012 50228 4052
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 49708 3508 49748 3548
rect 49900 3508 49940 3548
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 52204 4432 52244 4472
rect 52396 4096 52436 4136
rect 50860 3676 50900 3716
rect 50764 3424 50804 3464
rect 50476 3340 50516 3380
rect 51532 4012 51572 4052
rect 52588 4852 52628 4892
rect 52492 3676 52532 3716
rect 53068 4012 53108 4052
rect 53548 3676 53588 3716
rect 55084 4852 55124 4892
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 80716 3592 80756 3632
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 50860 1996 50900 2036
rect 80908 3508 80948 3548
rect 80908 1828 80948 1868
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 80716 1492 80756 1532
rect 90537 1420 90577 1460
rect 90929 1439 90969 1479
rect 91121 1439 91161 1479
rect 91313 1439 91353 1479
rect 90729 1156 90769 1196
rect 50188 1072 50228 1112
rect 35500 988 35540 1028
rect 38188 988 38228 1028
rect 27052 904 27092 944
rect 28300 904 28340 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 29251 38200 29260 38240
rect 29300 38200 29740 38240
rect 29780 38200 29789 38240
rect 33283 38200 33292 38240
rect 33332 38200 33868 38240
rect 33908 38200 33917 38240
rect 5539 37988 5597 37989
rect 835 37948 844 37988
rect 884 37948 5548 37988
rect 5588 37948 5597 37988
rect 5539 37947 5597 37948
rect 8515 37988 8573 37989
rect 8515 37948 8524 37988
rect 8564 37948 23884 37988
rect 23924 37948 24652 37988
rect 24692 37948 24701 37988
rect 33955 37948 33964 37988
rect 34004 37948 35692 37988
rect 35732 37948 35741 37988
rect 8515 37947 8573 37948
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 26659 37780 26668 37820
rect 26708 37780 27724 37820
rect 27764 37780 29260 37820
rect 29300 37780 29309 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 0 37568 80 37588
rect 0 37528 652 37568
rect 692 37528 701 37568
rect 24451 37528 24460 37568
rect 24500 37528 30412 37568
rect 30452 37528 32908 37568
rect 32948 37528 32957 37568
rect 0 37508 80 37528
rect 19747 37444 19756 37484
rect 19796 37444 20428 37484
rect 20468 37444 44044 37484
rect 44084 37444 44093 37484
rect 20995 37360 21004 37400
rect 21044 37360 21772 37400
rect 21812 37360 21821 37400
rect 22243 37360 22252 37400
rect 22292 37360 24556 37400
rect 24596 37360 24844 37400
rect 24884 37360 28108 37400
rect 28148 37360 28157 37400
rect 28963 37360 28972 37400
rect 29012 37360 29932 37400
rect 29972 37360 29981 37400
rect 30883 37360 30892 37400
rect 30932 37360 31468 37400
rect 31508 37360 34444 37400
rect 34484 37360 34493 37400
rect 36547 37360 36556 37400
rect 36596 37360 37420 37400
rect 37460 37360 38380 37400
rect 38420 37360 38429 37400
rect 38563 37360 38572 37400
rect 38612 37360 69292 37400
rect 69332 37360 69341 37400
rect 29932 37316 29972 37360
rect 38572 37316 38612 37360
rect 22531 37276 22540 37316
rect 22580 37276 27532 37316
rect 27572 37276 27581 37316
rect 29932 37276 32044 37316
rect 32084 37276 32093 37316
rect 33955 37276 33964 37316
rect 34004 37276 38612 37316
rect 22339 37192 22348 37232
rect 22388 37192 23404 37232
rect 23444 37192 24172 37232
rect 24212 37192 24221 37232
rect 27619 37192 27628 37232
rect 27668 37192 29740 37232
rect 29780 37192 32620 37232
rect 32660 37192 32669 37232
rect 33091 37192 33100 37232
rect 33140 37192 35308 37232
rect 35348 37192 36460 37232
rect 36500 37192 36509 37232
rect 36835 37192 36844 37232
rect 36884 37192 39916 37232
rect 39956 37192 39965 37232
rect 23779 37108 23788 37148
rect 23828 37108 24076 37148
rect 24116 37108 26132 37148
rect 26659 37108 26668 37148
rect 26708 37108 27436 37148
rect 27476 37108 28012 37148
rect 28052 37108 28061 37148
rect 26092 37064 26132 37108
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 23107 37024 23116 37064
rect 23156 37024 23980 37064
rect 24020 37024 25612 37064
rect 25652 37024 25996 37064
rect 26036 37024 26045 37064
rect 26092 37024 26860 37064
rect 26900 37024 27244 37064
rect 27284 37024 28204 37064
rect 28244 37024 30028 37064
rect 30068 37024 30077 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 24451 36940 24460 36980
rect 24500 36940 26092 36980
rect 26132 36940 26141 36980
rect 27331 36940 27340 36980
rect 27380 36940 27820 36980
rect 27860 36940 27869 36980
rect 87820 36940 92428 36980
rect 92468 36940 92477 36980
rect 27340 36896 27380 36940
rect 24163 36856 24172 36896
rect 24212 36856 24844 36896
rect 24884 36856 24893 36896
rect 25123 36856 25132 36896
rect 25172 36856 25516 36896
rect 25556 36856 27380 36896
rect 33100 36856 37804 36896
rect 37844 36856 37853 36896
rect 33100 36812 33140 36856
rect 87820 36812 87860 36940
rect 13891 36772 13900 36812
rect 13940 36772 23692 36812
rect 23732 36772 23741 36812
rect 24643 36772 24652 36812
rect 24692 36772 25324 36812
rect 25364 36772 26380 36812
rect 26420 36772 26429 36812
rect 27235 36772 27244 36812
rect 27284 36772 33140 36812
rect 81571 36772 81580 36812
rect 81620 36772 87860 36812
rect 89356 36856 92753 36896
rect 92793 36856 92802 36896
rect 0 36728 80 36748
rect 27244 36728 27284 36772
rect 89356 36728 89396 36856
rect 0 36688 7084 36728
rect 7124 36688 7133 36728
rect 18691 36688 18700 36728
rect 18740 36688 20524 36728
rect 20564 36688 20573 36728
rect 21859 36688 21868 36728
rect 21908 36688 23020 36728
rect 23060 36688 23069 36728
rect 24931 36688 24940 36728
rect 24980 36688 25708 36728
rect 25748 36688 25757 36728
rect 25804 36688 27284 36728
rect 28003 36688 28012 36728
rect 28052 36688 29260 36728
rect 29300 36688 29309 36728
rect 30019 36688 30028 36728
rect 30068 36688 30604 36728
rect 30644 36688 30653 36728
rect 35683 36688 35692 36728
rect 35732 36688 36940 36728
rect 36980 36688 39628 36728
rect 39668 36688 39677 36728
rect 40099 36688 40108 36728
rect 40148 36688 41068 36728
rect 41108 36688 42796 36728
rect 42836 36688 42845 36728
rect 80419 36688 80428 36728
rect 80468 36688 89396 36728
rect 89452 36772 91025 36812
rect 91065 36772 91074 36812
rect 0 36668 80 36688
rect 25804 36644 25844 36688
rect 39628 36644 39668 36688
rect 89452 36644 89492 36772
rect 22435 36604 22444 36644
rect 22484 36604 23884 36644
rect 23924 36604 25612 36644
rect 25652 36604 25844 36644
rect 25987 36604 25996 36644
rect 26036 36604 27148 36644
rect 27188 36604 27532 36644
rect 27572 36604 27581 36644
rect 39628 36604 40972 36644
rect 41012 36604 41021 36644
rect 83299 36604 83308 36644
rect 83348 36604 89492 36644
rect 90028 36688 92177 36728
rect 92217 36688 92226 36728
rect 21379 36520 21388 36560
rect 21428 36520 21676 36560
rect 21716 36520 22540 36560
rect 22580 36520 22589 36560
rect 27427 36520 27436 36560
rect 27476 36520 27820 36560
rect 27860 36520 27869 36560
rect 32899 36520 32908 36560
rect 32948 36520 37460 36560
rect 40291 36520 40300 36560
rect 40340 36520 42316 36560
rect 42356 36520 42365 36560
rect 37420 36476 37460 36520
rect 90028 36476 90068 36688
rect 23299 36436 23308 36476
rect 23348 36436 24652 36476
rect 24692 36436 24701 36476
rect 28003 36436 28012 36476
rect 28052 36436 28972 36476
rect 29012 36436 29021 36476
rect 31555 36436 31564 36476
rect 31604 36436 32332 36476
rect 32372 36436 33868 36476
rect 33908 36436 35692 36476
rect 35732 36436 35741 36476
rect 37420 36436 41932 36476
rect 41972 36436 41981 36476
rect 71971 36436 71980 36476
rect 72020 36436 90068 36476
rect 37795 36352 37804 36392
rect 37844 36352 39628 36392
rect 39668 36352 39677 36392
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 26467 36268 26476 36308
rect 26516 36268 26860 36308
rect 26900 36268 26909 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 21763 36184 21772 36224
rect 21812 36184 22444 36224
rect 22484 36184 22493 36224
rect 26755 36184 26764 36224
rect 26804 36184 27724 36224
rect 27764 36184 28108 36224
rect 28148 36184 28492 36224
rect 28532 36184 28541 36224
rect 31939 36184 31948 36224
rect 31988 36184 33004 36224
rect 33044 36184 35116 36224
rect 35156 36184 35165 36224
rect 33772 36140 33812 36184
rect 33763 36100 33772 36140
rect 33812 36100 33821 36140
rect 7075 36016 7084 36056
rect 7124 36016 32524 36056
rect 32564 36016 32573 36056
rect 34828 36016 35500 36056
rect 35540 36016 35549 36056
rect 36355 36016 36364 36056
rect 36404 36016 37708 36056
rect 37748 36016 39148 36056
rect 39188 36016 41164 36056
rect 41204 36016 41213 36056
rect 47971 36016 47980 36056
rect 48020 36016 71404 36056
rect 71444 36016 71980 36056
rect 72020 36016 72029 36056
rect 34828 35972 34868 36016
rect 44515 35972 44573 35973
rect 33379 35932 33388 35972
rect 33428 35932 34868 35972
rect 34915 35932 34924 35972
rect 34964 35932 35308 35972
rect 35348 35932 35732 35972
rect 36067 35932 36076 35972
rect 36116 35932 37132 35972
rect 37172 35932 37460 35972
rect 44430 35932 44524 35972
rect 44564 35932 44573 35972
rect 0 35888 80 35908
rect 35692 35888 35732 35932
rect 37420 35888 37460 35932
rect 44515 35931 44573 35932
rect 69187 35888 69245 35889
rect 0 35848 2380 35888
rect 2420 35848 2429 35888
rect 14179 35848 14188 35888
rect 14228 35848 16204 35888
rect 16244 35848 18508 35888
rect 18548 35848 19084 35888
rect 19124 35848 19660 35888
rect 19700 35848 19709 35888
rect 19939 35848 19948 35888
rect 19988 35848 19997 35888
rect 20611 35848 20620 35888
rect 20660 35848 20908 35888
rect 20948 35848 20957 35888
rect 25027 35848 25036 35888
rect 25076 35848 27100 35888
rect 27140 35848 33140 35888
rect 35683 35848 35692 35888
rect 35732 35848 36172 35888
rect 36212 35848 36221 35888
rect 37420 35848 37516 35888
rect 37556 35848 39724 35888
rect 39764 35848 39773 35888
rect 40003 35848 40012 35888
rect 40052 35848 40300 35888
rect 40340 35848 41356 35888
rect 41396 35848 43852 35888
rect 43892 35848 43901 35888
rect 45859 35848 45868 35888
rect 45908 35848 47020 35888
rect 47060 35848 47069 35888
rect 47203 35848 47212 35888
rect 47252 35848 48940 35888
rect 48980 35848 50668 35888
rect 50708 35848 51628 35888
rect 51668 35848 69196 35888
rect 69236 35848 69245 35888
rect 0 35828 80 35848
rect 19267 35804 19325 35805
rect 19948 35804 19988 35848
rect 22627 35804 22685 35805
rect 17539 35764 17548 35804
rect 17588 35764 18892 35804
rect 18932 35764 18941 35804
rect 19267 35764 19276 35804
rect 19316 35764 19988 35804
rect 22542 35764 22636 35804
rect 22676 35764 22685 35804
rect 33100 35804 33140 35848
rect 69187 35847 69245 35848
rect 35491 35804 35549 35805
rect 33100 35764 35500 35804
rect 35540 35764 35549 35804
rect 40195 35764 40204 35804
rect 40244 35764 40396 35804
rect 40436 35764 41260 35804
rect 41300 35764 43276 35804
rect 43316 35764 43325 35804
rect 43651 35764 43660 35804
rect 43700 35764 44140 35804
rect 44180 35764 45580 35804
rect 45620 35764 45629 35804
rect 50947 35764 50956 35804
rect 50996 35764 52012 35804
rect 52052 35764 52061 35804
rect 19267 35763 19325 35764
rect 22627 35763 22685 35764
rect 35491 35763 35549 35764
rect 13795 35680 13804 35720
rect 13844 35680 14092 35720
rect 14132 35680 15340 35720
rect 15380 35680 15389 35720
rect 18787 35680 18796 35720
rect 18836 35680 20044 35720
rect 20084 35680 20093 35720
rect 43939 35680 43948 35720
rect 43988 35680 44716 35720
rect 44756 35680 79180 35720
rect 79220 35680 79229 35720
rect 8131 35596 8140 35636
rect 8180 35596 35404 35636
rect 35444 35596 38380 35636
rect 38420 35596 38429 35636
rect 49315 35596 49324 35636
rect 49364 35596 51916 35636
rect 51956 35596 51965 35636
rect 19267 35552 19325 35553
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19182 35512 19276 35552
rect 19316 35512 19325 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 35788 35512 40588 35552
rect 40628 35512 40637 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 19267 35511 19325 35512
rect 8227 35468 8285 35469
rect 35788 35468 35828 35512
rect 931 35428 940 35468
rect 980 35428 7220 35468
rect 7180 35384 7220 35428
rect 8227 35428 8236 35468
rect 8276 35428 33388 35468
rect 33428 35428 33437 35468
rect 35779 35428 35788 35468
rect 35828 35428 35837 35468
rect 36163 35428 36172 35468
rect 36212 35428 44332 35468
rect 44372 35428 45964 35468
rect 46004 35428 46013 35468
rect 8227 35427 8285 35428
rect 35788 35384 35828 35428
rect 7180 35344 20908 35384
rect 20948 35344 20957 35384
rect 21091 35344 21100 35384
rect 21140 35344 21580 35384
rect 21620 35344 21629 35384
rect 27340 35344 35828 35384
rect 8035 35300 8093 35301
rect 27340 35300 27380 35344
rect 8035 35260 8044 35300
rect 8084 35260 27380 35300
rect 35203 35260 35212 35300
rect 35252 35260 35788 35300
rect 35828 35260 35837 35300
rect 37420 35260 47540 35300
rect 8035 35259 8093 35260
rect 37420 35216 37460 35260
rect 47500 35216 47540 35260
rect 13603 35176 13612 35216
rect 13652 35176 14092 35216
rect 14132 35176 14141 35216
rect 14659 35176 14668 35216
rect 14708 35176 16204 35216
rect 16244 35176 18124 35216
rect 18164 35176 18700 35216
rect 18740 35176 20140 35216
rect 20180 35176 20524 35216
rect 20564 35176 21964 35216
rect 22004 35176 22013 35216
rect 34531 35176 34540 35216
rect 34580 35176 37228 35216
rect 37268 35176 37460 35216
rect 44131 35176 44140 35216
rect 44180 35176 46348 35216
rect 46388 35176 47308 35216
rect 47348 35176 47357 35216
rect 47500 35176 65452 35216
rect 65492 35176 65501 35216
rect 8323 35132 8381 35133
rect 17443 35132 17501 35133
rect 8323 35092 8332 35132
rect 8372 35092 10636 35132
rect 10676 35092 10685 35132
rect 17443 35092 17452 35132
rect 17492 35092 18988 35132
rect 19028 35092 19564 35132
rect 19604 35092 21100 35132
rect 21140 35092 21149 35132
rect 31843 35092 31852 35132
rect 31892 35092 32812 35132
rect 32852 35092 36172 35132
rect 36212 35092 36221 35132
rect 42115 35092 42124 35132
rect 42164 35092 42796 35132
rect 42836 35092 45484 35132
rect 45524 35092 70156 35132
rect 70196 35092 70924 35132
rect 70964 35092 70973 35132
rect 8323 35091 8381 35092
rect 17443 35091 17501 35092
rect 0 34988 80 35068
rect 7843 35048 7901 35049
rect 7843 35008 7852 35048
rect 7892 35008 14476 35048
rect 14516 35008 17260 35048
rect 17300 35008 17309 35048
rect 19075 35008 19084 35048
rect 19124 35008 20140 35048
rect 20180 35008 20189 35048
rect 21379 35008 21388 35048
rect 21428 35008 22732 35048
rect 22772 35008 35116 35048
rect 35156 35008 35165 35048
rect 35395 35008 35404 35048
rect 35444 35008 36364 35048
rect 36404 35008 36413 35048
rect 47299 35008 47308 35048
rect 47348 35008 47540 35048
rect 48163 35008 48172 35048
rect 48212 35008 50764 35048
rect 50804 35008 53356 35048
rect 53396 35008 54028 35048
rect 54068 35008 54077 35048
rect 64387 35008 64396 35048
rect 64436 35008 81484 35048
rect 81524 35008 81533 35048
rect 7843 35007 7901 35008
rect 17251 34964 17309 34965
rect 47500 34964 47540 35008
rect 15331 34924 15340 34964
rect 15380 34924 17260 34964
rect 17300 34924 17309 34964
rect 20035 34924 20044 34964
rect 20084 34924 23116 34964
rect 23156 34924 23788 34964
rect 23828 34924 23837 34964
rect 43075 34924 43084 34964
rect 43124 34924 43468 34964
rect 43508 34924 47212 34964
rect 47252 34924 47261 34964
rect 47500 34924 49900 34964
rect 49940 34924 49949 34964
rect 52003 34924 52012 34964
rect 52052 34924 53836 34964
rect 53876 34924 54508 34964
rect 54548 34924 54557 34964
rect 17251 34923 17309 34924
rect 10627 34840 10636 34880
rect 10676 34840 20332 34880
rect 20372 34840 26284 34880
rect 26324 34840 26333 34880
rect 32515 34840 32524 34880
rect 32564 34840 32908 34880
rect 32948 34840 32957 34880
rect 33100 34840 35692 34880
rect 35732 34840 35741 34880
rect 51907 34840 51916 34880
rect 51956 34840 52972 34880
rect 53012 34840 53021 34880
rect 33100 34796 33140 34840
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 17347 34756 17356 34796
rect 17396 34756 18028 34796
rect 18068 34756 18077 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 18988 34756 33140 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 36355 34756 36364 34796
rect 36404 34756 36940 34796
rect 36980 34756 36989 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 49891 34756 49900 34796
rect 49940 34756 52492 34796
rect 52532 34756 53164 34796
rect 53204 34756 53213 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 7075 34712 7133 34713
rect 18988 34712 19028 34756
rect 7075 34672 7084 34712
rect 7124 34672 19028 34712
rect 26467 34672 26476 34712
rect 26516 34672 26764 34712
rect 26804 34672 30892 34712
rect 30932 34672 32716 34712
rect 32756 34672 36268 34712
rect 36308 34672 36317 34712
rect 47011 34672 47020 34712
rect 47060 34672 48076 34712
rect 48116 34672 49324 34712
rect 49364 34672 49373 34712
rect 7075 34671 7133 34672
rect 16579 34588 16588 34628
rect 16628 34588 19276 34628
rect 19316 34588 19325 34628
rect 21292 34588 25036 34628
rect 25076 34588 25085 34628
rect 27331 34588 27340 34628
rect 27380 34588 28876 34628
rect 28916 34588 31276 34628
rect 31316 34588 33388 34628
rect 33428 34588 33964 34628
rect 34004 34588 34013 34628
rect 4963 34504 4972 34544
rect 5012 34504 7276 34544
rect 7316 34504 7325 34544
rect 7555 34504 7564 34544
rect 7604 34504 12076 34544
rect 12116 34504 12125 34544
rect 12931 34504 12940 34544
rect 12980 34504 13420 34544
rect 13460 34504 13469 34544
rect 21292 34460 21332 34588
rect 35491 34544 35549 34545
rect 62371 34544 62429 34545
rect 35491 34504 35500 34544
rect 35540 34504 35692 34544
rect 35732 34504 38092 34544
rect 38132 34504 38141 34544
rect 42508 34504 49420 34544
rect 49460 34504 49469 34544
rect 49603 34504 49612 34544
rect 49652 34504 62380 34544
rect 62420 34504 62429 34544
rect 35491 34503 35549 34504
rect 17260 34420 19564 34460
rect 19604 34420 21292 34460
rect 21332 34420 21341 34460
rect 22531 34420 22540 34460
rect 22580 34420 25556 34460
rect 17260 34376 17300 34420
rect 25516 34376 25556 34420
rect 42508 34376 42548 34504
rect 62371 34503 62429 34504
rect 62572 34504 68044 34544
rect 68084 34504 68093 34544
rect 62572 34376 62612 34504
rect 5731 34336 5740 34376
rect 5780 34336 7852 34376
rect 7892 34336 17300 34376
rect 22243 34336 22252 34376
rect 22292 34336 24364 34376
rect 24404 34336 24413 34376
rect 25507 34336 25516 34376
rect 25556 34336 27052 34376
rect 27092 34336 29548 34376
rect 29588 34336 29597 34376
rect 30499 34336 30508 34376
rect 30548 34336 31564 34376
rect 31604 34336 32044 34376
rect 32084 34336 32428 34376
rect 32468 34336 32477 34376
rect 34339 34336 34348 34376
rect 34388 34336 42548 34376
rect 45187 34336 45196 34376
rect 45236 34336 62612 34376
rect 62755 34376 62813 34377
rect 62755 34336 62764 34376
rect 62804 34336 64204 34376
rect 64244 34336 64253 34376
rect 64579 34336 64588 34376
rect 64628 34336 66316 34376
rect 66356 34336 68908 34376
rect 68948 34336 70156 34376
rect 70196 34336 70636 34376
rect 70676 34336 70685 34376
rect 22252 34292 22292 34336
rect 62755 34335 62813 34336
rect 20995 34252 21004 34292
rect 21044 34252 22292 34292
rect 27139 34252 27148 34292
rect 27188 34252 29740 34292
rect 29780 34252 30028 34292
rect 30068 34252 30604 34292
rect 30644 34252 30653 34292
rect 77740 34252 82060 34292
rect 82100 34252 82109 34292
rect 0 34148 80 34228
rect 10243 34208 10301 34209
rect 77740 34208 77780 34252
rect 4867 34168 4876 34208
rect 4916 34168 7372 34208
rect 7412 34168 7421 34208
rect 10158 34168 10252 34208
rect 10292 34168 10301 34208
rect 13315 34168 13324 34208
rect 13364 34168 14380 34208
rect 14420 34168 15820 34208
rect 15860 34168 15869 34208
rect 15916 34168 18796 34208
rect 18836 34168 18845 34208
rect 31651 34168 31660 34208
rect 31700 34168 34540 34208
rect 34580 34168 36556 34208
rect 36596 34168 36605 34208
rect 38083 34168 38092 34208
rect 38132 34168 42220 34208
rect 42260 34168 50860 34208
rect 50900 34168 50909 34208
rect 52291 34168 52300 34208
rect 52340 34168 62764 34208
rect 62804 34168 62813 34208
rect 68515 34168 68524 34208
rect 68564 34168 77780 34208
rect 10243 34167 10301 34168
rect 7267 34084 7276 34124
rect 7316 34084 11212 34124
rect 11252 34084 11261 34124
rect 15916 34040 15956 34168
rect 17260 34084 23060 34124
rect 30211 34084 30220 34124
rect 30260 34084 36652 34124
rect 36692 34084 36701 34124
rect 62956 34084 82252 34124
rect 82292 34084 82301 34124
rect 17260 34040 17300 34084
rect 23020 34040 23060 34084
rect 62956 34040 62996 34084
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 5155 34000 5164 34040
rect 5204 34000 9964 34040
rect 10004 34000 10444 34040
rect 10484 34000 10493 34040
rect 13219 34000 13228 34040
rect 13268 34000 13516 34040
rect 13556 34000 15956 34040
rect 16003 34000 16012 34040
rect 16052 34000 17300 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 23020 34000 33196 34040
rect 33236 34000 33245 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 43363 34000 43372 34040
rect 43412 34000 46348 34040
rect 46388 34000 48940 34040
rect 48980 34000 49228 34040
rect 49268 34000 49277 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 50851 34000 50860 34040
rect 50900 34000 52492 34040
rect 52532 34000 61516 34040
rect 61556 34000 61565 34040
rect 62467 34000 62476 34040
rect 62516 34000 62996 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 8323 33916 8332 33956
rect 8372 33916 25228 33956
rect 25268 33916 25277 33956
rect 36931 33916 36940 33956
rect 36980 33916 38764 33956
rect 38804 33916 38813 33956
rect 40291 33916 40300 33956
rect 40340 33916 43988 33956
rect 46915 33916 46924 33956
rect 46964 33916 47636 33956
rect 43948 33872 43988 33916
rect 8227 33832 8236 33872
rect 8276 33832 26188 33872
rect 26228 33832 26237 33872
rect 36643 33832 36652 33872
rect 36692 33832 41164 33872
rect 41204 33832 43276 33872
rect 43316 33832 43325 33872
rect 43948 33832 47540 33872
rect 10339 33748 10348 33788
rect 10388 33748 13228 33788
rect 13268 33748 13277 33788
rect 15811 33748 15820 33788
rect 15860 33748 23980 33788
rect 24020 33748 24029 33788
rect 7939 33664 7948 33704
rect 7988 33664 16012 33704
rect 16052 33664 16061 33704
rect 47500 33536 47540 33832
rect 47596 33620 47636 33916
rect 62476 33872 62516 34000
rect 49411 33832 49420 33872
rect 49460 33832 52300 33872
rect 52340 33832 52349 33872
rect 54019 33832 54028 33872
rect 54068 33832 62516 33872
rect 64579 33832 64588 33872
rect 64628 33832 74188 33872
rect 74228 33832 74237 33872
rect 77740 33832 80908 33872
rect 80948 33832 80957 33872
rect 54691 33788 54749 33789
rect 53155 33748 53164 33788
rect 53204 33748 54700 33788
rect 54740 33748 54749 33788
rect 54691 33747 54749 33748
rect 51331 33664 51340 33704
rect 51380 33664 52780 33704
rect 52820 33664 52829 33704
rect 61507 33664 61516 33704
rect 61556 33664 64396 33704
rect 64436 33664 64445 33704
rect 47596 33580 49132 33620
rect 49172 33580 51052 33620
rect 51092 33580 55180 33620
rect 55220 33580 55229 33620
rect 77740 33536 77780 33832
rect 47500 33496 77780 33536
rect 0 33308 80 33388
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 99811 33200 99869 33201
rect 99920 33200 100000 33220
rect 80803 33160 80812 33200
rect 80852 33160 83116 33200
rect 83156 33160 83165 33200
rect 99811 33160 99820 33200
rect 99860 33160 100000 33200
rect 99811 33159 99869 33160
rect 99920 33140 100000 33160
rect 5539 32948 5597 32949
rect 5454 32908 5548 32948
rect 5588 32908 5597 32948
rect 5539 32907 5597 32908
rect 45571 32656 45580 32696
rect 45620 32656 78508 32696
rect 78548 32656 80140 32696
rect 80180 32656 80189 32696
rect 81187 32656 81196 32696
rect 81236 32656 81868 32696
rect 81908 32656 81917 32696
rect 69091 32612 69149 32613
rect 5251 32572 5260 32612
rect 5300 32572 35212 32612
rect 35252 32572 35261 32612
rect 52003 32572 52012 32612
rect 52052 32572 69100 32612
rect 69140 32572 69149 32612
rect 72643 32572 72652 32612
rect 72692 32572 85421 32612
rect 69091 32571 69149 32572
rect 0 32468 80 32548
rect 8131 32528 8189 32529
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 8131 32488 8140 32528
rect 8180 32488 36460 32528
rect 36500 32488 36509 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 8131 32487 8189 32488
rect 68803 32444 68861 32445
rect 6403 32404 6412 32444
rect 6452 32404 37612 32444
rect 37652 32404 37661 32444
rect 43651 32404 43660 32444
rect 43700 32404 68812 32444
rect 68852 32404 68861 32444
rect 68803 32403 68861 32404
rect 4579 32320 4588 32360
rect 4628 32320 4972 32360
rect 5012 32320 5021 32360
rect 2947 32068 2956 32108
rect 2996 32068 4396 32108
rect 4436 32068 5356 32108
rect 5396 32068 13900 32108
rect 13940 32068 13949 32108
rect 50371 31772 50429 31773
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 50286 31732 50380 31772
rect 50420 31732 50429 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 50371 31731 50429 31732
rect 0 31628 80 31708
rect 7747 31688 7805 31689
rect 7747 31648 7756 31688
rect 7796 31648 17548 31688
rect 17588 31648 18233 31688
rect 18273 31648 18282 31688
rect 79171 31648 79180 31688
rect 79220 31648 81964 31688
rect 82004 31648 82013 31688
rect 7747 31647 7805 31648
rect 10243 31604 10301 31605
rect 5827 31564 5836 31604
rect 5876 31564 10252 31604
rect 10292 31564 15161 31604
rect 15201 31564 15210 31604
rect 10243 31563 10301 31564
rect 5923 31480 5932 31520
rect 5972 31480 16313 31520
rect 16353 31480 16492 31520
rect 16532 31480 16541 31520
rect 80323 31396 80332 31436
rect 80372 31396 81388 31436
rect 81428 31396 81437 31436
rect 97323 31435 97365 31444
rect 97323 31395 97324 31435
rect 97364 31395 97365 31435
rect 97323 31386 97365 31395
rect 3811 31312 3820 31352
rect 3860 31312 4588 31352
rect 4628 31312 4637 31352
rect 81091 31312 81100 31352
rect 81140 31312 81676 31352
rect 81716 31312 81725 31352
rect 80995 31060 81004 31100
rect 81044 31060 83212 31100
rect 83252 31060 85421 31100
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 83107 30892 83116 30932
rect 83156 30892 85421 30932
rect 0 30788 80 30868
rect 83491 30848 83549 30849
rect 80035 30808 80044 30848
rect 80084 30808 80716 30848
rect 80756 30808 82924 30848
rect 82964 30808 83500 30848
rect 83540 30808 83549 30848
rect 83491 30807 83549 30808
rect 4483 30724 4492 30764
rect 4532 30724 5836 30764
rect 5876 30724 5885 30764
rect 4579 30640 4588 30680
rect 4628 30640 5068 30680
rect 5108 30640 5117 30680
rect 78595 30556 78604 30596
rect 78644 30556 79180 30596
rect 79220 30556 79229 30596
rect 3427 30472 3436 30512
rect 3476 30472 4204 30512
rect 4244 30472 4253 30512
rect 81379 30472 81388 30512
rect 81428 30472 82060 30512
rect 82100 30472 82109 30512
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 80035 30220 80044 30260
rect 80084 30220 81772 30260
rect 81812 30220 81821 30260
rect 79651 30136 79660 30176
rect 79700 30136 79948 30176
rect 79988 30136 80620 30176
rect 80660 30136 80669 30176
rect 0 29948 80 30028
rect 81667 29800 81676 29840
rect 81716 29800 83308 29840
rect 83348 29800 83357 29840
rect 80611 29632 80620 29672
rect 80660 29632 81196 29672
rect 81236 29632 81245 29672
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 97323 29397 97365 29406
rect 97323 29357 97324 29397
rect 97364 29357 97365 29397
rect 97323 29348 97365 29357
rect 80803 29212 80812 29252
rect 80852 29212 81388 29252
rect 81428 29212 81437 29252
rect 0 29108 80 29188
rect 5155 29128 5164 29168
rect 5204 29128 5836 29168
rect 5876 29128 5885 29168
rect 4483 29044 4492 29084
rect 4532 29044 4876 29084
rect 4916 29044 4925 29084
rect 3811 28960 3820 29000
rect 3860 28960 5452 29000
rect 5492 28960 5501 29000
rect 78787 28960 78796 29000
rect 78836 28960 79372 29000
rect 79412 28960 79421 29000
rect 3427 28876 3436 28916
rect 3476 28876 4876 28916
rect 4916 28876 4925 28916
rect 79171 28876 79180 28916
rect 79220 28876 81196 28916
rect 81236 28876 81245 28916
rect 84931 28748 84989 28749
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 80323 28708 80332 28748
rect 80372 28708 83212 28748
rect 83252 28708 84940 28748
rect 84980 28708 84989 28748
rect 84931 28707 84989 28708
rect 0 28268 80 28348
rect 7843 28328 7901 28329
rect 4771 28288 4780 28328
rect 4820 28288 7852 28328
rect 7892 28288 7901 28328
rect 80227 28288 80236 28328
rect 80276 28288 81580 28328
rect 81620 28288 81629 28328
rect 7843 28287 7901 28288
rect 4867 28204 4876 28244
rect 4916 28204 5356 28244
rect 5396 28204 5405 28244
rect 83299 28204 83308 28244
rect 83348 28204 85421 28244
rect 4483 28120 4492 28160
rect 4532 28120 4541 28160
rect 4492 28076 4532 28120
rect 4492 28036 4916 28076
rect 4876 27992 4916 28036
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 4867 27952 4876 27992
rect 4916 27952 4925 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 79747 27700 79756 27740
rect 79796 27700 80524 27740
rect 80564 27700 83308 27740
rect 83348 27700 83357 27740
rect 0 27428 80 27508
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 80131 26860 80140 26900
rect 80180 26860 80524 26900
rect 80564 26860 80573 26900
rect 80131 26692 80140 26732
rect 80180 26692 80428 26732
rect 80468 26692 82636 26732
rect 82676 26692 82685 26732
rect 0 26588 80 26668
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 80611 26144 80669 26145
rect 3427 26104 3436 26144
rect 3476 26104 4204 26144
rect 4244 26104 4253 26144
rect 80526 26104 80620 26144
rect 80660 26104 81196 26144
rect 81236 26104 81245 26144
rect 80611 26103 80669 26104
rect 3619 25936 3628 25976
rect 3668 25936 8021 25976
rect 4483 25852 4492 25892
rect 4532 25852 5836 25892
rect 5876 25852 5885 25892
rect 0 25748 80 25828
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 81283 25600 81292 25640
rect 81332 25600 81676 25640
rect 81716 25600 81725 25640
rect 80611 25432 80620 25472
rect 80660 25432 80948 25472
rect 80908 25304 80948 25432
rect 4579 25264 4588 25304
rect 4628 25264 5068 25304
rect 5108 25264 5117 25304
rect 80899 25264 80908 25304
rect 80948 25264 81868 25304
rect 81908 25264 81917 25304
rect 80515 25180 80524 25220
rect 80564 25180 81580 25220
rect 81620 25180 81629 25220
rect 80611 25136 80669 25137
rect 80526 25096 80620 25136
rect 80660 25096 80669 25136
rect 80611 25095 80669 25096
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 0 24908 80 24928
rect 931 24800 989 24801
rect 835 24760 844 24800
rect 884 24760 940 24800
rect 980 24760 989 24800
rect 931 24759 989 24760
rect 81571 24508 81580 24548
rect 81620 24508 82676 24548
rect 82636 24464 82676 24508
rect 82627 24424 82636 24464
rect 82676 24424 92572 24464
rect 92612 24424 92621 24464
rect 82723 24340 82732 24380
rect 82772 24340 90460 24380
rect 90500 24340 90509 24380
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 0 24068 80 24088
rect 835 24044 893 24045
rect 750 24004 844 24044
rect 884 24004 893 24044
rect 5155 24004 5164 24044
rect 5204 24004 5836 24044
rect 5876 24004 5885 24044
rect 81667 24004 81676 24044
rect 81716 24004 83212 24044
rect 83252 24004 87916 24044
rect 87956 24004 87965 24044
rect 835 24003 893 24004
rect 82915 23876 82973 23877
rect 99907 23876 99965 23877
rect 82915 23836 82924 23876
rect 82964 23836 99916 23876
rect 99956 23836 99965 23876
rect 82915 23835 82973 23836
rect 99907 23835 99965 23836
rect 81475 23752 81484 23792
rect 81524 23752 82060 23792
rect 82100 23752 82109 23792
rect 3427 23668 3436 23708
rect 3476 23668 4204 23708
rect 4244 23668 4253 23708
rect 80611 23668 80620 23708
rect 80660 23668 81196 23708
rect 81236 23668 82444 23708
rect 82484 23668 85420 23708
rect 85460 23668 85469 23708
rect 4012 23500 4876 23540
rect 4916 23500 4925 23540
rect 4012 23372 4052 23500
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 3907 23332 3916 23372
rect 3956 23332 4052 23372
rect 4492 23332 5164 23372
rect 5204 23332 5740 23372
rect 5780 23332 5789 23372
rect 0 23288 80 23308
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 0 23228 80 23248
rect 4492 23204 4532 23332
rect 4579 23248 4588 23288
rect 4628 23248 5836 23288
rect 5876 23248 5885 23288
rect 4483 23164 4492 23204
rect 4532 23164 4541 23204
rect 4780 23164 5260 23204
rect 5300 23164 5309 23204
rect 4780 23120 4820 23164
rect 3523 23080 3532 23120
rect 3572 23080 4588 23120
rect 4628 23080 4637 23120
rect 4771 23080 4780 23120
rect 4820 23080 4829 23120
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 0 22448 80 22468
rect 0 22408 652 22448
rect 692 22408 701 22448
rect 3331 22408 3340 22448
rect 3380 22408 3628 22448
rect 3668 22408 3677 22448
rect 0 22388 80 22408
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 5059 21904 5068 21944
rect 5108 21904 8021 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 3331 21652 3340 21692
rect 3380 21652 5356 21692
rect 5396 21652 5405 21692
rect 0 21608 80 21628
rect 6403 21608 6461 21609
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 3427 21568 3436 21608
rect 3476 21568 6412 21608
rect 6452 21568 6461 21608
rect 0 21548 80 21568
rect 6403 21567 6461 21568
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 81475 20980 81484 21020
rect 81524 20980 84460 21020
rect 84500 20980 84509 21020
rect 5731 20896 5740 20936
rect 5780 20896 8021 20936
rect 82051 20812 82060 20852
rect 82100 20812 82140 20852
rect 0 20768 80 20788
rect 82060 20768 82100 20812
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 4195 20728 4204 20768
rect 4244 20728 4972 20768
rect 5012 20728 5021 20768
rect 79459 20728 79468 20768
rect 79508 20728 83308 20768
rect 83348 20728 83357 20768
rect 0 20708 80 20728
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 82723 20056 82732 20096
rect 82772 20056 96748 20096
rect 96788 20056 96797 20096
rect 3907 19972 3916 20012
rect 3956 19972 5068 20012
rect 5108 19972 5836 20012
rect 5876 19972 5885 20012
rect 0 19928 80 19948
rect 99920 19928 100000 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 4003 19888 4012 19928
rect 4052 19888 4300 19928
rect 4340 19888 4349 19928
rect 98563 19888 98572 19928
rect 98612 19888 100000 19928
rect 0 19868 80 19888
rect 99920 19868 100000 19888
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 2947 19048 2956 19088
rect 2996 19048 4012 19088
rect 4052 19048 5836 19088
rect 5876 19048 8021 19088
rect 0 19028 80 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 5923 18880 5932 18920
rect 5972 18880 8021 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 2275 18628 2284 18668
rect 2324 18628 3244 18668
rect 3284 18628 4972 18668
rect 5012 18628 5021 18668
rect 2179 18544 2188 18584
rect 2228 18544 2572 18584
rect 2612 18544 2621 18584
rect 3907 18544 3916 18584
rect 3956 18544 4204 18584
rect 4244 18544 4684 18584
rect 4724 18544 4733 18584
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 75811 17956 75820 17996
rect 75860 17956 98860 17996
rect 98900 17956 98909 17996
rect 2563 17872 2572 17912
rect 2612 17872 2860 17912
rect 2900 17872 5068 17912
rect 5108 17872 8021 17912
rect 2467 17788 2476 17828
rect 2516 17788 3820 17828
rect 3860 17788 3869 17828
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 0 17348 80 17368
rect 2083 17284 2092 17324
rect 2132 17284 3916 17324
rect 3956 17300 4724 17324
rect 3956 17284 4659 17300
rect 4584 17260 4659 17284
rect 4699 17260 4724 17300
rect 1315 17200 1324 17240
rect 1364 17200 2284 17240
rect 2324 17200 3052 17240
rect 3092 17200 3101 17240
rect 3907 16864 3916 16904
rect 3956 16864 8021 16904
rect 78403 16780 78412 16820
rect 78452 16780 80620 16820
rect 80660 16780 81388 16820
rect 81428 16780 81437 16820
rect 7843 16763 7901 16764
rect 7660 16736 7852 16763
rect 5827 16696 5836 16736
rect 5876 16723 7852 16736
rect 7892 16723 8040 16763
rect 5876 16696 7700 16723
rect 7843 16722 7901 16723
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 5923 16528 5932 16568
rect 5972 16528 8021 16568
rect 0 16508 80 16528
rect 1795 16444 1804 16484
rect 1844 16444 2572 16484
rect 2612 16444 3244 16484
rect 3284 16444 3916 16484
rect 3956 16444 3965 16484
rect 76963 16232 77021 16233
rect 76963 16192 76972 16232
rect 77012 16192 78508 16232
rect 78548 16192 78557 16232
rect 76963 16191 77021 16192
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 0 15728 80 15748
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 0 15668 80 15688
rect 4483 15604 4492 15644
rect 4532 15604 5836 15644
rect 5876 15604 5885 15644
rect 4579 15520 4588 15560
rect 4628 15520 5932 15560
rect 5972 15520 5981 15560
rect 1219 15476 1277 15477
rect 1134 15436 1228 15476
rect 1268 15436 1277 15476
rect 3427 15436 3436 15476
rect 3476 15436 4204 15476
rect 4244 15436 4253 15476
rect 1219 15435 1277 15436
rect 835 15352 844 15392
rect 884 15352 1516 15392
rect 1556 15352 1565 15392
rect 2947 15352 2956 15392
rect 2996 15352 4108 15392
rect 4148 15352 4157 15392
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 0 14888 80 14908
rect 0 14848 1036 14888
rect 1076 14848 1085 14888
rect 1603 14848 1612 14888
rect 1652 14848 1900 14888
rect 1940 14848 3244 14888
rect 3284 14848 8021 14888
rect 0 14828 80 14848
rect 2083 14680 2092 14720
rect 2132 14680 4684 14720
rect 4724 14680 4876 14720
rect 4916 14680 6412 14720
rect 6452 14680 6461 14720
rect 3811 14512 3820 14552
rect 3860 14512 4588 14552
rect 4628 14512 4637 14552
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 4195 14176 4204 14216
rect 4244 14176 5068 14216
rect 5108 14176 5117 14216
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 0 13988 80 14008
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 1219 13168 1228 13208
rect 1268 13168 1420 13208
rect 1460 13168 3724 13208
rect 3764 13168 3773 13208
rect 4675 13168 4684 13208
rect 4724 13168 4876 13208
rect 4916 13168 4925 13208
rect 0 13148 80 13168
rect 1987 13000 1996 13040
rect 2036 13000 2572 13040
rect 2612 13000 4204 13040
rect 4244 13000 4253 13040
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 7660 12821 8040 12861
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 7660 12788 7700 12821
rect 2755 12748 2764 12788
rect 2804 12748 5740 12788
rect 5780 12748 7700 12788
rect 3907 12664 3916 12704
rect 3956 12664 5836 12704
rect 5876 12664 8021 12704
rect 835 12580 844 12620
rect 884 12580 1420 12620
rect 1460 12580 1469 12620
rect 1795 12496 1804 12536
rect 1844 12496 2476 12536
rect 2516 12496 4972 12536
rect 5012 12496 8021 12536
rect 0 12368 80 12388
rect 0 12328 1036 12368
rect 1076 12328 1085 12368
rect 2947 12328 2956 12368
rect 2996 12328 3916 12368
rect 3956 12328 5836 12368
rect 5876 12328 8021 12368
rect 0 12308 80 12328
rect 1699 12244 1708 12284
rect 1748 12244 3244 12284
rect 3284 12244 7700 12284
rect 7660 12242 7700 12244
rect 7660 12202 8040 12242
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 5251 11992 5260 12032
rect 5300 11992 8021 12032
rect 4291 11656 4300 11696
rect 4340 11656 5260 11696
rect 5300 11656 5309 11696
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 3715 11488 3724 11528
rect 3764 11488 4684 11528
rect 4724 11488 4876 11528
rect 4916 11488 4925 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 835 10900 844 10940
rect 884 10900 1804 10940
rect 1844 10900 1853 10940
rect 643 10732 652 10772
rect 692 10732 701 10772
rect 0 10688 80 10708
rect 652 10688 692 10732
rect 0 10648 692 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 835 10228 844 10268
rect 884 10228 1900 10268
rect 1940 10228 1949 10268
rect 2659 10144 2668 10184
rect 2708 10144 2900 10184
rect 2947 10144 2956 10184
rect 2996 10144 4588 10184
rect 4628 10144 4972 10184
rect 5012 10144 5164 10184
rect 5204 10144 5213 10184
rect 2860 10100 2900 10144
rect 2860 10060 4204 10100
rect 4244 10060 5836 10100
rect 5876 10060 5885 10100
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 0 9788 80 9808
rect 835 9428 893 9429
rect 750 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 98760 9379 98860 9419
rect 98900 9379 98909 9419
rect 81379 9220 81388 9260
rect 81428 9251 82484 9260
rect 81428 9220 82840 9251
rect 82444 9211 82840 9220
rect 98731 9213 98789 9214
rect 98731 9173 98740 9213
rect 98780 9173 98789 9213
rect 98731 9172 98789 9173
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 82819 9083 82877 9084
rect 82819 9043 82828 9083
rect 82868 9043 82877 9083
rect 82819 9042 82877 9043
rect 98731 9045 98789 9046
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 98731 9005 98740 9045
rect 98780 9005 98789 9045
rect 98731 9004 98789 9005
rect 0 8948 80 8968
rect 98851 8877 98909 8878
rect 98760 8837 98860 8877
rect 98900 8837 98909 8877
rect 98851 8836 98909 8837
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 0 8168 80 8188
rect 0 8128 556 8168
rect 596 8128 605 8168
rect 4579 8128 4588 8168
rect 4628 8128 5740 8168
rect 5780 8128 5789 8168
rect 0 8108 80 8128
rect 3427 7960 3436 8000
rect 3476 7960 4300 8000
rect 4340 7960 4349 8000
rect 4675 7960 4684 8000
rect 4724 7960 5164 8000
rect 5204 7960 5213 8000
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 0 7328 80 7348
rect 40867 7328 40925 7329
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 40867 7288 40876 7328
rect 40929 7288 41011 7328
rect 0 7268 80 7288
rect 40867 7287 40925 7288
rect 26323 7204 26332 7244
rect 26372 7204 26420 7244
rect 26380 7160 26420 7204
rect 2179 7120 2188 7160
rect 2228 7120 25612 7160
rect 25652 7120 25661 7160
rect 26380 7120 71404 7160
rect 71444 7120 71453 7160
rect 7939 7036 7948 7076
rect 7988 7036 33772 7076
rect 33812 7036 33821 7076
rect 37507 7036 37516 7076
rect 37556 7036 37900 7076
rect 37940 7036 82732 7076
rect 82772 7036 82781 7076
rect 5923 6952 5932 6992
rect 5972 6952 23788 6992
rect 23828 6952 23837 6992
rect 7747 6824 7805 6825
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 7747 6784 7756 6824
rect 7796 6784 17452 6824
rect 17492 6784 17501 6824
rect 33379 6784 33388 6824
rect 33428 6784 37612 6824
rect 37652 6784 37661 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 7747 6783 7805 6784
rect 1795 6700 1804 6740
rect 1844 6700 49036 6740
rect 49076 6700 49085 6740
rect 72739 6656 72797 6657
rect 82339 6656 82397 6657
rect 1891 6616 1900 6656
rect 1940 6616 37460 6656
rect 37603 6616 37612 6656
rect 37652 6616 72748 6656
rect 72788 6616 72797 6656
rect 80515 6616 80524 6656
rect 80564 6616 82348 6656
rect 82388 6616 82397 6656
rect 8131 6572 8189 6573
rect 8131 6532 8140 6572
rect 8180 6532 36172 6572
rect 36212 6532 36221 6572
rect 8131 6531 8189 6532
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 1411 6448 1420 6488
rect 1460 6448 31756 6488
rect 31796 6448 31805 6488
rect 0 6428 80 6448
rect 37420 6236 37460 6616
rect 72739 6615 72797 6616
rect 82339 6615 82397 6616
rect 98947 6656 99005 6657
rect 99920 6656 100000 6676
rect 98947 6616 98956 6656
rect 98996 6616 100000 6656
rect 98947 6615 99005 6616
rect 99920 6596 100000 6616
rect 68803 6488 68861 6489
rect 44515 6448 44524 6488
rect 44564 6448 68812 6488
rect 68852 6448 68861 6488
rect 68803 6447 68861 6448
rect 77740 6448 78508 6488
rect 78548 6448 78557 6488
rect 77740 6320 77780 6448
rect 40771 6280 40780 6320
rect 40820 6280 41068 6320
rect 41108 6280 77780 6320
rect 37420 6196 49612 6236
rect 49652 6196 49661 6236
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 35395 5816 35453 5817
rect 35310 5776 35404 5816
rect 35444 5776 35453 5816
rect 35395 5775 35453 5776
rect 29251 5692 29260 5732
rect 29300 5692 34924 5732
rect 34964 5692 34973 5732
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 18691 5608 18700 5648
rect 18740 5608 21580 5648
rect 21620 5608 23980 5648
rect 24020 5608 24029 5648
rect 34627 5608 34636 5648
rect 34676 5608 35020 5648
rect 35060 5608 35069 5648
rect 0 5588 80 5608
rect 1123 5524 1132 5564
rect 1172 5524 35116 5564
rect 35156 5524 35165 5564
rect 931 5440 940 5480
rect 980 5440 35404 5480
rect 35444 5440 35453 5480
rect 40579 5440 40588 5480
rect 40628 5440 72652 5480
rect 72692 5440 72701 5480
rect 4771 5356 4780 5396
rect 4820 5356 18700 5396
rect 18740 5356 18749 5396
rect 23212 5356 26284 5396
rect 26324 5356 26333 5396
rect 32707 5356 32716 5396
rect 32756 5356 49420 5396
rect 49460 5356 49469 5396
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 5059 5272 5068 5312
rect 5108 5272 17932 5312
rect 17972 5272 17981 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 8515 5228 8573 5229
rect 23212 5228 23252 5356
rect 35203 5312 35261 5313
rect 23683 5272 23692 5312
rect 23732 5272 24652 5312
rect 24692 5272 24701 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 35118 5272 35212 5312
rect 35252 5272 35261 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 35203 5271 35261 5272
rect 35011 5228 35069 5229
rect 69187 5228 69245 5229
rect 8515 5188 8524 5228
rect 8564 5188 23252 5228
rect 23299 5188 23308 5228
rect 23348 5188 24748 5228
rect 24788 5188 24797 5228
rect 35011 5188 35020 5228
rect 35060 5188 35788 5228
rect 35828 5188 35837 5228
rect 52195 5188 52204 5228
rect 52244 5188 69196 5228
rect 69236 5188 69245 5228
rect 8515 5187 8573 5188
rect 35011 5187 35069 5188
rect 69187 5187 69245 5188
rect 7075 5144 7133 5145
rect 39427 5144 39485 5145
rect 71491 5144 71549 5145
rect 7075 5104 7084 5144
rect 7124 5104 35980 5144
rect 36020 5104 36029 5144
rect 39342 5104 39436 5144
rect 39476 5104 39485 5144
rect 49987 5104 49996 5144
rect 50036 5104 71500 5144
rect 71540 5104 71549 5144
rect 7075 5103 7133 5104
rect 39427 5103 39485 5104
rect 71491 5103 71549 5104
rect 46339 5020 46348 5060
rect 46388 5020 47596 5060
rect 47636 5020 48364 5060
rect 48404 5020 48413 5060
rect 53923 5020 53932 5060
rect 53972 5020 79468 5060
rect 79508 5020 79517 5060
rect 73507 4976 73565 4977
rect 7075 4936 7084 4976
rect 7124 4936 42892 4976
rect 42932 4936 42941 4976
rect 43843 4936 43852 4976
rect 43892 4936 46732 4976
rect 46772 4936 47980 4976
rect 48020 4936 48029 4976
rect 49507 4936 49516 4976
rect 49556 4936 73516 4976
rect 73556 4936 73565 4976
rect 73507 4935 73565 4936
rect 45187 4852 45196 4892
rect 45236 4852 47540 4892
rect 48067 4852 48076 4892
rect 48116 4852 52588 4892
rect 52628 4852 55084 4892
rect 55124 4852 55133 4892
rect 0 4808 80 4828
rect 35011 4808 35069 4809
rect 47500 4808 47540 4852
rect 53731 4808 53789 4809
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 1027 4768 1036 4808
rect 1076 4768 32716 4808
rect 32756 4768 32765 4808
rect 32899 4768 32908 4808
rect 32948 4768 33292 4808
rect 33332 4768 33341 4808
rect 33475 4768 33484 4808
rect 33524 4768 34444 4808
rect 34484 4768 34493 4808
rect 34926 4768 35020 4808
rect 35060 4768 35069 4808
rect 35491 4768 35500 4808
rect 35540 4768 36940 4808
rect 36980 4768 36989 4808
rect 37420 4768 37804 4808
rect 37844 4768 37853 4808
rect 39235 4768 39244 4808
rect 39284 4768 40684 4808
rect 40724 4768 40733 4808
rect 47500 4768 50380 4808
rect 50420 4768 53740 4808
rect 53780 4768 53789 4808
rect 0 4748 80 4768
rect 33484 4724 33524 4768
rect 35011 4767 35069 4768
rect 37420 4724 37460 4768
rect 53731 4767 53789 4768
rect 49699 4724 49757 4725
rect 18307 4684 18316 4724
rect 18356 4684 21100 4724
rect 21140 4684 21149 4724
rect 24355 4684 24364 4724
rect 24404 4684 24748 4724
rect 24788 4684 24797 4724
rect 32035 4684 32044 4724
rect 32084 4684 32428 4724
rect 32468 4684 33524 4724
rect 35203 4684 35212 4724
rect 35252 4684 37460 4724
rect 41923 4684 41932 4724
rect 41972 4684 42220 4724
rect 42260 4684 43852 4724
rect 43892 4684 43901 4724
rect 49614 4684 49708 4724
rect 49748 4684 49757 4724
rect 49699 4683 49757 4684
rect 22627 4600 22636 4640
rect 22676 4600 22924 4640
rect 22964 4600 25036 4640
rect 25076 4600 25085 4640
rect 26275 4600 26284 4640
rect 26324 4600 40876 4640
rect 40916 4600 40925 4640
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 24835 4516 24844 4556
rect 24884 4516 25708 4556
rect 25748 4516 25757 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 34627 4432 34636 4472
rect 34676 4432 35596 4472
rect 35636 4432 35645 4472
rect 42403 4432 42412 4472
rect 42452 4432 46828 4472
rect 46868 4432 52204 4472
rect 52244 4432 52253 4472
rect 31651 4348 31660 4388
rect 31700 4348 32140 4388
rect 32180 4348 32189 4388
rect 34435 4348 34444 4388
rect 34484 4348 36076 4388
rect 36116 4348 36125 4388
rect 47107 4348 47116 4388
rect 47156 4348 48076 4388
rect 48116 4348 48125 4388
rect 8131 4264 8140 4304
rect 8180 4264 34924 4304
rect 34964 4264 35596 4304
rect 35636 4264 36172 4304
rect 36212 4264 36221 4304
rect 49219 4264 49228 4304
rect 49268 4264 49900 4304
rect 49940 4264 49949 4304
rect 8323 4220 8381 4221
rect 8323 4180 8332 4220
rect 8372 4180 18508 4220
rect 18548 4180 18557 4220
rect 18691 4180 18700 4220
rect 18740 4180 19276 4220
rect 19316 4180 19325 4220
rect 20899 4180 20908 4220
rect 20948 4180 22444 4220
rect 22484 4180 22493 4220
rect 24643 4180 24652 4220
rect 24692 4180 27148 4220
rect 27188 4180 27436 4220
rect 27476 4180 27485 4220
rect 34531 4180 34540 4220
rect 34580 4180 37036 4220
rect 37076 4180 37085 4220
rect 40483 4180 40492 4220
rect 40532 4180 42316 4220
rect 42356 4180 44140 4220
rect 44180 4180 45196 4220
rect 45236 4180 45245 4220
rect 45379 4180 45388 4220
rect 45428 4180 46348 4220
rect 46388 4180 46732 4220
rect 46772 4180 46781 4220
rect 8323 4179 8381 4180
rect 32611 4136 32669 4137
rect 35203 4136 35261 4137
rect 35395 4136 35453 4137
rect 36739 4136 36797 4137
rect 5155 4096 5164 4136
rect 5204 4096 18124 4136
rect 18164 4096 20428 4136
rect 20468 4096 21772 4136
rect 21812 4096 22540 4136
rect 22580 4096 22589 4136
rect 25123 4096 25132 4136
rect 25172 4096 25612 4136
rect 25652 4096 27724 4136
rect 27764 4096 27773 4136
rect 32526 4096 32620 4136
rect 32660 4096 32669 4136
rect 33091 4096 33100 4136
rect 33140 4096 34828 4136
rect 34868 4096 34877 4136
rect 35107 4096 35116 4136
rect 35156 4096 35212 4136
rect 35252 4096 35261 4136
rect 35310 4096 35404 4136
rect 35444 4096 35453 4136
rect 36654 4096 36748 4136
rect 36788 4096 36797 4136
rect 32611 4095 32669 4096
rect 35203 4095 35261 4096
rect 35395 4095 35453 4096
rect 36739 4095 36797 4096
rect 37507 4136 37565 4137
rect 69091 4136 69149 4137
rect 37507 4096 37516 4136
rect 37556 4096 38860 4136
rect 38900 4096 41164 4136
rect 41204 4096 41213 4136
rect 41731 4096 41740 4136
rect 41780 4096 44044 4136
rect 44084 4096 49612 4136
rect 49652 4096 49804 4136
rect 49844 4096 52396 4136
rect 52436 4096 69100 4136
rect 69140 4096 69149 4136
rect 37507 4095 37565 4096
rect 69091 4095 69149 4096
rect 17260 4012 17356 4052
rect 17396 4012 19564 4052
rect 19604 4012 20716 4052
rect 20756 4012 21676 4052
rect 21716 4012 21725 4052
rect 29923 4012 29932 4052
rect 29972 4012 36076 4052
rect 36116 4012 36125 4052
rect 36835 4012 36844 4052
rect 36884 4012 37612 4052
rect 37652 4012 37661 4052
rect 40003 4012 40012 4052
rect 40052 4012 42220 4052
rect 42260 4012 42892 4052
rect 42932 4012 42941 4052
rect 46723 4012 46732 4052
rect 46772 4012 48940 4052
rect 48980 4012 50188 4052
rect 50228 4012 51532 4052
rect 51572 4012 53068 4052
rect 53108 4012 53117 4052
rect 0 3968 80 3988
rect 17260 3968 17300 4012
rect 36844 3968 36884 4012
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 17251 3928 17260 3968
rect 17300 3928 17309 3968
rect 18499 3928 18508 3968
rect 18548 3928 20908 3968
rect 20948 3928 20957 3968
rect 21571 3928 21580 3968
rect 21620 3928 23212 3968
rect 23252 3928 23692 3968
rect 23732 3928 23741 3968
rect 31747 3928 31756 3968
rect 31796 3928 33196 3968
rect 33236 3928 36884 3968
rect 37699 3928 37708 3968
rect 37748 3928 39148 3968
rect 39188 3928 39628 3968
rect 39668 3928 39677 3968
rect 40867 3928 40876 3968
rect 40916 3928 43180 3968
rect 43220 3928 43229 3968
rect 0 3908 80 3928
rect 8035 3884 8093 3885
rect 8035 3844 8044 3884
rect 8084 3844 27380 3884
rect 29731 3844 29740 3884
rect 29780 3844 39532 3884
rect 39572 3844 39581 3884
rect 8035 3843 8093 3844
rect 27340 3800 27380 3844
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 27340 3760 34484 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 37123 3760 37132 3800
rect 37172 3760 37996 3800
rect 38036 3760 39052 3800
rect 39092 3760 49228 3800
rect 49268 3760 49277 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 34444 3716 34484 3760
rect 4099 3676 4108 3716
rect 4148 3676 17356 3716
rect 17396 3676 17405 3716
rect 22435 3676 22444 3716
rect 22484 3676 32236 3716
rect 32276 3676 32285 3716
rect 34444 3676 35788 3716
rect 35828 3676 40108 3716
rect 40148 3676 40157 3716
rect 46915 3676 46924 3716
rect 46964 3676 50860 3716
rect 50900 3676 52492 3716
rect 52532 3676 53548 3716
rect 53588 3676 53597 3716
rect 32707 3592 32716 3632
rect 32756 3592 33100 3632
rect 33140 3592 33149 3632
rect 34051 3592 34060 3632
rect 34100 3592 35692 3632
rect 35732 3592 35884 3632
rect 35924 3592 35933 3632
rect 49315 3592 49324 3632
rect 49364 3592 80716 3632
rect 80756 3592 80765 3632
rect 23683 3508 23692 3548
rect 23732 3508 25516 3548
rect 25556 3508 25565 3548
rect 27235 3508 27244 3548
rect 27284 3508 29740 3548
rect 29780 3508 29789 3548
rect 33859 3508 33868 3548
rect 33908 3508 34348 3548
rect 34388 3508 35788 3548
rect 35828 3508 35837 3548
rect 40963 3508 40972 3548
rect 41012 3508 44236 3548
rect 44276 3508 44716 3548
rect 44756 3508 44765 3548
rect 47299 3508 47308 3548
rect 47348 3508 47540 3548
rect 49219 3508 49228 3548
rect 49268 3508 49708 3548
rect 49748 3508 49757 3548
rect 49891 3508 49900 3548
rect 49940 3508 80908 3548
rect 80948 3508 80957 3548
rect 47500 3464 47540 3508
rect 8227 3424 8236 3464
rect 8276 3424 24556 3464
rect 24596 3424 28588 3464
rect 28628 3424 28637 3464
rect 32131 3424 32140 3464
rect 32180 3424 39148 3464
rect 39188 3424 39197 3464
rect 39523 3424 39532 3464
rect 39572 3424 39916 3464
rect 39956 3424 43084 3464
rect 43124 3424 43133 3464
rect 44515 3424 44524 3464
rect 44564 3424 47116 3464
rect 47156 3424 47165 3464
rect 47500 3424 48364 3464
rect 48404 3424 50764 3464
rect 50804 3424 50813 3464
rect 739 3340 748 3380
rect 788 3340 32620 3380
rect 32660 3340 37708 3380
rect 37748 3340 37757 3380
rect 47779 3340 47788 3380
rect 47828 3340 50476 3380
rect 50516 3340 50525 3380
rect 21283 3256 21292 3296
rect 21332 3256 21868 3296
rect 21908 3256 21917 3296
rect 8227 3212 8285 3213
rect 8227 3172 8236 3212
rect 8276 3172 30412 3212
rect 30452 3172 31180 3212
rect 31220 3172 31229 3212
rect 8227 3171 8285 3172
rect 0 3128 80 3148
rect 0 3088 652 3128
rect 692 3088 701 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 35683 3004 35692 3044
rect 35732 3004 39052 3044
rect 39092 3004 46444 3044
rect 46484 3004 46493 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 27235 2920 27244 2960
rect 27284 2920 27724 2960
rect 27764 2920 28780 2960
rect 28820 2920 32620 2960
rect 32660 2920 32669 2960
rect 46147 2920 46156 2960
rect 46196 2920 46732 2960
rect 46772 2920 47116 2960
rect 47156 2920 47165 2960
rect 8323 2836 8332 2876
rect 8372 2836 25996 2876
rect 26036 2836 28108 2876
rect 28148 2836 28157 2876
rect 20611 2752 20620 2792
rect 20660 2752 21484 2792
rect 21524 2752 22732 2792
rect 22772 2752 22781 2792
rect 20515 2668 20524 2708
rect 20564 2668 23500 2708
rect 23540 2668 24268 2708
rect 24308 2668 24317 2708
rect 39427 2668 39436 2708
rect 39476 2668 43852 2708
rect 43892 2668 44908 2708
rect 44948 2668 45100 2708
rect 45140 2668 45149 2708
rect 27139 2584 27148 2624
rect 27188 2584 27628 2624
rect 27668 2584 28012 2624
rect 28052 2584 30700 2624
rect 30740 2584 33196 2624
rect 33236 2584 33245 2624
rect 33475 2584 33484 2624
rect 33524 2584 34828 2624
rect 34868 2584 36076 2624
rect 36116 2584 36125 2624
rect 37891 2584 37900 2624
rect 37940 2584 38860 2624
rect 38900 2584 38909 2624
rect 39715 2584 39724 2624
rect 39764 2584 40108 2624
rect 40148 2584 41356 2624
rect 41396 2584 41405 2624
rect 47395 2584 47404 2624
rect 47444 2584 48172 2624
rect 48212 2584 48364 2624
rect 48404 2584 48413 2624
rect 38179 2500 38188 2540
rect 38228 2500 39628 2540
rect 39668 2500 39820 2540
rect 39860 2500 40972 2540
rect 41012 2500 41021 2540
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 0 2228 80 2248
rect 66211 2204 66269 2205
rect 46243 2164 46252 2204
rect 46292 2164 47212 2204
rect 47252 2164 48940 2204
rect 48980 2164 66220 2204
rect 66260 2164 66269 2204
rect 66211 2163 66269 2164
rect 30307 2080 30316 2120
rect 30356 2080 32044 2120
rect 32084 2080 32524 2120
rect 32564 2080 32573 2120
rect 34627 2080 34636 2120
rect 34676 2080 35404 2120
rect 35444 2080 35453 2120
rect 41347 2080 41356 2120
rect 41396 2080 44236 2120
rect 44276 2080 44285 2120
rect 24643 1996 24652 2036
rect 24692 1996 25036 2036
rect 25076 1996 27148 2036
rect 27188 1996 27197 2036
rect 28099 1996 28108 2036
rect 28148 1996 29740 2036
rect 29780 1996 30892 2036
rect 30932 1996 37900 2036
rect 37940 1996 37949 2036
rect 41260 1996 43948 2036
rect 43988 1996 44140 2036
rect 44180 1996 44189 2036
rect 45187 1996 45196 2036
rect 45236 1996 47500 2036
rect 47540 1996 47549 2036
rect 48451 1996 48460 2036
rect 48500 1996 50860 2036
rect 50900 1996 50909 2036
rect 41260 1952 41300 1996
rect 24355 1912 24364 1952
rect 24404 1912 26956 1952
rect 26996 1912 27005 1952
rect 28579 1912 28588 1952
rect 28628 1912 33484 1952
rect 33524 1912 33533 1952
rect 36931 1912 36940 1952
rect 36980 1912 37020 1952
rect 40579 1912 40588 1952
rect 40628 1912 41260 1952
rect 41300 1912 41309 1952
rect 43075 1912 43084 1952
rect 43124 1912 45292 1952
rect 45332 1912 45868 1952
rect 45908 1912 46252 1952
rect 46292 1912 46301 1952
rect 36940 1868 36980 1912
rect 26083 1828 26092 1868
rect 26132 1828 30028 1868
rect 30068 1828 33964 1868
rect 34004 1828 39724 1868
rect 39764 1828 42220 1868
rect 42260 1828 42269 1868
rect 80899 1828 80908 1868
rect 80948 1828 91316 1868
rect 23971 1744 23980 1784
rect 24020 1744 25900 1784
rect 25940 1744 25949 1784
rect 27340 1744 29260 1784
rect 29300 1744 29309 1784
rect 35203 1744 35212 1784
rect 35252 1744 37748 1784
rect 27340 1700 27380 1744
rect 37708 1700 37748 1744
rect 26947 1660 26956 1700
rect 26996 1660 27380 1700
rect 28291 1660 28300 1700
rect 28340 1660 32332 1700
rect 32372 1660 34636 1700
rect 34676 1660 34685 1700
rect 37699 1660 37708 1700
rect 37748 1660 38572 1700
rect 38612 1660 38621 1700
rect 39235 1576 39244 1616
rect 39284 1576 90740 1616
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 80707 1492 80716 1532
rect 80756 1492 89972 1532
rect 89932 1448 89972 1492
rect 90700 1479 90740 1576
rect 91075 1479 91133 1480
rect 91276 1479 91316 1828
rect 90124 1448 90537 1460
rect 36739 1408 36748 1448
rect 36788 1408 44812 1448
rect 44852 1408 47308 1448
rect 47348 1408 47788 1448
rect 47828 1408 47837 1448
rect 89932 1420 90537 1448
rect 90577 1420 90586 1460
rect 90700 1439 90929 1479
rect 90969 1439 90978 1479
rect 91075 1439 91084 1479
rect 91161 1439 91219 1479
rect 91276 1439 91313 1479
rect 91353 1439 91362 1479
rect 91075 1438 91133 1439
rect 89932 1408 90164 1420
rect 28387 1324 28396 1364
rect 28436 1324 30796 1364
rect 30836 1324 35116 1364
rect 35156 1324 35165 1364
rect 35587 1324 35596 1364
rect 35636 1324 37324 1364
rect 37364 1324 37373 1364
rect 38851 1324 38860 1364
rect 38900 1324 40108 1364
rect 40148 1324 40157 1364
rect 40675 1156 40684 1196
rect 40724 1156 90729 1196
rect 90769 1156 90778 1196
rect 32419 1072 32428 1112
rect 32468 1072 35020 1112
rect 35060 1072 35308 1112
rect 35348 1072 35357 1112
rect 38467 1072 38476 1112
rect 38516 1072 40204 1112
rect 40244 1072 40253 1112
rect 40483 1072 40492 1112
rect 40532 1072 42604 1112
rect 42644 1072 42653 1112
rect 44323 1072 44332 1112
rect 44372 1072 46540 1112
rect 46580 1072 46589 1112
rect 47587 1072 47596 1112
rect 47636 1072 50188 1112
rect 50228 1072 50237 1112
rect 32515 988 32524 1028
rect 32564 988 32716 1028
rect 32756 988 34924 1028
rect 34964 988 35500 1028
rect 35540 988 38188 1028
rect 38228 988 38237 1028
rect 27043 904 27052 944
rect 27092 904 28300 944
rect 28340 904 28349 944
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 5548 37948 5588 37988
rect 8524 37948 8564 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 44524 35932 44564 35972
rect 69196 35848 69236 35888
rect 19276 35764 19316 35804
rect 22636 35764 22676 35804
rect 35500 35764 35540 35804
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19276 35512 19316 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 8236 35428 8276 35468
rect 8044 35260 8084 35300
rect 8332 35092 8372 35132
rect 17452 35092 17492 35132
rect 7852 35008 7892 35048
rect 17260 34924 17300 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 7084 34672 7124 34712
rect 35500 34504 35540 34544
rect 62380 34504 62420 34544
rect 62764 34336 62804 34376
rect 10252 34168 10292 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 54700 33748 54740 33788
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 99820 33160 99860 33200
rect 5548 32908 5588 32948
rect 69100 32572 69140 32612
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8140 32488 8180 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 68812 32404 68852 32444
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 50380 31732 50420 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 7756 31648 7796 31688
rect 10252 31564 10292 31604
rect 97324 31395 97364 31435
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 83500 30808 83540 30848
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 97324 29357 97364 29397
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 84940 28708 84980 28748
rect 7852 28288 7892 28328
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 80620 26104 80660 26144
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 80620 25096 80660 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 940 24760 980 24800
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 844 24004 884 24044
rect 82924 23836 82964 23876
rect 99916 23836 99956 23876
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 6412 21568 6452 21608
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 7852 16723 7892 16763
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 76972 16192 77012 16232
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 1228 15436 1268 15476
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 844 9388 884 9428
rect 98740 9173 98780 9213
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 82828 9043 82868 9083
rect 98740 9005 98780 9045
rect 98860 8837 98900 8877
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 40876 7288 40889 7328
rect 40889 7288 40916 7328
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 7756 6784 7796 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 72748 6616 72788 6656
rect 82348 6616 82388 6656
rect 8140 6532 8180 6572
rect 98956 6616 98996 6656
rect 68812 6448 68852 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 35404 5776 35444 5816
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 35212 5272 35252 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 8524 5188 8564 5228
rect 35020 5188 35060 5228
rect 69196 5188 69236 5228
rect 7084 5104 7124 5144
rect 39436 5104 39476 5144
rect 71500 5104 71540 5144
rect 73516 4936 73556 4976
rect 35020 4768 35060 4808
rect 53740 4768 53780 4808
rect 49708 4684 49748 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 8332 4180 8372 4220
rect 32620 4096 32660 4136
rect 35212 4096 35252 4136
rect 35404 4096 35444 4136
rect 36748 4096 36788 4136
rect 37516 4096 37556 4136
rect 69100 4096 69140 4136
rect 8044 3844 8084 3884
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 8236 3172 8276 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 66220 2164 66260 2204
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 91084 1439 91121 1479
rect 91121 1439 91124 1479
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 5548 37988 5588 37997
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 5548 35981 5588 37948
rect 8524 37988 8564 37997
rect 5547 35972 5589 35981
rect 5547 35932 5548 35972
rect 5588 35932 5589 35972
rect 5547 35923 5589 35932
rect 843 35804 885 35813
rect 843 35764 844 35804
rect 884 35764 885 35804
rect 843 35755 885 35764
rect 844 24044 884 35755
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 5548 32948 5588 35923
rect 8236 35468 8276 35477
rect 8044 35300 8084 35309
rect 7852 35048 7892 35057
rect 5548 32899 5588 32908
rect 7084 34712 7124 34721
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 844 23995 884 24004
rect 940 24800 980 24809
rect 844 9428 884 9437
rect 844 4733 884 9388
rect 843 4724 885 4733
rect 843 4684 844 4724
rect 884 4684 885 4724
rect 843 4675 885 4684
rect 940 4145 980 24760
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 6412 21608 6452 21617
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 1228 15476 1268 15485
rect 1228 5069 1268 15436
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 6412 7505 6452 21568
rect 6411 7496 6453 7505
rect 6411 7456 6412 7496
rect 6452 7456 6453 7496
rect 6411 7447 6453 7456
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 7084 5144 7124 34672
rect 7756 31688 7796 31697
rect 7756 6824 7796 31648
rect 7852 28328 7892 35008
rect 7947 30344 7989 30353
rect 7947 30304 7948 30344
rect 7988 30304 7989 30344
rect 7947 30295 7989 30304
rect 7852 28279 7892 28288
rect 7948 17300 7988 30295
rect 7852 17260 7988 17300
rect 7852 16763 7892 17260
rect 7852 16714 7892 16723
rect 7756 6775 7796 6784
rect 7084 5095 7124 5104
rect 1227 5060 1269 5069
rect 1227 5020 1228 5060
rect 1268 5020 1269 5060
rect 1227 5011 1269 5020
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 939 4136 981 4145
rect 939 4096 940 4136
rect 980 4096 981 4136
rect 939 4087 981 4096
rect 8044 3884 8084 35260
rect 8140 32528 8180 32537
rect 8140 6572 8180 32488
rect 8140 6523 8180 6532
rect 8044 3835 8084 3844
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 8236 3212 8276 35428
rect 8332 35132 8372 35141
rect 8332 4220 8372 35092
rect 8524 5228 8564 37948
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 44523 35972 44565 35981
rect 44523 35932 44524 35972
rect 44564 35932 44565 35972
rect 44523 35923 44565 35932
rect 44524 35838 44564 35923
rect 69196 35888 69236 35897
rect 19276 35804 19316 35813
rect 19276 35552 19316 35764
rect 22635 35804 22677 35813
rect 22635 35764 22636 35804
rect 22676 35764 22677 35804
rect 22635 35755 22677 35764
rect 35500 35804 35540 35813
rect 22636 35670 22676 35755
rect 19276 35503 19316 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 17452 35132 17492 35141
rect 17260 34964 17300 34973
rect 17452 34964 17492 35092
rect 17300 34924 17492 34964
rect 17260 34915 17300 34924
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 35500 34544 35540 35764
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 35500 34495 35540 34504
rect 62380 34544 62420 34553
rect 62420 34504 62804 34544
rect 62380 34495 62420 34504
rect 62764 34376 62804 34504
rect 62764 34327 62804 34336
rect 10252 34208 10292 34217
rect 10252 31604 10292 34168
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 54700 33788 54740 33797
rect 54700 32453 54740 33748
rect 69100 32612 69140 32621
rect 54699 32444 54741 32453
rect 54699 32404 54700 32444
rect 54740 32404 54741 32444
rect 54699 32395 54741 32404
rect 68812 32444 68852 32453
rect 10252 31555 10292 31564
rect 50380 31772 50420 31781
rect 50380 30941 50420 31732
rect 50379 30932 50421 30941
rect 50379 30892 50380 30932
rect 50420 30892 50421 30932
rect 50379 30883 50421 30892
rect 53739 7832 53781 7841
rect 53739 7792 53740 7832
rect 53780 7792 53781 7832
rect 53739 7783 53781 7792
rect 40875 7496 40917 7505
rect 40875 7456 40876 7496
rect 40916 7456 40917 7496
rect 40875 7447 40917 7456
rect 40876 7328 40916 7447
rect 40876 7279 40916 7288
rect 35404 5816 35444 5825
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 35212 5312 35252 5321
rect 8524 5179 8564 5188
rect 35020 5228 35060 5237
rect 35020 4808 35060 5188
rect 35020 4759 35060 4768
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 8332 4171 8372 4180
rect 32619 4136 32661 4145
rect 32619 4096 32620 4136
rect 32660 4096 32661 4136
rect 32619 4087 32661 4096
rect 35212 4136 35252 5272
rect 35212 4087 35252 4096
rect 35404 4136 35444 5776
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 39435 5144 39477 5153
rect 39435 5104 39436 5144
rect 39476 5104 39477 5144
rect 39435 5095 39477 5104
rect 39436 5010 39476 5095
rect 53740 4808 53780 7783
rect 68812 6488 68852 32404
rect 68812 6439 68852 6448
rect 66219 5816 66261 5825
rect 66219 5776 66220 5816
rect 66260 5776 66261 5816
rect 66219 5767 66261 5776
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 53740 4759 53780 4768
rect 49707 4724 49749 4733
rect 49707 4684 49708 4724
rect 49748 4684 49749 4724
rect 49707 4675 49749 4684
rect 49708 4590 49748 4675
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 35404 4087 35444 4096
rect 36748 4136 36788 4145
rect 32620 4002 32660 4087
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 8236 3163 8276 3172
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 36748 1709 36788 4096
rect 37515 4136 37557 4145
rect 37515 4096 37516 4136
rect 37556 4096 37557 4136
rect 37515 4087 37557 4096
rect 37516 4002 37556 4087
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 66220 2204 66260 5767
rect 69100 4136 69140 32572
rect 69196 5228 69236 35848
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 99820 33200 99860 33209
rect 99860 33160 99956 33200
rect 99820 33151 99860 33160
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 97324 31445 97364 31530
rect 83499 31436 83541 31445
rect 83499 31396 83500 31436
rect 83540 31396 83541 31436
rect 83499 31387 83541 31396
rect 97323 31436 97365 31445
rect 97323 31395 97324 31436
rect 97364 31395 97365 31436
rect 97323 31387 97365 31395
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 83500 30848 83540 31387
rect 97324 31386 97364 31387
rect 83500 30799 83540 30808
rect 76971 30344 77013 30353
rect 76971 30304 76972 30344
rect 77012 30304 77013 30344
rect 76971 30295 77013 30304
rect 76972 16232 77012 30295
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 97324 29397 97364 29406
rect 97324 28757 97364 29357
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 84939 28748 84981 28757
rect 84939 28708 84940 28748
rect 84980 28708 84981 28748
rect 84939 28699 84981 28708
rect 97323 28748 97365 28757
rect 97323 28708 97324 28748
rect 97364 28708 97365 28748
rect 97323 28699 97365 28708
rect 84940 28614 84980 28699
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 80620 26144 80660 26153
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 80620 25136 80660 26104
rect 80620 25087 80660 25096
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 82924 23876 82964 23885
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 82924 17300 82964 23836
rect 99916 23876 99956 33160
rect 99916 23827 99956 23836
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 82828 17260 82964 17300
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 76972 16183 77012 16192
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 82828 9083 82868 17260
rect 98740 9213 98780 9222
rect 82828 9034 82868 9043
rect 98572 9173 98740 9176
rect 98572 9136 98780 9173
rect 72747 8924 72789 8933
rect 72747 8884 72748 8924
rect 72788 8884 72789 8924
rect 72747 8875 72789 8884
rect 71499 7916 71541 7925
rect 71499 7876 71500 7916
rect 71540 7876 71541 7916
rect 71499 7867 71541 7876
rect 69196 5179 69236 5188
rect 71500 5144 71540 7867
rect 72748 6656 72788 8875
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 98572 8009 98612 9136
rect 98740 9045 98780 9054
rect 98740 8933 98780 9005
rect 98739 8924 98781 8933
rect 98739 8884 98740 8924
rect 98780 8884 98781 8924
rect 98739 8875 98781 8884
rect 98860 8877 98900 8886
rect 73515 8000 73557 8009
rect 73515 7960 73516 8000
rect 73556 7960 73557 8000
rect 73515 7951 73557 7960
rect 98571 8000 98613 8009
rect 98571 7960 98572 8000
rect 98612 7960 98613 8000
rect 98571 7951 98613 7960
rect 72748 6607 72788 6616
rect 71500 5095 71540 5104
rect 73516 4976 73556 7951
rect 98860 7925 98900 8837
rect 98859 7916 98901 7925
rect 98859 7876 98860 7916
rect 98900 7876 98901 7916
rect 98859 7867 98901 7876
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 82347 6656 82389 6665
rect 82347 6616 82348 6656
rect 82388 6616 82389 6656
rect 82347 6607 82389 6616
rect 98955 6656 98997 6665
rect 98955 6616 98956 6656
rect 98996 6616 98997 6656
rect 98955 6607 98997 6616
rect 82348 6522 82388 6607
rect 98956 6522 98996 6607
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 73516 4927 73556 4936
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 69100 4087 69140 4096
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 66220 2155 66260 2164
rect 36747 1700 36789 1709
rect 36747 1660 36748 1700
rect 36788 1660 36789 1700
rect 36747 1651 36789 1660
rect 91083 1700 91125 1709
rect 91083 1660 91084 1700
rect 91124 1660 91125 1700
rect 91083 1651 91125 1660
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 91084 1479 91124 1651
rect 91084 1430 91124 1439
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 5548 35932 5588 35972
rect 844 35764 884 35804
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 844 4684 884 4724
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 6412 7456 6452 7496
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 7948 30304 7988 30344
rect 1228 5020 1268 5060
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 940 4096 980 4136
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 44524 35932 44564 35972
rect 22636 35764 22676 35804
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 54700 32404 54740 32444
rect 50380 30892 50420 30932
rect 53740 7792 53780 7832
rect 40876 7456 40916 7496
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 32620 4096 32660 4136
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 39436 5104 39476 5144
rect 66220 5776 66260 5816
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 49708 4684 49748 4724
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 37516 4096 37556 4136
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 83500 31396 83540 31436
rect 97324 31435 97364 31436
rect 97324 31396 97364 31435
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 76972 30304 77012 30344
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 84940 28708 84980 28748
rect 97324 28708 97364 28748
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 72748 8884 72788 8924
rect 71500 7876 71540 7916
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 98740 8884 98780 8924
rect 73516 7960 73556 8000
rect 98572 7960 98612 8000
rect 98860 7876 98900 7916
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 82348 6616 82388 6656
rect 98956 6616 98996 6656
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 36748 1660 36788 1700
rect 91084 1660 91124 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
<< metal5 >>
rect 4343 38576 4390 38618
rect 4514 38576 4558 38618
rect 4682 38576 4729 38618
rect 4343 38536 4352 38576
rect 4514 38536 4516 38576
rect 4556 38536 4558 38576
rect 4720 38536 4729 38576
rect 4343 38494 4390 38536
rect 4514 38494 4558 38536
rect 4682 38494 4729 38536
rect 19463 38576 19510 38618
rect 19634 38576 19678 38618
rect 19802 38576 19849 38618
rect 19463 38536 19472 38576
rect 19634 38536 19636 38576
rect 19676 38536 19678 38576
rect 19840 38536 19849 38576
rect 19463 38494 19510 38536
rect 19634 38494 19678 38536
rect 19802 38494 19849 38536
rect 34583 38576 34630 38618
rect 34754 38576 34798 38618
rect 34922 38576 34969 38618
rect 34583 38536 34592 38576
rect 34754 38536 34756 38576
rect 34796 38536 34798 38576
rect 34960 38536 34969 38576
rect 34583 38494 34630 38536
rect 34754 38494 34798 38536
rect 34922 38494 34969 38536
rect 49703 38576 49750 38618
rect 49874 38576 49918 38618
rect 50042 38576 50089 38618
rect 49703 38536 49712 38576
rect 49874 38536 49876 38576
rect 49916 38536 49918 38576
rect 50080 38536 50089 38576
rect 49703 38494 49750 38536
rect 49874 38494 49918 38536
rect 50042 38494 50089 38536
rect 64823 38576 64870 38618
rect 64994 38576 65038 38618
rect 65162 38576 65209 38618
rect 64823 38536 64832 38576
rect 64994 38536 64996 38576
rect 65036 38536 65038 38576
rect 65200 38536 65209 38576
rect 64823 38494 64870 38536
rect 64994 38494 65038 38536
rect 65162 38494 65209 38536
rect 79943 38576 79990 38618
rect 80114 38576 80158 38618
rect 80282 38576 80329 38618
rect 79943 38536 79952 38576
rect 80114 38536 80116 38576
rect 80156 38536 80158 38576
rect 80320 38536 80329 38576
rect 79943 38494 79990 38536
rect 80114 38494 80158 38536
rect 80282 38494 80329 38536
rect 3103 37820 3150 37862
rect 3274 37820 3318 37862
rect 3442 37820 3489 37862
rect 3103 37780 3112 37820
rect 3274 37780 3276 37820
rect 3316 37780 3318 37820
rect 3480 37780 3489 37820
rect 3103 37738 3150 37780
rect 3274 37738 3318 37780
rect 3442 37738 3489 37780
rect 18223 37820 18270 37862
rect 18394 37820 18438 37862
rect 18562 37820 18609 37862
rect 18223 37780 18232 37820
rect 18394 37780 18396 37820
rect 18436 37780 18438 37820
rect 18600 37780 18609 37820
rect 18223 37738 18270 37780
rect 18394 37738 18438 37780
rect 18562 37738 18609 37780
rect 33343 37820 33390 37862
rect 33514 37820 33558 37862
rect 33682 37820 33729 37862
rect 33343 37780 33352 37820
rect 33514 37780 33516 37820
rect 33556 37780 33558 37820
rect 33720 37780 33729 37820
rect 33343 37738 33390 37780
rect 33514 37738 33558 37780
rect 33682 37738 33729 37780
rect 48463 37820 48510 37862
rect 48634 37820 48678 37862
rect 48802 37820 48849 37862
rect 48463 37780 48472 37820
rect 48634 37780 48636 37820
rect 48676 37780 48678 37820
rect 48840 37780 48849 37820
rect 48463 37738 48510 37780
rect 48634 37738 48678 37780
rect 48802 37738 48849 37780
rect 63583 37820 63630 37862
rect 63754 37820 63798 37862
rect 63922 37820 63969 37862
rect 63583 37780 63592 37820
rect 63754 37780 63756 37820
rect 63796 37780 63798 37820
rect 63960 37780 63969 37820
rect 63583 37738 63630 37780
rect 63754 37738 63798 37780
rect 63922 37738 63969 37780
rect 78703 37820 78750 37862
rect 78874 37820 78918 37862
rect 79042 37820 79089 37862
rect 78703 37780 78712 37820
rect 78874 37780 78876 37820
rect 78916 37780 78918 37820
rect 79080 37780 79089 37820
rect 78703 37738 78750 37780
rect 78874 37738 78918 37780
rect 79042 37738 79089 37780
rect 4343 37064 4390 37106
rect 4514 37064 4558 37106
rect 4682 37064 4729 37106
rect 4343 37024 4352 37064
rect 4514 37024 4516 37064
rect 4556 37024 4558 37064
rect 4720 37024 4729 37064
rect 4343 36982 4390 37024
rect 4514 36982 4558 37024
rect 4682 36982 4729 37024
rect 19463 37064 19510 37106
rect 19634 37064 19678 37106
rect 19802 37064 19849 37106
rect 19463 37024 19472 37064
rect 19634 37024 19636 37064
rect 19676 37024 19678 37064
rect 19840 37024 19849 37064
rect 19463 36982 19510 37024
rect 19634 36982 19678 37024
rect 19802 36982 19849 37024
rect 34583 37064 34630 37106
rect 34754 37064 34798 37106
rect 34922 37064 34969 37106
rect 34583 37024 34592 37064
rect 34754 37024 34756 37064
rect 34796 37024 34798 37064
rect 34960 37024 34969 37064
rect 34583 36982 34630 37024
rect 34754 36982 34798 37024
rect 34922 36982 34969 37024
rect 49703 37064 49750 37106
rect 49874 37064 49918 37106
rect 50042 37064 50089 37106
rect 49703 37024 49712 37064
rect 49874 37024 49876 37064
rect 49916 37024 49918 37064
rect 50080 37024 50089 37064
rect 49703 36982 49750 37024
rect 49874 36982 49918 37024
rect 50042 36982 50089 37024
rect 64823 37064 64870 37106
rect 64994 37064 65038 37106
rect 65162 37064 65209 37106
rect 64823 37024 64832 37064
rect 64994 37024 64996 37064
rect 65036 37024 65038 37064
rect 65200 37024 65209 37064
rect 64823 36982 64870 37024
rect 64994 36982 65038 37024
rect 65162 36982 65209 37024
rect 79943 37064 79990 37106
rect 80114 37064 80158 37106
rect 80282 37064 80329 37106
rect 79943 37024 79952 37064
rect 80114 37024 80116 37064
rect 80156 37024 80158 37064
rect 80320 37024 80329 37064
rect 79943 36982 79990 37024
rect 80114 36982 80158 37024
rect 80282 36982 80329 37024
rect 3103 36308 3150 36350
rect 3274 36308 3318 36350
rect 3442 36308 3489 36350
rect 3103 36268 3112 36308
rect 3274 36268 3276 36308
rect 3316 36268 3318 36308
rect 3480 36268 3489 36308
rect 3103 36226 3150 36268
rect 3274 36226 3318 36268
rect 3442 36226 3489 36268
rect 18223 36308 18270 36350
rect 18394 36308 18438 36350
rect 18562 36308 18609 36350
rect 18223 36268 18232 36308
rect 18394 36268 18396 36308
rect 18436 36268 18438 36308
rect 18600 36268 18609 36308
rect 18223 36226 18270 36268
rect 18394 36226 18438 36268
rect 18562 36226 18609 36268
rect 33343 36308 33390 36350
rect 33514 36308 33558 36350
rect 33682 36308 33729 36350
rect 33343 36268 33352 36308
rect 33514 36268 33516 36308
rect 33556 36268 33558 36308
rect 33720 36268 33729 36308
rect 33343 36226 33390 36268
rect 33514 36226 33558 36268
rect 33682 36226 33729 36268
rect 48463 36308 48510 36350
rect 48634 36308 48678 36350
rect 48802 36308 48849 36350
rect 48463 36268 48472 36308
rect 48634 36268 48636 36308
rect 48676 36268 48678 36308
rect 48840 36268 48849 36308
rect 48463 36226 48510 36268
rect 48634 36226 48678 36268
rect 48802 36226 48849 36268
rect 63583 36308 63630 36350
rect 63754 36308 63798 36350
rect 63922 36308 63969 36350
rect 63583 36268 63592 36308
rect 63754 36268 63756 36308
rect 63796 36268 63798 36308
rect 63960 36268 63969 36308
rect 63583 36226 63630 36268
rect 63754 36226 63798 36268
rect 63922 36226 63969 36268
rect 78703 36308 78750 36350
rect 78874 36308 78918 36350
rect 79042 36308 79089 36350
rect 78703 36268 78712 36308
rect 78874 36268 78876 36308
rect 78916 36268 78918 36308
rect 79080 36268 79089 36308
rect 78703 36226 78750 36268
rect 78874 36226 78918 36268
rect 79042 36226 79089 36268
rect 5539 35932 5548 35972
rect 5588 35932 44524 35972
rect 44564 35932 44573 35972
rect 835 35764 844 35804
rect 884 35764 22636 35804
rect 22676 35764 22685 35804
rect 4343 35552 4390 35594
rect 4514 35552 4558 35594
rect 4682 35552 4729 35594
rect 4343 35512 4352 35552
rect 4514 35512 4516 35552
rect 4556 35512 4558 35552
rect 4720 35512 4729 35552
rect 4343 35470 4390 35512
rect 4514 35470 4558 35512
rect 4682 35470 4729 35512
rect 19463 35552 19510 35594
rect 19634 35552 19678 35594
rect 19802 35552 19849 35594
rect 19463 35512 19472 35552
rect 19634 35512 19636 35552
rect 19676 35512 19678 35552
rect 19840 35512 19849 35552
rect 19463 35470 19510 35512
rect 19634 35470 19678 35512
rect 19802 35470 19849 35512
rect 34583 35552 34630 35594
rect 34754 35552 34798 35594
rect 34922 35552 34969 35594
rect 34583 35512 34592 35552
rect 34754 35512 34756 35552
rect 34796 35512 34798 35552
rect 34960 35512 34969 35552
rect 34583 35470 34630 35512
rect 34754 35470 34798 35512
rect 34922 35470 34969 35512
rect 49703 35552 49750 35594
rect 49874 35552 49918 35594
rect 50042 35552 50089 35594
rect 49703 35512 49712 35552
rect 49874 35512 49876 35552
rect 49916 35512 49918 35552
rect 50080 35512 50089 35552
rect 49703 35470 49750 35512
rect 49874 35470 49918 35512
rect 50042 35470 50089 35512
rect 64823 35552 64870 35594
rect 64994 35552 65038 35594
rect 65162 35552 65209 35594
rect 64823 35512 64832 35552
rect 64994 35512 64996 35552
rect 65036 35512 65038 35552
rect 65200 35512 65209 35552
rect 64823 35470 64870 35512
rect 64994 35470 65038 35512
rect 65162 35470 65209 35512
rect 79943 35552 79990 35594
rect 80114 35552 80158 35594
rect 80282 35552 80329 35594
rect 79943 35512 79952 35552
rect 80114 35512 80116 35552
rect 80156 35512 80158 35552
rect 80320 35512 80329 35552
rect 79943 35470 79990 35512
rect 80114 35470 80158 35512
rect 80282 35470 80329 35512
rect 3103 34796 3150 34838
rect 3274 34796 3318 34838
rect 3442 34796 3489 34838
rect 3103 34756 3112 34796
rect 3274 34756 3276 34796
rect 3316 34756 3318 34796
rect 3480 34756 3489 34796
rect 3103 34714 3150 34756
rect 3274 34714 3318 34756
rect 3442 34714 3489 34756
rect 18223 34796 18270 34838
rect 18394 34796 18438 34838
rect 18562 34796 18609 34838
rect 18223 34756 18232 34796
rect 18394 34756 18396 34796
rect 18436 34756 18438 34796
rect 18600 34756 18609 34796
rect 18223 34714 18270 34756
rect 18394 34714 18438 34756
rect 18562 34714 18609 34756
rect 33343 34796 33390 34838
rect 33514 34796 33558 34838
rect 33682 34796 33729 34838
rect 33343 34756 33352 34796
rect 33514 34756 33516 34796
rect 33556 34756 33558 34796
rect 33720 34756 33729 34796
rect 33343 34714 33390 34756
rect 33514 34714 33558 34756
rect 33682 34714 33729 34756
rect 48463 34796 48510 34838
rect 48634 34796 48678 34838
rect 48802 34796 48849 34838
rect 48463 34756 48472 34796
rect 48634 34756 48636 34796
rect 48676 34756 48678 34796
rect 48840 34756 48849 34796
rect 48463 34714 48510 34756
rect 48634 34714 48678 34756
rect 48802 34714 48849 34756
rect 63583 34796 63630 34838
rect 63754 34796 63798 34838
rect 63922 34796 63969 34838
rect 63583 34756 63592 34796
rect 63754 34756 63756 34796
rect 63796 34756 63798 34796
rect 63960 34756 63969 34796
rect 63583 34714 63630 34756
rect 63754 34714 63798 34756
rect 63922 34714 63969 34756
rect 78703 34796 78750 34838
rect 78874 34796 78918 34838
rect 79042 34796 79089 34838
rect 78703 34756 78712 34796
rect 78874 34756 78876 34796
rect 78916 34756 78918 34796
rect 79080 34756 79089 34796
rect 78703 34714 78750 34756
rect 78874 34714 78918 34756
rect 79042 34714 79089 34756
rect 93796 34222 94236 34296
rect 93796 34098 93870 34222
rect 93994 34098 94038 34222
rect 94162 34098 94236 34222
rect 4343 34040 4390 34082
rect 4514 34040 4558 34082
rect 4682 34040 4729 34082
rect 4343 34000 4352 34040
rect 4514 34000 4516 34040
rect 4556 34000 4558 34040
rect 4720 34000 4729 34040
rect 4343 33958 4390 34000
rect 4514 33958 4558 34000
rect 4682 33958 4729 34000
rect 19463 34040 19510 34082
rect 19634 34040 19678 34082
rect 19802 34040 19849 34082
rect 19463 34000 19472 34040
rect 19634 34000 19636 34040
rect 19676 34000 19678 34040
rect 19840 34000 19849 34040
rect 19463 33958 19510 34000
rect 19634 33958 19678 34000
rect 19802 33958 19849 34000
rect 34583 34040 34630 34082
rect 34754 34040 34798 34082
rect 34922 34040 34969 34082
rect 34583 34000 34592 34040
rect 34754 34000 34756 34040
rect 34796 34000 34798 34040
rect 34960 34000 34969 34040
rect 34583 33958 34630 34000
rect 34754 33958 34798 34000
rect 34922 33958 34969 34000
rect 49703 34040 49750 34082
rect 49874 34040 49918 34082
rect 50042 34040 50089 34082
rect 49703 34000 49712 34040
rect 49874 34000 49876 34040
rect 49916 34000 49918 34040
rect 50080 34000 50089 34040
rect 49703 33958 49750 34000
rect 49874 33958 49918 34000
rect 50042 33958 50089 34000
rect 64823 34040 64870 34082
rect 64994 34040 65038 34082
rect 65162 34040 65209 34082
rect 64823 34000 64832 34040
rect 64994 34000 64996 34040
rect 65036 34000 65038 34040
rect 65200 34000 65209 34040
rect 64823 33958 64870 34000
rect 64994 33958 65038 34000
rect 65162 33958 65209 34000
rect 79943 34040 79990 34082
rect 80114 34040 80158 34082
rect 80282 34040 80329 34082
rect 79943 34000 79952 34040
rect 80114 34000 80116 34040
rect 80156 34000 80158 34040
rect 80320 34000 80329 34040
rect 79943 33958 79990 34000
rect 80114 33958 80158 34000
rect 80282 33958 80329 34000
rect 93796 34054 94236 34098
rect 93796 33930 93870 34054
rect 93994 33930 94038 34054
rect 94162 33930 94236 34054
rect 93796 33856 94236 33930
rect 3103 33284 3150 33326
rect 3274 33284 3318 33326
rect 3442 33284 3489 33326
rect 3103 33244 3112 33284
rect 3274 33244 3276 33284
rect 3316 33244 3318 33284
rect 3480 33244 3489 33284
rect 3103 33202 3150 33244
rect 3274 33202 3318 33244
rect 3442 33202 3489 33244
rect 78703 33284 78750 33326
rect 78874 33284 78918 33326
rect 79042 33284 79089 33326
rect 78703 33244 78712 33284
rect 78874 33244 78876 33284
rect 78916 33244 78918 33284
rect 79080 33244 79089 33284
rect 78703 33202 78750 33244
rect 78874 33202 78918 33244
rect 79042 33202 79089 33244
rect 4343 32528 4390 32570
rect 4514 32528 4558 32570
rect 4682 32528 4729 32570
rect 4343 32488 4352 32528
rect 4514 32488 4516 32528
rect 4556 32488 4558 32528
rect 4720 32488 4729 32528
rect 4343 32446 4390 32488
rect 4514 32446 4558 32488
rect 4682 32446 4729 32488
rect 79943 32528 79990 32570
rect 80114 32528 80158 32570
rect 80282 32528 80329 32570
rect 79943 32488 79952 32528
rect 80114 32488 80116 32528
rect 80156 32488 80158 32528
rect 80320 32488 80329 32528
rect 54691 32404 54700 32444
rect 54740 32404 67298 32444
rect 79943 32446 79990 32488
rect 80114 32446 80158 32488
rect 80282 32446 80329 32488
rect 3103 31772 3150 31814
rect 3274 31772 3318 31814
rect 3442 31772 3489 31814
rect 3103 31732 3112 31772
rect 3274 31732 3276 31772
rect 3316 31732 3318 31772
rect 3480 31732 3489 31772
rect 3103 31690 3150 31732
rect 3274 31690 3318 31732
rect 3442 31690 3489 31732
rect 78703 31772 78750 31814
rect 78874 31772 78918 31814
rect 79042 31772 79089 31814
rect 78703 31732 78712 31772
rect 78874 31732 78876 31772
rect 78916 31732 78918 31772
rect 79080 31732 79089 31772
rect 78703 31690 78750 31732
rect 78874 31690 78918 31732
rect 79042 31690 79089 31732
rect 83491 31396 83500 31436
rect 83540 31396 97324 31436
rect 97364 31396 97373 31436
rect 4343 31016 4390 31058
rect 4514 31016 4558 31058
rect 4682 31016 4729 31058
rect 4343 30976 4352 31016
rect 4514 30976 4516 31016
rect 4556 30976 4558 31016
rect 4720 30976 4729 31016
rect 4343 30934 4390 30976
rect 4514 30934 4558 30976
rect 4682 30934 4729 30976
rect 79943 31016 79990 31058
rect 80114 31016 80158 31058
rect 80282 31016 80329 31058
rect 79943 30976 79952 31016
rect 80114 30976 80116 31016
rect 80156 30976 80158 31016
rect 80320 30976 80329 31016
rect 50371 30892 50380 30932
rect 50420 30892 66386 30932
rect 79943 30934 79990 30976
rect 80114 30934 80158 30976
rect 80282 30934 80329 30976
rect 7939 30304 7948 30344
rect 7988 30304 76972 30344
rect 77012 30304 77021 30344
rect 3103 30260 3150 30302
rect 3274 30260 3318 30302
rect 3442 30260 3489 30302
rect 3103 30220 3112 30260
rect 3274 30220 3276 30260
rect 3316 30220 3318 30260
rect 3480 30220 3489 30260
rect 3103 30178 3150 30220
rect 3274 30178 3318 30220
rect 3442 30178 3489 30220
rect 78703 30260 78750 30302
rect 78874 30260 78918 30302
rect 79042 30260 79089 30302
rect 78703 30220 78712 30260
rect 78874 30220 78876 30260
rect 78916 30220 78918 30260
rect 79080 30220 79089 30260
rect 78703 30178 78750 30220
rect 78874 30178 78918 30220
rect 79042 30178 79089 30220
rect 4343 29504 4390 29546
rect 4514 29504 4558 29546
rect 4682 29504 4729 29546
rect 4343 29464 4352 29504
rect 4514 29464 4516 29504
rect 4556 29464 4558 29504
rect 4720 29464 4729 29504
rect 4343 29422 4390 29464
rect 4514 29422 4558 29464
rect 4682 29422 4729 29464
rect 79943 29504 79990 29546
rect 80114 29504 80158 29546
rect 80282 29504 80329 29546
rect 79943 29464 79952 29504
rect 80114 29464 80116 29504
rect 80156 29464 80158 29504
rect 80320 29464 80329 29504
rect 79943 29422 79990 29464
rect 80114 29422 80158 29464
rect 80282 29422 80329 29464
rect 95036 29462 95476 29536
rect 95036 29338 95110 29462
rect 95234 29338 95278 29462
rect 95402 29338 95476 29462
rect 95036 29294 95476 29338
rect 95036 29170 95110 29294
rect 95234 29170 95278 29294
rect 95402 29170 95476 29294
rect 95036 29096 95476 29170
rect 18196 29022 18636 29096
rect 18196 28898 18270 29022
rect 18394 28898 18438 29022
rect 18562 28898 18636 29022
rect 18196 28854 18636 28898
rect 3103 28748 3150 28790
rect 3274 28748 3318 28790
rect 3442 28748 3489 28790
rect 3103 28708 3112 28748
rect 3274 28708 3276 28748
rect 3316 28708 3318 28748
rect 3480 28708 3489 28748
rect 3103 28666 3150 28708
rect 3274 28666 3318 28708
rect 3442 28666 3489 28708
rect 18196 28730 18270 28854
rect 18394 28730 18438 28854
rect 18562 28730 18636 28854
rect 18196 28656 18636 28730
rect 33316 29022 33756 29096
rect 33316 28898 33390 29022
rect 33514 28898 33558 29022
rect 33682 28898 33756 29022
rect 33316 28854 33756 28898
rect 33316 28730 33390 28854
rect 33514 28730 33558 28854
rect 33682 28730 33756 28854
rect 33316 28656 33756 28730
rect 48436 29022 48876 29096
rect 48436 28898 48510 29022
rect 48634 28898 48678 29022
rect 48802 28898 48876 29022
rect 48436 28854 48876 28898
rect 48436 28730 48510 28854
rect 48634 28730 48678 28854
rect 48802 28730 48876 28854
rect 48436 28656 48876 28730
rect 63556 29022 63996 29096
rect 63556 28898 63630 29022
rect 63754 28898 63798 29022
rect 63922 28898 63996 29022
rect 63556 28854 63996 28898
rect 63556 28730 63630 28854
rect 63754 28730 63798 28854
rect 63922 28730 63996 28854
rect 63556 28656 63996 28730
rect 78703 28748 78750 28790
rect 78874 28748 78918 28790
rect 79042 28748 79089 28790
rect 78703 28708 78712 28748
rect 78874 28708 78876 28748
rect 78916 28708 78918 28748
rect 79080 28708 79089 28748
rect 84931 28708 84940 28748
rect 84980 28708 97324 28748
rect 97364 28708 97373 28748
rect 78703 28666 78750 28708
rect 78874 28666 78918 28708
rect 79042 28666 79089 28708
rect 93796 28222 94236 28296
rect 93796 28098 93870 28222
rect 93994 28098 94038 28222
rect 94162 28098 94236 28222
rect 93796 28054 94236 28098
rect 4343 27992 4390 28034
rect 4514 27992 4558 28034
rect 4682 27992 4729 28034
rect 4343 27952 4352 27992
rect 4514 27952 4516 27992
rect 4556 27952 4558 27992
rect 4720 27952 4729 27992
rect 4343 27910 4390 27952
rect 4514 27910 4558 27952
rect 4682 27910 4729 27952
rect 79943 27992 79990 28034
rect 80114 27992 80158 28034
rect 80282 27992 80329 28034
rect 79943 27952 79952 27992
rect 80114 27952 80116 27992
rect 80156 27952 80158 27992
rect 80320 27952 80329 27992
rect 79943 27910 79990 27952
rect 80114 27910 80158 27952
rect 80282 27910 80329 27952
rect 93796 27930 93870 28054
rect 93994 27930 94038 28054
rect 94162 27930 94236 28054
rect 93796 27856 94236 27930
rect 3103 27236 3150 27278
rect 3274 27236 3318 27278
rect 3442 27236 3489 27278
rect 3103 27196 3112 27236
rect 3274 27196 3276 27236
rect 3316 27196 3318 27236
rect 3480 27196 3489 27236
rect 3103 27154 3150 27196
rect 3274 27154 3318 27196
rect 3442 27154 3489 27196
rect 78703 27236 78750 27278
rect 78874 27236 78918 27278
rect 79042 27236 79089 27278
rect 78703 27196 78712 27236
rect 78874 27196 78876 27236
rect 78916 27196 78918 27236
rect 79080 27196 79089 27236
rect 78703 27154 78750 27196
rect 78874 27154 78918 27196
rect 79042 27154 79089 27196
rect 4343 26480 4390 26522
rect 4514 26480 4558 26522
rect 4682 26480 4729 26522
rect 4343 26440 4352 26480
rect 4514 26440 4516 26480
rect 4556 26440 4558 26480
rect 4720 26440 4729 26480
rect 4343 26398 4390 26440
rect 4514 26398 4558 26440
rect 4682 26398 4729 26440
rect 79943 26480 79990 26522
rect 80114 26480 80158 26522
rect 80282 26480 80329 26522
rect 79943 26440 79952 26480
rect 80114 26440 80116 26480
rect 80156 26440 80158 26480
rect 80320 26440 80329 26480
rect 79943 26398 79990 26440
rect 80114 26398 80158 26440
rect 80282 26398 80329 26440
rect 3103 25724 3150 25766
rect 3274 25724 3318 25766
rect 3442 25724 3489 25766
rect 3103 25684 3112 25724
rect 3274 25684 3276 25724
rect 3316 25684 3318 25724
rect 3480 25684 3489 25724
rect 3103 25642 3150 25684
rect 3274 25642 3318 25684
rect 3442 25642 3489 25684
rect 78703 25724 78750 25766
rect 78874 25724 78918 25766
rect 79042 25724 79089 25766
rect 78703 25684 78712 25724
rect 78874 25684 78876 25724
rect 78916 25684 78918 25724
rect 79080 25684 79089 25724
rect 78703 25642 78750 25684
rect 78874 25642 78918 25684
rect 79042 25642 79089 25684
rect 4343 24968 4390 25010
rect 4514 24968 4558 25010
rect 4682 24968 4729 25010
rect 4343 24928 4352 24968
rect 4514 24928 4516 24968
rect 4556 24928 4558 24968
rect 4720 24928 4729 24968
rect 4343 24886 4390 24928
rect 4514 24886 4558 24928
rect 4682 24886 4729 24928
rect 79943 24968 79990 25010
rect 80114 24968 80158 25010
rect 80282 24968 80329 25010
rect 79943 24928 79952 24968
rect 80114 24928 80116 24968
rect 80156 24928 80158 24968
rect 80320 24928 80329 24968
rect 79943 24886 79990 24928
rect 80114 24886 80158 24928
rect 80282 24886 80329 24928
rect 19436 24262 19876 24336
rect 3103 24212 3150 24254
rect 3274 24212 3318 24254
rect 3442 24212 3489 24254
rect 3103 24172 3112 24212
rect 3274 24172 3276 24212
rect 3316 24172 3318 24212
rect 3480 24172 3489 24212
rect 3103 24130 3150 24172
rect 3274 24130 3318 24172
rect 3442 24130 3489 24172
rect 19436 24138 19510 24262
rect 19634 24138 19678 24262
rect 19802 24138 19876 24262
rect 19436 24094 19876 24138
rect 19436 23970 19510 24094
rect 19634 23970 19678 24094
rect 19802 23970 19876 24094
rect 19436 23896 19876 23970
rect 34556 24262 34996 24336
rect 34556 24138 34630 24262
rect 34754 24138 34798 24262
rect 34922 24138 34996 24262
rect 34556 24094 34996 24138
rect 34556 23970 34630 24094
rect 34754 23970 34798 24094
rect 34922 23970 34996 24094
rect 34556 23896 34996 23970
rect 49676 24262 50116 24336
rect 49676 24138 49750 24262
rect 49874 24138 49918 24262
rect 50042 24138 50116 24262
rect 49676 24094 50116 24138
rect 49676 23970 49750 24094
rect 49874 23970 49918 24094
rect 50042 23970 50116 24094
rect 49676 23896 50116 23970
rect 64796 24262 65236 24336
rect 64796 24138 64870 24262
rect 64994 24138 65038 24262
rect 65162 24138 65236 24262
rect 64796 24094 65236 24138
rect 78703 24212 78750 24254
rect 78874 24212 78918 24254
rect 79042 24212 79089 24254
rect 78703 24172 78712 24212
rect 78874 24172 78876 24212
rect 78916 24172 78918 24212
rect 79080 24172 79089 24212
rect 78703 24130 78750 24172
rect 78874 24130 78918 24172
rect 79042 24130 79089 24172
rect 64796 23970 64870 24094
rect 64994 23970 65038 24094
rect 65162 23970 65236 24094
rect 64796 23896 65236 23970
rect 4343 23456 4390 23498
rect 4514 23456 4558 23498
rect 4682 23456 4729 23498
rect 4343 23416 4352 23456
rect 4514 23416 4516 23456
rect 4556 23416 4558 23456
rect 4720 23416 4729 23456
rect 4343 23374 4390 23416
rect 4514 23374 4558 23416
rect 4682 23374 4729 23416
rect 79943 23456 79990 23498
rect 80114 23456 80158 23498
rect 80282 23456 80329 23498
rect 79943 23416 79952 23456
rect 80114 23416 80116 23456
rect 80156 23416 80158 23456
rect 80320 23416 80329 23456
rect 79943 23374 79990 23416
rect 80114 23374 80158 23416
rect 80282 23374 80329 23416
rect 18196 23022 18636 23096
rect 18196 22898 18270 23022
rect 18394 22898 18438 23022
rect 18562 22898 18636 23022
rect 18196 22854 18636 22898
rect 3103 22700 3150 22742
rect 3274 22700 3318 22742
rect 3442 22700 3489 22742
rect 3103 22660 3112 22700
rect 3274 22660 3276 22700
rect 3316 22660 3318 22700
rect 3480 22660 3489 22700
rect 3103 22618 3150 22660
rect 3274 22618 3318 22660
rect 3442 22618 3489 22660
rect 18196 22730 18270 22854
rect 18394 22730 18438 22854
rect 18562 22730 18636 22854
rect 18196 22656 18636 22730
rect 33316 23022 33756 23096
rect 33316 22898 33390 23022
rect 33514 22898 33558 23022
rect 33682 22898 33756 23022
rect 33316 22854 33756 22898
rect 33316 22730 33390 22854
rect 33514 22730 33558 22854
rect 33682 22730 33756 22854
rect 33316 22656 33756 22730
rect 48436 23022 48876 23096
rect 48436 22898 48510 23022
rect 48634 22898 48678 23022
rect 48802 22898 48876 23022
rect 48436 22854 48876 22898
rect 48436 22730 48510 22854
rect 48634 22730 48678 22854
rect 48802 22730 48876 22854
rect 48436 22656 48876 22730
rect 63556 23022 63996 23096
rect 63556 22898 63630 23022
rect 63754 22898 63798 23022
rect 63922 22898 63996 23022
rect 63556 22854 63996 22898
rect 63556 22730 63630 22854
rect 63754 22730 63798 22854
rect 63922 22730 63996 22854
rect 63556 22656 63996 22730
rect 78703 22700 78750 22742
rect 78874 22700 78918 22742
rect 79042 22700 79089 22742
rect 78703 22660 78712 22700
rect 78874 22660 78876 22700
rect 78916 22660 78918 22700
rect 79080 22660 79089 22700
rect 78703 22618 78750 22660
rect 78874 22618 78918 22660
rect 79042 22618 79089 22660
rect 4343 21944 4390 21986
rect 4514 21944 4558 21986
rect 4682 21944 4729 21986
rect 4343 21904 4352 21944
rect 4514 21904 4516 21944
rect 4556 21904 4558 21944
rect 4720 21904 4729 21944
rect 4343 21862 4390 21904
rect 4514 21862 4558 21904
rect 4682 21862 4729 21904
rect 79943 21944 79990 21986
rect 80114 21944 80158 21986
rect 80282 21944 80329 21986
rect 79943 21904 79952 21944
rect 80114 21904 80116 21944
rect 80156 21904 80158 21944
rect 80320 21904 80329 21944
rect 79943 21862 79990 21904
rect 80114 21862 80158 21904
rect 80282 21862 80329 21904
rect 95063 21944 95110 21986
rect 95234 21944 95278 21986
rect 95402 21944 95449 21986
rect 95063 21904 95072 21944
rect 95234 21904 95236 21944
rect 95276 21904 95278 21944
rect 95440 21904 95449 21944
rect 95063 21862 95110 21904
rect 95234 21862 95278 21904
rect 95402 21862 95449 21904
rect 3103 21188 3150 21230
rect 3274 21188 3318 21230
rect 3442 21188 3489 21230
rect 3103 21148 3112 21188
rect 3274 21148 3276 21188
rect 3316 21148 3318 21188
rect 3480 21148 3489 21188
rect 3103 21106 3150 21148
rect 3274 21106 3318 21148
rect 3442 21106 3489 21148
rect 78703 21188 78750 21230
rect 78874 21188 78918 21230
rect 79042 21188 79089 21230
rect 78703 21148 78712 21188
rect 78874 21148 78876 21188
rect 78916 21148 78918 21188
rect 79080 21148 79089 21188
rect 78703 21106 78750 21148
rect 78874 21106 78918 21148
rect 79042 21106 79089 21148
rect 93823 21188 93870 21230
rect 93994 21188 94038 21230
rect 94162 21188 94209 21230
rect 93823 21148 93832 21188
rect 93994 21148 93996 21188
rect 94036 21148 94038 21188
rect 94200 21148 94209 21188
rect 93823 21106 93870 21148
rect 93994 21106 94038 21148
rect 94162 21106 94209 21148
rect 4343 20432 4390 20474
rect 4514 20432 4558 20474
rect 4682 20432 4729 20474
rect 4343 20392 4352 20432
rect 4514 20392 4516 20432
rect 4556 20392 4558 20432
rect 4720 20392 4729 20432
rect 4343 20350 4390 20392
rect 4514 20350 4558 20392
rect 4682 20350 4729 20392
rect 79943 20432 79990 20474
rect 80114 20432 80158 20474
rect 80282 20432 80329 20474
rect 79943 20392 79952 20432
rect 80114 20392 80116 20432
rect 80156 20392 80158 20432
rect 80320 20392 80329 20432
rect 79943 20350 79990 20392
rect 80114 20350 80158 20392
rect 80282 20350 80329 20392
rect 95063 20432 95110 20474
rect 95234 20432 95278 20474
rect 95402 20432 95449 20474
rect 95063 20392 95072 20432
rect 95234 20392 95236 20432
rect 95276 20392 95278 20432
rect 95440 20392 95449 20432
rect 95063 20350 95110 20392
rect 95234 20350 95278 20392
rect 95402 20350 95449 20392
rect 3103 19676 3150 19718
rect 3274 19676 3318 19718
rect 3442 19676 3489 19718
rect 3103 19636 3112 19676
rect 3274 19636 3276 19676
rect 3316 19636 3318 19676
rect 3480 19636 3489 19676
rect 3103 19594 3150 19636
rect 3274 19594 3318 19636
rect 3442 19594 3489 19636
rect 78703 19676 78750 19718
rect 78874 19676 78918 19718
rect 79042 19676 79089 19718
rect 78703 19636 78712 19676
rect 78874 19636 78876 19676
rect 78916 19636 78918 19676
rect 79080 19636 79089 19676
rect 78703 19594 78750 19636
rect 78874 19594 78918 19636
rect 79042 19594 79089 19636
rect 93823 19676 93870 19718
rect 93994 19676 94038 19718
rect 94162 19676 94209 19718
rect 93823 19636 93832 19676
rect 93994 19636 93996 19676
rect 94036 19636 94038 19676
rect 94200 19636 94209 19676
rect 93823 19594 93870 19636
rect 93994 19594 94038 19636
rect 94162 19594 94209 19636
rect 4343 18920 4390 18962
rect 4514 18920 4558 18962
rect 4682 18920 4729 18962
rect 4343 18880 4352 18920
rect 4514 18880 4516 18920
rect 4556 18880 4558 18920
rect 4720 18880 4729 18920
rect 4343 18838 4390 18880
rect 4514 18838 4558 18880
rect 4682 18838 4729 18880
rect 79943 18920 79990 18962
rect 80114 18920 80158 18962
rect 80282 18920 80329 18962
rect 79943 18880 79952 18920
rect 80114 18880 80116 18920
rect 80156 18880 80158 18920
rect 80320 18880 80329 18920
rect 79943 18838 79990 18880
rect 80114 18838 80158 18880
rect 80282 18838 80329 18880
rect 19436 18262 19876 18336
rect 3103 18164 3150 18206
rect 3274 18164 3318 18206
rect 3442 18164 3489 18206
rect 3103 18124 3112 18164
rect 3274 18124 3276 18164
rect 3316 18124 3318 18164
rect 3480 18124 3489 18164
rect 3103 18082 3150 18124
rect 3274 18082 3318 18124
rect 3442 18082 3489 18124
rect 19436 18138 19510 18262
rect 19634 18138 19678 18262
rect 19802 18138 19876 18262
rect 19436 18094 19876 18138
rect 19436 17970 19510 18094
rect 19634 17970 19678 18094
rect 19802 17970 19876 18094
rect 19436 17896 19876 17970
rect 34556 18262 34996 18336
rect 34556 18138 34630 18262
rect 34754 18138 34798 18262
rect 34922 18138 34996 18262
rect 34556 18094 34996 18138
rect 34556 17970 34630 18094
rect 34754 17970 34798 18094
rect 34922 17970 34996 18094
rect 34556 17896 34996 17970
rect 49676 18262 50116 18336
rect 49676 18138 49750 18262
rect 49874 18138 49918 18262
rect 50042 18138 50116 18262
rect 49676 18094 50116 18138
rect 49676 17970 49750 18094
rect 49874 17970 49918 18094
rect 50042 17970 50116 18094
rect 49676 17896 50116 17970
rect 64796 18262 65236 18336
rect 64796 18138 64870 18262
rect 64994 18138 65038 18262
rect 65162 18138 65236 18262
rect 64796 18094 65236 18138
rect 64796 17970 64870 18094
rect 64994 17970 65038 18094
rect 65162 17970 65236 18094
rect 78703 18164 78750 18206
rect 78874 18164 78918 18206
rect 79042 18164 79089 18206
rect 78703 18124 78712 18164
rect 78874 18124 78876 18164
rect 78916 18124 78918 18164
rect 79080 18124 79089 18164
rect 78703 18082 78750 18124
rect 78874 18082 78918 18124
rect 79042 18082 79089 18124
rect 64796 17896 65236 17970
rect 4343 17408 4390 17450
rect 4514 17408 4558 17450
rect 4682 17408 4729 17450
rect 4343 17368 4352 17408
rect 4514 17368 4516 17408
rect 4556 17368 4558 17408
rect 4720 17368 4729 17408
rect 4343 17326 4390 17368
rect 4514 17326 4558 17368
rect 4682 17326 4729 17368
rect 79943 17408 79990 17450
rect 80114 17408 80158 17450
rect 80282 17408 80329 17450
rect 79943 17368 79952 17408
rect 80114 17368 80116 17408
rect 80156 17368 80158 17408
rect 80320 17368 80329 17408
rect 79943 17326 79990 17368
rect 80114 17326 80158 17368
rect 80282 17326 80329 17368
rect 18196 17022 18636 17096
rect 18196 16898 18270 17022
rect 18394 16898 18438 17022
rect 18562 16898 18636 17022
rect 18196 16854 18636 16898
rect 18196 16730 18270 16854
rect 18394 16730 18438 16854
rect 18562 16730 18636 16854
rect 3103 16652 3150 16694
rect 3274 16652 3318 16694
rect 3442 16652 3489 16694
rect 18196 16656 18636 16730
rect 33316 17022 33756 17096
rect 33316 16898 33390 17022
rect 33514 16898 33558 17022
rect 33682 16898 33756 17022
rect 33316 16854 33756 16898
rect 33316 16730 33390 16854
rect 33514 16730 33558 16854
rect 33682 16730 33756 16854
rect 33316 16656 33756 16730
rect 48436 17022 48876 17096
rect 48436 16898 48510 17022
rect 48634 16898 48678 17022
rect 48802 16898 48876 17022
rect 48436 16854 48876 16898
rect 48436 16730 48510 16854
rect 48634 16730 48678 16854
rect 48802 16730 48876 16854
rect 48436 16656 48876 16730
rect 63556 17022 63996 17096
rect 63556 16898 63630 17022
rect 63754 16898 63798 17022
rect 63922 16898 63996 17022
rect 63556 16854 63996 16898
rect 63556 16730 63630 16854
rect 63754 16730 63798 16854
rect 63922 16730 63996 16854
rect 63556 16656 63996 16730
rect 3103 16612 3112 16652
rect 3274 16612 3276 16652
rect 3316 16612 3318 16652
rect 3480 16612 3489 16652
rect 3103 16570 3150 16612
rect 3274 16570 3318 16612
rect 3442 16570 3489 16612
rect 78703 16652 78750 16694
rect 78874 16652 78918 16694
rect 79042 16652 79089 16694
rect 78703 16612 78712 16652
rect 78874 16612 78876 16652
rect 78916 16612 78918 16652
rect 79080 16612 79089 16652
rect 78703 16570 78750 16612
rect 78874 16570 78918 16612
rect 79042 16570 79089 16612
rect 4343 15896 4390 15938
rect 4514 15896 4558 15938
rect 4682 15896 4729 15938
rect 4343 15856 4352 15896
rect 4514 15856 4516 15896
rect 4556 15856 4558 15896
rect 4720 15856 4729 15896
rect 4343 15814 4390 15856
rect 4514 15814 4558 15856
rect 4682 15814 4729 15856
rect 79943 15896 79990 15938
rect 80114 15896 80158 15938
rect 80282 15896 80329 15938
rect 79943 15856 79952 15896
rect 80114 15856 80116 15896
rect 80156 15856 80158 15896
rect 80320 15856 80329 15896
rect 79943 15814 79990 15856
rect 80114 15814 80158 15856
rect 80282 15814 80329 15856
rect 3103 15140 3150 15182
rect 3274 15140 3318 15182
rect 3442 15140 3489 15182
rect 3103 15100 3112 15140
rect 3274 15100 3276 15140
rect 3316 15100 3318 15140
rect 3480 15100 3489 15140
rect 3103 15058 3150 15100
rect 3274 15058 3318 15100
rect 3442 15058 3489 15100
rect 78703 15140 78750 15182
rect 78874 15140 78918 15182
rect 79042 15140 79089 15182
rect 78703 15100 78712 15140
rect 78874 15100 78876 15140
rect 78916 15100 78918 15140
rect 79080 15100 79089 15140
rect 78703 15058 78750 15100
rect 78874 15058 78918 15100
rect 79042 15058 79089 15100
rect 4343 14384 4390 14426
rect 4514 14384 4558 14426
rect 4682 14384 4729 14426
rect 4343 14344 4352 14384
rect 4514 14344 4516 14384
rect 4556 14344 4558 14384
rect 4720 14344 4729 14384
rect 4343 14302 4390 14344
rect 4514 14302 4558 14344
rect 4682 14302 4729 14344
rect 79943 14384 79990 14426
rect 80114 14384 80158 14426
rect 80282 14384 80329 14426
rect 79943 14344 79952 14384
rect 80114 14344 80116 14384
rect 80156 14344 80158 14384
rect 80320 14344 80329 14384
rect 79943 14302 79990 14344
rect 80114 14302 80158 14344
rect 80282 14302 80329 14344
rect 3103 13628 3150 13670
rect 3274 13628 3318 13670
rect 3442 13628 3489 13670
rect 3103 13588 3112 13628
rect 3274 13588 3276 13628
rect 3316 13588 3318 13628
rect 3480 13588 3489 13628
rect 3103 13546 3150 13588
rect 3274 13546 3318 13588
rect 3442 13546 3489 13588
rect 78703 13628 78750 13670
rect 78874 13628 78918 13670
rect 79042 13628 79089 13670
rect 78703 13588 78712 13628
rect 78874 13588 78876 13628
rect 78916 13588 78918 13628
rect 79080 13588 79089 13628
rect 78703 13546 78750 13588
rect 78874 13546 78918 13588
rect 79042 13546 79089 13588
rect 4343 12872 4390 12914
rect 4514 12872 4558 12914
rect 4682 12872 4729 12914
rect 4343 12832 4352 12872
rect 4514 12832 4516 12872
rect 4556 12832 4558 12872
rect 4720 12832 4729 12872
rect 4343 12790 4390 12832
rect 4514 12790 4558 12832
rect 4682 12790 4729 12832
rect 79943 12872 79990 12914
rect 80114 12872 80158 12914
rect 80282 12872 80329 12914
rect 79943 12832 79952 12872
rect 80114 12832 80116 12872
rect 80156 12832 80158 12872
rect 80320 12832 80329 12872
rect 79943 12790 79990 12832
rect 80114 12790 80158 12832
rect 80282 12790 80329 12832
rect 19436 12262 19876 12336
rect 3103 12116 3150 12158
rect 3274 12116 3318 12158
rect 3442 12116 3489 12158
rect 3103 12076 3112 12116
rect 3274 12076 3276 12116
rect 3316 12076 3318 12116
rect 3480 12076 3489 12116
rect 3103 12034 3150 12076
rect 3274 12034 3318 12076
rect 3442 12034 3489 12076
rect 19436 12138 19510 12262
rect 19634 12138 19678 12262
rect 19802 12138 19876 12262
rect 19436 12094 19876 12138
rect 19436 11970 19510 12094
rect 19634 11970 19678 12094
rect 19802 11970 19876 12094
rect 19436 11896 19876 11970
rect 34556 12262 34996 12336
rect 34556 12138 34630 12262
rect 34754 12138 34798 12262
rect 34922 12138 34996 12262
rect 34556 12094 34996 12138
rect 34556 11970 34630 12094
rect 34754 11970 34798 12094
rect 34922 11970 34996 12094
rect 34556 11896 34996 11970
rect 49676 12262 50116 12336
rect 49676 12138 49750 12262
rect 49874 12138 49918 12262
rect 50042 12138 50116 12262
rect 49676 12094 50116 12138
rect 49676 11970 49750 12094
rect 49874 11970 49918 12094
rect 50042 11970 50116 12094
rect 49676 11896 50116 11970
rect 64796 12262 65236 12336
rect 64796 12138 64870 12262
rect 64994 12138 65038 12262
rect 65162 12138 65236 12262
rect 95036 12262 95476 12336
rect 64796 12094 65236 12138
rect 64796 11970 64870 12094
rect 64994 11970 65038 12094
rect 65162 11970 65236 12094
rect 78703 12116 78750 12158
rect 78874 12116 78918 12158
rect 79042 12116 79089 12158
rect 78703 12076 78712 12116
rect 78874 12076 78876 12116
rect 78916 12076 78918 12116
rect 79080 12076 79089 12116
rect 78703 12034 78750 12076
rect 78874 12034 78918 12076
rect 79042 12034 79089 12076
rect 95036 12138 95110 12262
rect 95234 12138 95278 12262
rect 95402 12138 95476 12262
rect 95036 12094 95476 12138
rect 64796 11896 65236 11970
rect 95036 11970 95110 12094
rect 95234 11970 95278 12094
rect 95402 11970 95476 12094
rect 95036 11896 95476 11970
rect 4343 11360 4390 11402
rect 4514 11360 4558 11402
rect 4682 11360 4729 11402
rect 4343 11320 4352 11360
rect 4514 11320 4516 11360
rect 4556 11320 4558 11360
rect 4720 11320 4729 11360
rect 4343 11278 4390 11320
rect 4514 11278 4558 11320
rect 4682 11278 4729 11320
rect 79943 11360 79990 11402
rect 80114 11360 80158 11402
rect 80282 11360 80329 11402
rect 79943 11320 79952 11360
rect 80114 11320 80116 11360
rect 80156 11320 80158 11360
rect 80320 11320 80329 11360
rect 79943 11278 79990 11320
rect 80114 11278 80158 11320
rect 80282 11278 80329 11320
rect 18196 11022 18636 11096
rect 18196 10898 18270 11022
rect 18394 10898 18438 11022
rect 18562 10898 18636 11022
rect 18196 10854 18636 10898
rect 18196 10730 18270 10854
rect 18394 10730 18438 10854
rect 18562 10730 18636 10854
rect 18196 10656 18636 10730
rect 33316 11022 33756 11096
rect 33316 10898 33390 11022
rect 33514 10898 33558 11022
rect 33682 10898 33756 11022
rect 33316 10854 33756 10898
rect 33316 10730 33390 10854
rect 33514 10730 33558 10854
rect 33682 10730 33756 10854
rect 33316 10656 33756 10730
rect 48436 11022 48876 11096
rect 48436 10898 48510 11022
rect 48634 10898 48678 11022
rect 48802 10898 48876 11022
rect 48436 10854 48876 10898
rect 48436 10730 48510 10854
rect 48634 10730 48678 10854
rect 48802 10730 48876 10854
rect 48436 10656 48876 10730
rect 63556 11022 63996 11096
rect 63556 10898 63630 11022
rect 63754 10898 63798 11022
rect 63922 10898 63996 11022
rect 63556 10854 63996 10898
rect 63556 10730 63630 10854
rect 63754 10730 63798 10854
rect 63922 10730 63996 10854
rect 63556 10656 63996 10730
rect 93796 11022 94236 11096
rect 93796 10898 93870 11022
rect 93994 10898 94038 11022
rect 94162 10898 94236 11022
rect 93796 10854 94236 10898
rect 93796 10730 93870 10854
rect 93994 10730 94038 10854
rect 94162 10730 94236 10854
rect 93796 10656 94236 10730
rect 3103 10604 3150 10646
rect 3274 10604 3318 10646
rect 3442 10604 3489 10646
rect 3103 10564 3112 10604
rect 3274 10564 3276 10604
rect 3316 10564 3318 10604
rect 3480 10564 3489 10604
rect 3103 10522 3150 10564
rect 3274 10522 3318 10564
rect 3442 10522 3489 10564
rect 78703 10604 78750 10646
rect 78874 10604 78918 10646
rect 79042 10604 79089 10646
rect 78703 10564 78712 10604
rect 78874 10564 78876 10604
rect 78916 10564 78918 10604
rect 79080 10564 79089 10604
rect 78703 10522 78750 10564
rect 78874 10522 78918 10564
rect 79042 10522 79089 10564
rect 4343 9848 4390 9890
rect 4514 9848 4558 9890
rect 4682 9848 4729 9890
rect 4343 9808 4352 9848
rect 4514 9808 4516 9848
rect 4556 9808 4558 9848
rect 4720 9808 4729 9848
rect 4343 9766 4390 9808
rect 4514 9766 4558 9808
rect 4682 9766 4729 9808
rect 79943 9848 79990 9890
rect 80114 9848 80158 9890
rect 80282 9848 80329 9890
rect 79943 9808 79952 9848
rect 80114 9808 80116 9848
rect 80156 9808 80158 9848
rect 80320 9808 80329 9848
rect 79943 9766 79990 9808
rect 80114 9766 80158 9808
rect 80282 9766 80329 9808
rect 3103 9092 3150 9134
rect 3274 9092 3318 9134
rect 3442 9092 3489 9134
rect 3103 9052 3112 9092
rect 3274 9052 3276 9092
rect 3316 9052 3318 9092
rect 3480 9052 3489 9092
rect 3103 9010 3150 9052
rect 3274 9010 3318 9052
rect 3442 9010 3489 9052
rect 78703 9092 78750 9134
rect 78874 9092 78918 9134
rect 79042 9092 79089 9134
rect 78703 9052 78712 9092
rect 78874 9052 78876 9092
rect 78916 9052 78918 9092
rect 79080 9052 79089 9092
rect 78703 9010 78750 9052
rect 78874 9010 78918 9052
rect 79042 9010 79089 9052
rect 72739 8884 72748 8924
rect 72788 8884 98740 8924
rect 98780 8884 98789 8924
rect 4343 8336 4390 8378
rect 4514 8336 4558 8378
rect 4682 8336 4729 8378
rect 4343 8296 4352 8336
rect 4514 8296 4516 8336
rect 4556 8296 4558 8336
rect 4720 8296 4729 8336
rect 4343 8254 4390 8296
rect 4514 8254 4558 8296
rect 4682 8254 4729 8296
rect 79943 8336 79990 8378
rect 80114 8336 80158 8378
rect 80282 8336 80329 8378
rect 79943 8296 79952 8336
rect 80114 8296 80116 8336
rect 80156 8296 80158 8336
rect 80320 8296 80329 8336
rect 79943 8254 79990 8296
rect 80114 8254 80158 8296
rect 80282 8254 80329 8296
rect 73507 7960 73516 8000
rect 73556 7960 98572 8000
rect 98612 7960 98621 8000
rect 71491 7876 71500 7916
rect 71540 7876 98860 7916
rect 98900 7876 98909 7916
rect 53731 7792 53740 7832
rect 53780 7792 67298 7832
rect 3103 7580 3150 7622
rect 3274 7580 3318 7622
rect 3442 7580 3489 7622
rect 3103 7540 3112 7580
rect 3274 7540 3276 7580
rect 3316 7540 3318 7580
rect 3480 7540 3489 7580
rect 3103 7498 3150 7540
rect 3274 7498 3318 7540
rect 3442 7498 3489 7540
rect 78703 7580 78750 7622
rect 78874 7580 78918 7622
rect 79042 7580 79089 7622
rect 78703 7540 78712 7580
rect 78874 7540 78876 7580
rect 78916 7540 78918 7580
rect 79080 7540 79089 7580
rect 78703 7498 78750 7540
rect 78874 7498 78918 7540
rect 79042 7498 79089 7540
rect 6403 7456 6412 7496
rect 6452 7456 40876 7496
rect 40916 7456 40925 7496
rect 4343 6824 4390 6866
rect 4514 6824 4558 6866
rect 4682 6824 4729 6866
rect 4343 6784 4352 6824
rect 4514 6784 4516 6824
rect 4556 6784 4558 6824
rect 4720 6784 4729 6824
rect 4343 6742 4390 6784
rect 4514 6742 4558 6784
rect 4682 6742 4729 6784
rect 79943 6824 79990 6866
rect 80114 6824 80158 6866
rect 80282 6824 80329 6866
rect 79943 6784 79952 6824
rect 80114 6784 80116 6824
rect 80156 6784 80158 6824
rect 80320 6784 80329 6824
rect 79943 6742 79990 6784
rect 80114 6742 80158 6784
rect 80282 6742 80329 6784
rect 82339 6616 82348 6656
rect 82388 6616 98956 6656
rect 98996 6616 99005 6656
rect 95036 6262 95476 6336
rect 95036 6138 95110 6262
rect 95234 6138 95278 6262
rect 95402 6138 95476 6262
rect 3103 6068 3150 6110
rect 3274 6068 3318 6110
rect 3442 6068 3489 6110
rect 3103 6028 3112 6068
rect 3274 6028 3276 6068
rect 3316 6028 3318 6068
rect 3480 6028 3489 6068
rect 3103 5986 3150 6028
rect 3274 5986 3318 6028
rect 3442 5986 3489 6028
rect 78703 6068 78750 6110
rect 78874 6068 78918 6110
rect 79042 6068 79089 6110
rect 78703 6028 78712 6068
rect 78874 6028 78876 6068
rect 78916 6028 78918 6068
rect 79080 6028 79089 6068
rect 78703 5986 78750 6028
rect 78874 5986 78918 6028
rect 79042 5986 79089 6028
rect 95036 6094 95476 6138
rect 95036 5970 95110 6094
rect 95234 5970 95278 6094
rect 95402 5970 95476 6094
rect 95036 5896 95476 5970
rect 66211 5776 66220 5816
rect 66260 5776 66386 5816
rect 4343 5312 4390 5354
rect 4514 5312 4558 5354
rect 4682 5312 4729 5354
rect 4343 5272 4352 5312
rect 4514 5272 4516 5312
rect 4556 5272 4558 5312
rect 4720 5272 4729 5312
rect 4343 5230 4390 5272
rect 4514 5230 4558 5272
rect 4682 5230 4729 5272
rect 19463 5312 19510 5354
rect 19634 5312 19678 5354
rect 19802 5312 19849 5354
rect 19463 5272 19472 5312
rect 19634 5272 19636 5312
rect 19676 5272 19678 5312
rect 19840 5272 19849 5312
rect 19463 5230 19510 5272
rect 19634 5230 19678 5272
rect 19802 5230 19849 5272
rect 34583 5312 34630 5354
rect 34754 5312 34798 5354
rect 34922 5312 34969 5354
rect 34583 5272 34592 5312
rect 34754 5272 34756 5312
rect 34796 5272 34798 5312
rect 34960 5272 34969 5312
rect 34583 5230 34630 5272
rect 34754 5230 34798 5272
rect 34922 5230 34969 5272
rect 49703 5312 49750 5354
rect 49874 5312 49918 5354
rect 50042 5312 50089 5354
rect 49703 5272 49712 5312
rect 49874 5272 49876 5312
rect 49916 5272 49918 5312
rect 50080 5272 50089 5312
rect 49703 5230 49750 5272
rect 49874 5230 49918 5272
rect 50042 5230 50089 5272
rect 64823 5312 64870 5354
rect 64994 5312 65038 5354
rect 65162 5312 65209 5354
rect 64823 5272 64832 5312
rect 64994 5272 64996 5312
rect 65036 5272 65038 5312
rect 65200 5272 65209 5312
rect 64823 5230 64870 5272
rect 64994 5230 65038 5272
rect 65162 5230 65209 5272
rect 79943 5312 79990 5354
rect 80114 5312 80158 5354
rect 80282 5312 80329 5354
rect 79943 5272 79952 5312
rect 80114 5272 80116 5312
rect 80156 5272 80158 5312
rect 80320 5272 80329 5312
rect 79943 5230 79990 5272
rect 80114 5230 80158 5272
rect 80282 5230 80329 5272
rect 27340 5104 39436 5144
rect 39476 5104 39485 5144
rect 27340 5060 27380 5104
rect 1219 5020 1228 5060
rect 1268 5020 27380 5060
rect 93796 5022 94236 5096
rect 93796 4898 93870 5022
rect 93994 4898 94038 5022
rect 94162 4898 94236 5022
rect 93796 4854 94236 4898
rect 93796 4730 93870 4854
rect 93994 4730 94038 4854
rect 94162 4730 94236 4854
rect 835 4684 844 4724
rect 884 4684 49708 4724
rect 49748 4684 49757 4724
rect 93796 4656 94236 4730
rect 3103 4556 3150 4598
rect 3274 4556 3318 4598
rect 3442 4556 3489 4598
rect 3103 4516 3112 4556
rect 3274 4516 3276 4556
rect 3316 4516 3318 4556
rect 3480 4516 3489 4556
rect 3103 4474 3150 4516
rect 3274 4474 3318 4516
rect 3442 4474 3489 4516
rect 18223 4556 18270 4598
rect 18394 4556 18438 4598
rect 18562 4556 18609 4598
rect 18223 4516 18232 4556
rect 18394 4516 18396 4556
rect 18436 4516 18438 4556
rect 18600 4516 18609 4556
rect 18223 4474 18270 4516
rect 18394 4474 18438 4516
rect 18562 4474 18609 4516
rect 33343 4556 33390 4598
rect 33514 4556 33558 4598
rect 33682 4556 33729 4598
rect 33343 4516 33352 4556
rect 33514 4516 33516 4556
rect 33556 4516 33558 4556
rect 33720 4516 33729 4556
rect 33343 4474 33390 4516
rect 33514 4474 33558 4516
rect 33682 4474 33729 4516
rect 48463 4556 48510 4598
rect 48634 4556 48678 4598
rect 48802 4556 48849 4598
rect 48463 4516 48472 4556
rect 48634 4516 48636 4556
rect 48676 4516 48678 4556
rect 48840 4516 48849 4556
rect 48463 4474 48510 4516
rect 48634 4474 48678 4516
rect 48802 4474 48849 4516
rect 63583 4556 63630 4598
rect 63754 4556 63798 4598
rect 63922 4556 63969 4598
rect 63583 4516 63592 4556
rect 63754 4516 63756 4556
rect 63796 4516 63798 4556
rect 63960 4516 63969 4556
rect 63583 4474 63630 4516
rect 63754 4474 63798 4516
rect 63922 4474 63969 4516
rect 78703 4556 78750 4598
rect 78874 4556 78918 4598
rect 79042 4556 79089 4598
rect 78703 4516 78712 4556
rect 78874 4516 78876 4556
rect 78916 4516 78918 4556
rect 79080 4516 79089 4556
rect 78703 4474 78750 4516
rect 78874 4474 78918 4516
rect 79042 4474 79089 4516
rect 931 4096 940 4136
rect 980 4096 32620 4136
rect 32660 4096 37516 4136
rect 37556 4096 37565 4136
rect 4343 3800 4390 3842
rect 4514 3800 4558 3842
rect 4682 3800 4729 3842
rect 4343 3760 4352 3800
rect 4514 3760 4516 3800
rect 4556 3760 4558 3800
rect 4720 3760 4729 3800
rect 4343 3718 4390 3760
rect 4514 3718 4558 3760
rect 4682 3718 4729 3760
rect 19463 3800 19510 3842
rect 19634 3800 19678 3842
rect 19802 3800 19849 3842
rect 19463 3760 19472 3800
rect 19634 3760 19636 3800
rect 19676 3760 19678 3800
rect 19840 3760 19849 3800
rect 19463 3718 19510 3760
rect 19634 3718 19678 3760
rect 19802 3718 19849 3760
rect 34583 3800 34630 3842
rect 34754 3800 34798 3842
rect 34922 3800 34969 3842
rect 34583 3760 34592 3800
rect 34754 3760 34756 3800
rect 34796 3760 34798 3800
rect 34960 3760 34969 3800
rect 34583 3718 34630 3760
rect 34754 3718 34798 3760
rect 34922 3718 34969 3760
rect 49703 3800 49750 3842
rect 49874 3800 49918 3842
rect 50042 3800 50089 3842
rect 49703 3760 49712 3800
rect 49874 3760 49876 3800
rect 49916 3760 49918 3800
rect 50080 3760 50089 3800
rect 49703 3718 49750 3760
rect 49874 3718 49918 3760
rect 50042 3718 50089 3760
rect 64823 3800 64870 3842
rect 64994 3800 65038 3842
rect 65162 3800 65209 3842
rect 64823 3760 64832 3800
rect 64994 3760 64996 3800
rect 65036 3760 65038 3800
rect 65200 3760 65209 3800
rect 64823 3718 64870 3760
rect 64994 3718 65038 3760
rect 65162 3718 65209 3760
rect 79943 3800 79990 3842
rect 80114 3800 80158 3842
rect 80282 3800 80329 3842
rect 79943 3760 79952 3800
rect 80114 3760 80116 3800
rect 80156 3760 80158 3800
rect 80320 3760 80329 3800
rect 79943 3718 79990 3760
rect 80114 3718 80158 3760
rect 80282 3718 80329 3760
rect 3103 3044 3150 3086
rect 3274 3044 3318 3086
rect 3442 3044 3489 3086
rect 3103 3004 3112 3044
rect 3274 3004 3276 3044
rect 3316 3004 3318 3044
rect 3480 3004 3489 3044
rect 3103 2962 3150 3004
rect 3274 2962 3318 3004
rect 3442 2962 3489 3004
rect 18223 3044 18270 3086
rect 18394 3044 18438 3086
rect 18562 3044 18609 3086
rect 18223 3004 18232 3044
rect 18394 3004 18396 3044
rect 18436 3004 18438 3044
rect 18600 3004 18609 3044
rect 18223 2962 18270 3004
rect 18394 2962 18438 3004
rect 18562 2962 18609 3004
rect 33343 3044 33390 3086
rect 33514 3044 33558 3086
rect 33682 3044 33729 3086
rect 33343 3004 33352 3044
rect 33514 3004 33516 3044
rect 33556 3004 33558 3044
rect 33720 3004 33729 3044
rect 33343 2962 33390 3004
rect 33514 2962 33558 3004
rect 33682 2962 33729 3004
rect 48463 3044 48510 3086
rect 48634 3044 48678 3086
rect 48802 3044 48849 3086
rect 48463 3004 48472 3044
rect 48634 3004 48636 3044
rect 48676 3004 48678 3044
rect 48840 3004 48849 3044
rect 48463 2962 48510 3004
rect 48634 2962 48678 3004
rect 48802 2962 48849 3004
rect 63583 3044 63630 3086
rect 63754 3044 63798 3086
rect 63922 3044 63969 3086
rect 63583 3004 63592 3044
rect 63754 3004 63756 3044
rect 63796 3004 63798 3044
rect 63960 3004 63969 3044
rect 63583 2962 63630 3004
rect 63754 2962 63798 3004
rect 63922 2962 63969 3004
rect 78703 3044 78750 3086
rect 78874 3044 78918 3086
rect 79042 3044 79089 3086
rect 78703 3004 78712 3044
rect 78874 3004 78876 3044
rect 78916 3004 78918 3044
rect 79080 3004 79089 3044
rect 78703 2962 78750 3004
rect 78874 2962 78918 3004
rect 79042 2962 79089 3004
rect 4343 2288 4390 2330
rect 4514 2288 4558 2330
rect 4682 2288 4729 2330
rect 4343 2248 4352 2288
rect 4514 2248 4516 2288
rect 4556 2248 4558 2288
rect 4720 2248 4729 2288
rect 4343 2206 4390 2248
rect 4514 2206 4558 2248
rect 4682 2206 4729 2248
rect 19463 2288 19510 2330
rect 19634 2288 19678 2330
rect 19802 2288 19849 2330
rect 19463 2248 19472 2288
rect 19634 2248 19636 2288
rect 19676 2248 19678 2288
rect 19840 2248 19849 2288
rect 19463 2206 19510 2248
rect 19634 2206 19678 2248
rect 19802 2206 19849 2248
rect 34583 2288 34630 2330
rect 34754 2288 34798 2330
rect 34922 2288 34969 2330
rect 34583 2248 34592 2288
rect 34754 2248 34756 2288
rect 34796 2248 34798 2288
rect 34960 2248 34969 2288
rect 34583 2206 34630 2248
rect 34754 2206 34798 2248
rect 34922 2206 34969 2248
rect 49703 2288 49750 2330
rect 49874 2288 49918 2330
rect 50042 2288 50089 2330
rect 49703 2248 49712 2288
rect 49874 2248 49876 2288
rect 49916 2248 49918 2288
rect 50080 2248 50089 2288
rect 49703 2206 49750 2248
rect 49874 2206 49918 2248
rect 50042 2206 50089 2248
rect 64823 2288 64870 2330
rect 64994 2288 65038 2330
rect 65162 2288 65209 2330
rect 64823 2248 64832 2288
rect 64994 2248 64996 2288
rect 65036 2248 65038 2288
rect 65200 2248 65209 2288
rect 64823 2206 64870 2248
rect 64994 2206 65038 2248
rect 65162 2206 65209 2248
rect 79943 2288 79990 2330
rect 80114 2288 80158 2330
rect 80282 2288 80329 2330
rect 79943 2248 79952 2288
rect 80114 2248 80116 2288
rect 80156 2248 80158 2288
rect 80320 2248 80329 2288
rect 79943 2206 79990 2248
rect 80114 2206 80158 2248
rect 80282 2206 80329 2248
rect 36739 1660 36748 1700
rect 36788 1660 91084 1700
rect 91124 1660 91133 1700
rect 3103 1532 3150 1574
rect 3274 1532 3318 1574
rect 3442 1532 3489 1574
rect 3103 1492 3112 1532
rect 3274 1492 3276 1532
rect 3316 1492 3318 1532
rect 3480 1492 3489 1532
rect 3103 1450 3150 1492
rect 3274 1450 3318 1492
rect 3442 1450 3489 1492
rect 18223 1532 18270 1574
rect 18394 1532 18438 1574
rect 18562 1532 18609 1574
rect 18223 1492 18232 1532
rect 18394 1492 18396 1532
rect 18436 1492 18438 1532
rect 18600 1492 18609 1532
rect 18223 1450 18270 1492
rect 18394 1450 18438 1492
rect 18562 1450 18609 1492
rect 33343 1532 33390 1574
rect 33514 1532 33558 1574
rect 33682 1532 33729 1574
rect 33343 1492 33352 1532
rect 33514 1492 33516 1532
rect 33556 1492 33558 1532
rect 33720 1492 33729 1532
rect 33343 1450 33390 1492
rect 33514 1450 33558 1492
rect 33682 1450 33729 1492
rect 48463 1532 48510 1574
rect 48634 1532 48678 1574
rect 48802 1532 48849 1574
rect 48463 1492 48472 1532
rect 48634 1492 48636 1532
rect 48676 1492 48678 1532
rect 48840 1492 48849 1532
rect 48463 1450 48510 1492
rect 48634 1450 48678 1492
rect 48802 1450 48849 1492
rect 63583 1532 63630 1574
rect 63754 1532 63798 1574
rect 63922 1532 63969 1574
rect 63583 1492 63592 1532
rect 63754 1492 63756 1532
rect 63796 1492 63798 1532
rect 63960 1492 63969 1532
rect 63583 1450 63630 1492
rect 63754 1450 63798 1492
rect 63922 1450 63969 1492
rect 78703 1532 78750 1574
rect 78874 1532 78918 1574
rect 79042 1532 79089 1574
rect 78703 1492 78712 1532
rect 78874 1492 78876 1532
rect 78916 1492 78918 1532
rect 79080 1492 79089 1532
rect 78703 1450 78750 1492
rect 78874 1450 78918 1492
rect 79042 1450 79089 1492
rect 4343 776 4390 818
rect 4514 776 4558 818
rect 4682 776 4729 818
rect 4343 736 4352 776
rect 4514 736 4516 776
rect 4556 736 4558 776
rect 4720 736 4729 776
rect 4343 694 4390 736
rect 4514 694 4558 736
rect 4682 694 4729 736
rect 19463 776 19510 818
rect 19634 776 19678 818
rect 19802 776 19849 818
rect 19463 736 19472 776
rect 19634 736 19636 776
rect 19676 736 19678 776
rect 19840 736 19849 776
rect 19463 694 19510 736
rect 19634 694 19678 736
rect 19802 694 19849 736
rect 34583 776 34630 818
rect 34754 776 34798 818
rect 34922 776 34969 818
rect 34583 736 34592 776
rect 34754 736 34756 776
rect 34796 736 34798 776
rect 34960 736 34969 776
rect 34583 694 34630 736
rect 34754 694 34798 736
rect 34922 694 34969 736
rect 49703 776 49750 818
rect 49874 776 49918 818
rect 50042 776 50089 818
rect 49703 736 49712 776
rect 49874 736 49876 776
rect 49916 736 49918 776
rect 50080 736 50089 776
rect 49703 694 49750 736
rect 49874 694 49918 736
rect 50042 694 50089 736
rect 64823 776 64870 818
rect 64994 776 65038 818
rect 65162 776 65209 818
rect 64823 736 64832 776
rect 64994 736 64996 776
rect 65036 736 65038 776
rect 65200 736 65209 776
rect 64823 694 64870 736
rect 64994 694 65038 736
rect 65162 694 65209 736
rect 79943 776 79990 818
rect 80114 776 80158 818
rect 80282 776 80329 818
rect 79943 736 79952 776
rect 80114 736 80116 776
rect 80156 736 80158 776
rect 80320 736 80329 776
rect 79943 694 79990 736
rect 80114 694 80158 736
rect 80282 694 80329 736
<< via5 >>
rect 4390 38576 4514 38618
rect 4558 38576 4682 38618
rect 4390 38536 4392 38576
rect 4392 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4514 38576
rect 4558 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4680 38576
rect 4680 38536 4682 38576
rect 4390 38494 4514 38536
rect 4558 38494 4682 38536
rect 19510 38576 19634 38618
rect 19678 38576 19802 38618
rect 19510 38536 19512 38576
rect 19512 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19634 38576
rect 19678 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19800 38576
rect 19800 38536 19802 38576
rect 19510 38494 19634 38536
rect 19678 38494 19802 38536
rect 34630 38576 34754 38618
rect 34798 38576 34922 38618
rect 34630 38536 34632 38576
rect 34632 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34754 38576
rect 34798 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34920 38576
rect 34920 38536 34922 38576
rect 34630 38494 34754 38536
rect 34798 38494 34922 38536
rect 49750 38576 49874 38618
rect 49918 38576 50042 38618
rect 49750 38536 49752 38576
rect 49752 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49874 38576
rect 49918 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50040 38576
rect 50040 38536 50042 38576
rect 49750 38494 49874 38536
rect 49918 38494 50042 38536
rect 64870 38576 64994 38618
rect 65038 38576 65162 38618
rect 64870 38536 64872 38576
rect 64872 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64994 38576
rect 65038 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65160 38576
rect 65160 38536 65162 38576
rect 64870 38494 64994 38536
rect 65038 38494 65162 38536
rect 79990 38576 80114 38618
rect 80158 38576 80282 38618
rect 79990 38536 79992 38576
rect 79992 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80114 38576
rect 80158 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80280 38576
rect 80280 38536 80282 38576
rect 79990 38494 80114 38536
rect 80158 38494 80282 38536
rect 3150 37820 3274 37862
rect 3318 37820 3442 37862
rect 3150 37780 3152 37820
rect 3152 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3274 37820
rect 3318 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3440 37820
rect 3440 37780 3442 37820
rect 3150 37738 3274 37780
rect 3318 37738 3442 37780
rect 18270 37820 18394 37862
rect 18438 37820 18562 37862
rect 18270 37780 18272 37820
rect 18272 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18394 37820
rect 18438 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18560 37820
rect 18560 37780 18562 37820
rect 18270 37738 18394 37780
rect 18438 37738 18562 37780
rect 33390 37820 33514 37862
rect 33558 37820 33682 37862
rect 33390 37780 33392 37820
rect 33392 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33514 37820
rect 33558 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33680 37820
rect 33680 37780 33682 37820
rect 33390 37738 33514 37780
rect 33558 37738 33682 37780
rect 48510 37820 48634 37862
rect 48678 37820 48802 37862
rect 48510 37780 48512 37820
rect 48512 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48634 37820
rect 48678 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48800 37820
rect 48800 37780 48802 37820
rect 48510 37738 48634 37780
rect 48678 37738 48802 37780
rect 63630 37820 63754 37862
rect 63798 37820 63922 37862
rect 63630 37780 63632 37820
rect 63632 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63754 37820
rect 63798 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63920 37820
rect 63920 37780 63922 37820
rect 63630 37738 63754 37780
rect 63798 37738 63922 37780
rect 78750 37820 78874 37862
rect 78918 37820 79042 37862
rect 78750 37780 78752 37820
rect 78752 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78874 37820
rect 78918 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79040 37820
rect 79040 37780 79042 37820
rect 78750 37738 78874 37780
rect 78918 37738 79042 37780
rect 4390 37064 4514 37106
rect 4558 37064 4682 37106
rect 4390 37024 4392 37064
rect 4392 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4514 37064
rect 4558 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4680 37064
rect 4680 37024 4682 37064
rect 4390 36982 4514 37024
rect 4558 36982 4682 37024
rect 19510 37064 19634 37106
rect 19678 37064 19802 37106
rect 19510 37024 19512 37064
rect 19512 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19634 37064
rect 19678 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19800 37064
rect 19800 37024 19802 37064
rect 19510 36982 19634 37024
rect 19678 36982 19802 37024
rect 34630 37064 34754 37106
rect 34798 37064 34922 37106
rect 34630 37024 34632 37064
rect 34632 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34754 37064
rect 34798 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34920 37064
rect 34920 37024 34922 37064
rect 34630 36982 34754 37024
rect 34798 36982 34922 37024
rect 49750 37064 49874 37106
rect 49918 37064 50042 37106
rect 49750 37024 49752 37064
rect 49752 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49874 37064
rect 49918 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50040 37064
rect 50040 37024 50042 37064
rect 49750 36982 49874 37024
rect 49918 36982 50042 37024
rect 64870 37064 64994 37106
rect 65038 37064 65162 37106
rect 64870 37024 64872 37064
rect 64872 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64994 37064
rect 65038 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65160 37064
rect 65160 37024 65162 37064
rect 64870 36982 64994 37024
rect 65038 36982 65162 37024
rect 79990 37064 80114 37106
rect 80158 37064 80282 37106
rect 79990 37024 79992 37064
rect 79992 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80114 37064
rect 80158 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80280 37064
rect 80280 37024 80282 37064
rect 79990 36982 80114 37024
rect 80158 36982 80282 37024
rect 3150 36308 3274 36350
rect 3318 36308 3442 36350
rect 3150 36268 3152 36308
rect 3152 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3274 36308
rect 3318 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3440 36308
rect 3440 36268 3442 36308
rect 3150 36226 3274 36268
rect 3318 36226 3442 36268
rect 18270 36308 18394 36350
rect 18438 36308 18562 36350
rect 18270 36268 18272 36308
rect 18272 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18394 36308
rect 18438 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18560 36308
rect 18560 36268 18562 36308
rect 18270 36226 18394 36268
rect 18438 36226 18562 36268
rect 33390 36308 33514 36350
rect 33558 36308 33682 36350
rect 33390 36268 33392 36308
rect 33392 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33514 36308
rect 33558 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33680 36308
rect 33680 36268 33682 36308
rect 33390 36226 33514 36268
rect 33558 36226 33682 36268
rect 48510 36308 48634 36350
rect 48678 36308 48802 36350
rect 48510 36268 48512 36308
rect 48512 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48634 36308
rect 48678 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48800 36308
rect 48800 36268 48802 36308
rect 48510 36226 48634 36268
rect 48678 36226 48802 36268
rect 63630 36308 63754 36350
rect 63798 36308 63922 36350
rect 63630 36268 63632 36308
rect 63632 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63754 36308
rect 63798 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63920 36308
rect 63920 36268 63922 36308
rect 63630 36226 63754 36268
rect 63798 36226 63922 36268
rect 78750 36308 78874 36350
rect 78918 36308 79042 36350
rect 78750 36268 78752 36308
rect 78752 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78874 36308
rect 78918 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79040 36308
rect 79040 36268 79042 36308
rect 78750 36226 78874 36268
rect 78918 36226 79042 36268
rect 4390 35552 4514 35594
rect 4558 35552 4682 35594
rect 4390 35512 4392 35552
rect 4392 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4514 35552
rect 4558 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4680 35552
rect 4680 35512 4682 35552
rect 4390 35470 4514 35512
rect 4558 35470 4682 35512
rect 19510 35552 19634 35594
rect 19678 35552 19802 35594
rect 19510 35512 19512 35552
rect 19512 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19634 35552
rect 19678 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19800 35552
rect 19800 35512 19802 35552
rect 19510 35470 19634 35512
rect 19678 35470 19802 35512
rect 34630 35552 34754 35594
rect 34798 35552 34922 35594
rect 34630 35512 34632 35552
rect 34632 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34754 35552
rect 34798 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34920 35552
rect 34920 35512 34922 35552
rect 34630 35470 34754 35512
rect 34798 35470 34922 35512
rect 49750 35552 49874 35594
rect 49918 35552 50042 35594
rect 49750 35512 49752 35552
rect 49752 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49874 35552
rect 49918 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50040 35552
rect 50040 35512 50042 35552
rect 49750 35470 49874 35512
rect 49918 35470 50042 35512
rect 64870 35552 64994 35594
rect 65038 35552 65162 35594
rect 64870 35512 64872 35552
rect 64872 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64994 35552
rect 65038 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65160 35552
rect 65160 35512 65162 35552
rect 64870 35470 64994 35512
rect 65038 35470 65162 35512
rect 79990 35552 80114 35594
rect 80158 35552 80282 35594
rect 79990 35512 79992 35552
rect 79992 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80114 35552
rect 80158 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80280 35552
rect 80280 35512 80282 35552
rect 79990 35470 80114 35512
rect 80158 35470 80282 35512
rect 3150 34796 3274 34838
rect 3318 34796 3442 34838
rect 3150 34756 3152 34796
rect 3152 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3274 34796
rect 3318 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3440 34796
rect 3440 34756 3442 34796
rect 3150 34714 3274 34756
rect 3318 34714 3442 34756
rect 18270 34796 18394 34838
rect 18438 34796 18562 34838
rect 18270 34756 18272 34796
rect 18272 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18394 34796
rect 18438 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18560 34796
rect 18560 34756 18562 34796
rect 18270 34714 18394 34756
rect 18438 34714 18562 34756
rect 33390 34796 33514 34838
rect 33558 34796 33682 34838
rect 33390 34756 33392 34796
rect 33392 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33514 34796
rect 33558 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33680 34796
rect 33680 34756 33682 34796
rect 33390 34714 33514 34756
rect 33558 34714 33682 34756
rect 48510 34796 48634 34838
rect 48678 34796 48802 34838
rect 48510 34756 48512 34796
rect 48512 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48634 34796
rect 48678 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48800 34796
rect 48800 34756 48802 34796
rect 48510 34714 48634 34756
rect 48678 34714 48802 34756
rect 63630 34796 63754 34838
rect 63798 34796 63922 34838
rect 63630 34756 63632 34796
rect 63632 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63754 34796
rect 63798 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63920 34796
rect 63920 34756 63922 34796
rect 63630 34714 63754 34756
rect 63798 34714 63922 34756
rect 78750 34796 78874 34838
rect 78918 34796 79042 34838
rect 78750 34756 78752 34796
rect 78752 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78874 34796
rect 78918 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79040 34796
rect 79040 34756 79042 34796
rect 78750 34714 78874 34756
rect 78918 34714 79042 34756
rect 93870 34098 93994 34222
rect 94038 34098 94162 34222
rect 4390 34040 4514 34082
rect 4558 34040 4682 34082
rect 4390 34000 4392 34040
rect 4392 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4514 34040
rect 4558 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4680 34040
rect 4680 34000 4682 34040
rect 4390 33958 4514 34000
rect 4558 33958 4682 34000
rect 19510 34040 19634 34082
rect 19678 34040 19802 34082
rect 19510 34000 19512 34040
rect 19512 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19634 34040
rect 19678 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19800 34040
rect 19800 34000 19802 34040
rect 19510 33958 19634 34000
rect 19678 33958 19802 34000
rect 34630 34040 34754 34082
rect 34798 34040 34922 34082
rect 34630 34000 34632 34040
rect 34632 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34754 34040
rect 34798 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34920 34040
rect 34920 34000 34922 34040
rect 34630 33958 34754 34000
rect 34798 33958 34922 34000
rect 49750 34040 49874 34082
rect 49918 34040 50042 34082
rect 49750 34000 49752 34040
rect 49752 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49874 34040
rect 49918 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50040 34040
rect 50040 34000 50042 34040
rect 49750 33958 49874 34000
rect 49918 33958 50042 34000
rect 64870 34040 64994 34082
rect 65038 34040 65162 34082
rect 64870 34000 64872 34040
rect 64872 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64994 34040
rect 65038 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65160 34040
rect 65160 34000 65162 34040
rect 64870 33958 64994 34000
rect 65038 33958 65162 34000
rect 79990 34040 80114 34082
rect 80158 34040 80282 34082
rect 79990 34000 79992 34040
rect 79992 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80114 34040
rect 80158 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80280 34040
rect 80280 34000 80282 34040
rect 79990 33958 80114 34000
rect 80158 33958 80282 34000
rect 93870 33930 93994 34054
rect 94038 33930 94162 34054
rect 3150 33284 3274 33326
rect 3318 33284 3442 33326
rect 3150 33244 3152 33284
rect 3152 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3274 33284
rect 3318 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3440 33284
rect 3440 33244 3442 33284
rect 3150 33202 3274 33244
rect 3318 33202 3442 33244
rect 78750 33284 78874 33326
rect 78918 33284 79042 33326
rect 78750 33244 78752 33284
rect 78752 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78874 33284
rect 78918 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79040 33284
rect 79040 33244 79042 33284
rect 78750 33202 78874 33244
rect 78918 33202 79042 33244
rect 4390 32528 4514 32570
rect 4558 32528 4682 32570
rect 4390 32488 4392 32528
rect 4392 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4514 32528
rect 4558 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4680 32528
rect 4680 32488 4682 32528
rect 4390 32446 4514 32488
rect 4558 32446 4682 32488
rect 79990 32528 80114 32570
rect 80158 32528 80282 32570
rect 79990 32488 79992 32528
rect 79992 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80114 32528
rect 80158 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80280 32528
rect 80280 32488 80282 32528
rect 67298 32362 67422 32486
rect 79990 32446 80114 32488
rect 80158 32446 80282 32488
rect 3150 31772 3274 31814
rect 3318 31772 3442 31814
rect 3150 31732 3152 31772
rect 3152 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3274 31772
rect 3318 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3440 31772
rect 3440 31732 3442 31772
rect 3150 31690 3274 31732
rect 3318 31690 3442 31732
rect 78750 31772 78874 31814
rect 78918 31772 79042 31814
rect 78750 31732 78752 31772
rect 78752 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78874 31772
rect 78918 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79040 31772
rect 79040 31732 79042 31772
rect 78750 31690 78874 31732
rect 78918 31690 79042 31732
rect 4390 31016 4514 31058
rect 4558 31016 4682 31058
rect 4390 30976 4392 31016
rect 4392 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4514 31016
rect 4558 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4680 31016
rect 4680 30976 4682 31016
rect 4390 30934 4514 30976
rect 4558 30934 4682 30976
rect 79990 31016 80114 31058
rect 80158 31016 80282 31058
rect 79990 30976 79992 31016
rect 79992 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80114 31016
rect 80158 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80280 31016
rect 80280 30976 80282 31016
rect 66386 30850 66510 30974
rect 79990 30934 80114 30976
rect 80158 30934 80282 30976
rect 3150 30260 3274 30302
rect 3318 30260 3442 30302
rect 3150 30220 3152 30260
rect 3152 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3274 30260
rect 3318 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3440 30260
rect 3440 30220 3442 30260
rect 3150 30178 3274 30220
rect 3318 30178 3442 30220
rect 78750 30260 78874 30302
rect 78918 30260 79042 30302
rect 78750 30220 78752 30260
rect 78752 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78874 30260
rect 78918 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79040 30260
rect 79040 30220 79042 30260
rect 78750 30178 78874 30220
rect 78918 30178 79042 30220
rect 4390 29504 4514 29546
rect 4558 29504 4682 29546
rect 4390 29464 4392 29504
rect 4392 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4514 29504
rect 4558 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4680 29504
rect 4680 29464 4682 29504
rect 4390 29422 4514 29464
rect 4558 29422 4682 29464
rect 79990 29504 80114 29546
rect 80158 29504 80282 29546
rect 79990 29464 79992 29504
rect 79992 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80114 29504
rect 80158 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80280 29504
rect 80280 29464 80282 29504
rect 79990 29422 80114 29464
rect 80158 29422 80282 29464
rect 95110 29338 95234 29462
rect 95278 29338 95402 29462
rect 95110 29170 95234 29294
rect 95278 29170 95402 29294
rect 18270 28898 18394 29022
rect 18438 28898 18562 29022
rect 3150 28748 3274 28790
rect 3318 28748 3442 28790
rect 3150 28708 3152 28748
rect 3152 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3274 28748
rect 3318 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3440 28748
rect 3440 28708 3442 28748
rect 3150 28666 3274 28708
rect 3318 28666 3442 28708
rect 18270 28730 18394 28854
rect 18438 28730 18562 28854
rect 33390 28898 33514 29022
rect 33558 28898 33682 29022
rect 33390 28730 33514 28854
rect 33558 28730 33682 28854
rect 48510 28898 48634 29022
rect 48678 28898 48802 29022
rect 48510 28730 48634 28854
rect 48678 28730 48802 28854
rect 63630 28898 63754 29022
rect 63798 28898 63922 29022
rect 63630 28730 63754 28854
rect 63798 28730 63922 28854
rect 78750 28748 78874 28790
rect 78918 28748 79042 28790
rect 78750 28708 78752 28748
rect 78752 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78874 28748
rect 78918 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79040 28748
rect 79040 28708 79042 28748
rect 78750 28666 78874 28708
rect 78918 28666 79042 28708
rect 93870 28098 93994 28222
rect 94038 28098 94162 28222
rect 4390 27992 4514 28034
rect 4558 27992 4682 28034
rect 4390 27952 4392 27992
rect 4392 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4514 27992
rect 4558 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4680 27992
rect 4680 27952 4682 27992
rect 4390 27910 4514 27952
rect 4558 27910 4682 27952
rect 79990 27992 80114 28034
rect 80158 27992 80282 28034
rect 79990 27952 79992 27992
rect 79992 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80114 27992
rect 80158 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80280 27992
rect 80280 27952 80282 27992
rect 79990 27910 80114 27952
rect 80158 27910 80282 27952
rect 93870 27930 93994 28054
rect 94038 27930 94162 28054
rect 3150 27236 3274 27278
rect 3318 27236 3442 27278
rect 3150 27196 3152 27236
rect 3152 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3274 27236
rect 3318 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3440 27236
rect 3440 27196 3442 27236
rect 3150 27154 3274 27196
rect 3318 27154 3442 27196
rect 78750 27236 78874 27278
rect 78918 27236 79042 27278
rect 78750 27196 78752 27236
rect 78752 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78874 27236
rect 78918 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79040 27236
rect 79040 27196 79042 27236
rect 78750 27154 78874 27196
rect 78918 27154 79042 27196
rect 4390 26480 4514 26522
rect 4558 26480 4682 26522
rect 4390 26440 4392 26480
rect 4392 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4514 26480
rect 4558 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4680 26480
rect 4680 26440 4682 26480
rect 4390 26398 4514 26440
rect 4558 26398 4682 26440
rect 79990 26480 80114 26522
rect 80158 26480 80282 26522
rect 79990 26440 79992 26480
rect 79992 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80114 26480
rect 80158 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80280 26480
rect 80280 26440 80282 26480
rect 79990 26398 80114 26440
rect 80158 26398 80282 26440
rect 3150 25724 3274 25766
rect 3318 25724 3442 25766
rect 3150 25684 3152 25724
rect 3152 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3274 25724
rect 3318 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3440 25724
rect 3440 25684 3442 25724
rect 3150 25642 3274 25684
rect 3318 25642 3442 25684
rect 78750 25724 78874 25766
rect 78918 25724 79042 25766
rect 78750 25684 78752 25724
rect 78752 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78874 25724
rect 78918 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79040 25724
rect 79040 25684 79042 25724
rect 78750 25642 78874 25684
rect 78918 25642 79042 25684
rect 4390 24968 4514 25010
rect 4558 24968 4682 25010
rect 4390 24928 4392 24968
rect 4392 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4514 24968
rect 4558 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4680 24968
rect 4680 24928 4682 24968
rect 4390 24886 4514 24928
rect 4558 24886 4682 24928
rect 79990 24968 80114 25010
rect 80158 24968 80282 25010
rect 79990 24928 79992 24968
rect 79992 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80114 24968
rect 80158 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80280 24968
rect 80280 24928 80282 24968
rect 79990 24886 80114 24928
rect 80158 24886 80282 24928
rect 3150 24212 3274 24254
rect 3318 24212 3442 24254
rect 3150 24172 3152 24212
rect 3152 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3274 24212
rect 3318 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3440 24212
rect 3440 24172 3442 24212
rect 3150 24130 3274 24172
rect 3318 24130 3442 24172
rect 19510 24138 19634 24262
rect 19678 24138 19802 24262
rect 19510 23970 19634 24094
rect 19678 23970 19802 24094
rect 34630 24138 34754 24262
rect 34798 24138 34922 24262
rect 34630 23970 34754 24094
rect 34798 23970 34922 24094
rect 49750 24138 49874 24262
rect 49918 24138 50042 24262
rect 49750 23970 49874 24094
rect 49918 23970 50042 24094
rect 64870 24138 64994 24262
rect 65038 24138 65162 24262
rect 78750 24212 78874 24254
rect 78918 24212 79042 24254
rect 78750 24172 78752 24212
rect 78752 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78874 24212
rect 78918 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79040 24212
rect 79040 24172 79042 24212
rect 78750 24130 78874 24172
rect 78918 24130 79042 24172
rect 64870 23970 64994 24094
rect 65038 23970 65162 24094
rect 4390 23456 4514 23498
rect 4558 23456 4682 23498
rect 4390 23416 4392 23456
rect 4392 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4514 23456
rect 4558 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4680 23456
rect 4680 23416 4682 23456
rect 4390 23374 4514 23416
rect 4558 23374 4682 23416
rect 79990 23456 80114 23498
rect 80158 23456 80282 23498
rect 79990 23416 79992 23456
rect 79992 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80114 23456
rect 80158 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80280 23456
rect 80280 23416 80282 23456
rect 79990 23374 80114 23416
rect 80158 23374 80282 23416
rect 18270 22898 18394 23022
rect 18438 22898 18562 23022
rect 3150 22700 3274 22742
rect 3318 22700 3442 22742
rect 3150 22660 3152 22700
rect 3152 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3274 22700
rect 3318 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3440 22700
rect 3440 22660 3442 22700
rect 3150 22618 3274 22660
rect 3318 22618 3442 22660
rect 18270 22730 18394 22854
rect 18438 22730 18562 22854
rect 33390 22898 33514 23022
rect 33558 22898 33682 23022
rect 33390 22730 33514 22854
rect 33558 22730 33682 22854
rect 48510 22898 48634 23022
rect 48678 22898 48802 23022
rect 48510 22730 48634 22854
rect 48678 22730 48802 22854
rect 63630 22898 63754 23022
rect 63798 22898 63922 23022
rect 63630 22730 63754 22854
rect 63798 22730 63922 22854
rect 78750 22700 78874 22742
rect 78918 22700 79042 22742
rect 78750 22660 78752 22700
rect 78752 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78874 22700
rect 78918 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79040 22700
rect 79040 22660 79042 22700
rect 78750 22618 78874 22660
rect 78918 22618 79042 22660
rect 4390 21944 4514 21986
rect 4558 21944 4682 21986
rect 4390 21904 4392 21944
rect 4392 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4514 21944
rect 4558 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4680 21944
rect 4680 21904 4682 21944
rect 4390 21862 4514 21904
rect 4558 21862 4682 21904
rect 79990 21944 80114 21986
rect 80158 21944 80282 21986
rect 79990 21904 79992 21944
rect 79992 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80114 21944
rect 80158 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80280 21944
rect 80280 21904 80282 21944
rect 79990 21862 80114 21904
rect 80158 21862 80282 21904
rect 95110 21944 95234 21986
rect 95278 21944 95402 21986
rect 95110 21904 95112 21944
rect 95112 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95234 21944
rect 95278 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95400 21944
rect 95400 21904 95402 21944
rect 95110 21862 95234 21904
rect 95278 21862 95402 21904
rect 3150 21188 3274 21230
rect 3318 21188 3442 21230
rect 3150 21148 3152 21188
rect 3152 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3274 21188
rect 3318 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3440 21188
rect 3440 21148 3442 21188
rect 3150 21106 3274 21148
rect 3318 21106 3442 21148
rect 78750 21188 78874 21230
rect 78918 21188 79042 21230
rect 78750 21148 78752 21188
rect 78752 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78874 21188
rect 78918 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79040 21188
rect 79040 21148 79042 21188
rect 78750 21106 78874 21148
rect 78918 21106 79042 21148
rect 93870 21188 93994 21230
rect 94038 21188 94162 21230
rect 93870 21148 93872 21188
rect 93872 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93994 21188
rect 94038 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94160 21188
rect 94160 21148 94162 21188
rect 93870 21106 93994 21148
rect 94038 21106 94162 21148
rect 4390 20432 4514 20474
rect 4558 20432 4682 20474
rect 4390 20392 4392 20432
rect 4392 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4514 20432
rect 4558 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4680 20432
rect 4680 20392 4682 20432
rect 4390 20350 4514 20392
rect 4558 20350 4682 20392
rect 79990 20432 80114 20474
rect 80158 20432 80282 20474
rect 79990 20392 79992 20432
rect 79992 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80114 20432
rect 80158 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80280 20432
rect 80280 20392 80282 20432
rect 79990 20350 80114 20392
rect 80158 20350 80282 20392
rect 95110 20432 95234 20474
rect 95278 20432 95402 20474
rect 95110 20392 95112 20432
rect 95112 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95234 20432
rect 95278 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95400 20432
rect 95400 20392 95402 20432
rect 95110 20350 95234 20392
rect 95278 20350 95402 20392
rect 3150 19676 3274 19718
rect 3318 19676 3442 19718
rect 3150 19636 3152 19676
rect 3152 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3274 19676
rect 3318 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3440 19676
rect 3440 19636 3442 19676
rect 3150 19594 3274 19636
rect 3318 19594 3442 19636
rect 78750 19676 78874 19718
rect 78918 19676 79042 19718
rect 78750 19636 78752 19676
rect 78752 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78874 19676
rect 78918 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79040 19676
rect 79040 19636 79042 19676
rect 78750 19594 78874 19636
rect 78918 19594 79042 19636
rect 93870 19676 93994 19718
rect 94038 19676 94162 19718
rect 93870 19636 93872 19676
rect 93872 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93994 19676
rect 94038 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94160 19676
rect 94160 19636 94162 19676
rect 93870 19594 93994 19636
rect 94038 19594 94162 19636
rect 4390 18920 4514 18962
rect 4558 18920 4682 18962
rect 4390 18880 4392 18920
rect 4392 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4514 18920
rect 4558 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4680 18920
rect 4680 18880 4682 18920
rect 4390 18838 4514 18880
rect 4558 18838 4682 18880
rect 79990 18920 80114 18962
rect 80158 18920 80282 18962
rect 79990 18880 79992 18920
rect 79992 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80114 18920
rect 80158 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80280 18920
rect 80280 18880 80282 18920
rect 79990 18838 80114 18880
rect 80158 18838 80282 18880
rect 3150 18164 3274 18206
rect 3318 18164 3442 18206
rect 3150 18124 3152 18164
rect 3152 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3274 18164
rect 3318 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3440 18164
rect 3440 18124 3442 18164
rect 3150 18082 3274 18124
rect 3318 18082 3442 18124
rect 19510 18138 19634 18262
rect 19678 18138 19802 18262
rect 19510 17970 19634 18094
rect 19678 17970 19802 18094
rect 34630 18138 34754 18262
rect 34798 18138 34922 18262
rect 34630 17970 34754 18094
rect 34798 17970 34922 18094
rect 49750 18138 49874 18262
rect 49918 18138 50042 18262
rect 49750 17970 49874 18094
rect 49918 17970 50042 18094
rect 64870 18138 64994 18262
rect 65038 18138 65162 18262
rect 64870 17970 64994 18094
rect 65038 17970 65162 18094
rect 78750 18164 78874 18206
rect 78918 18164 79042 18206
rect 78750 18124 78752 18164
rect 78752 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78874 18164
rect 78918 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79040 18164
rect 79040 18124 79042 18164
rect 78750 18082 78874 18124
rect 78918 18082 79042 18124
rect 4390 17408 4514 17450
rect 4558 17408 4682 17450
rect 4390 17368 4392 17408
rect 4392 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4514 17408
rect 4558 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4680 17408
rect 4680 17368 4682 17408
rect 4390 17326 4514 17368
rect 4558 17326 4682 17368
rect 79990 17408 80114 17450
rect 80158 17408 80282 17450
rect 79990 17368 79992 17408
rect 79992 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80114 17408
rect 80158 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80280 17408
rect 80280 17368 80282 17408
rect 79990 17326 80114 17368
rect 80158 17326 80282 17368
rect 18270 16898 18394 17022
rect 18438 16898 18562 17022
rect 18270 16730 18394 16854
rect 18438 16730 18562 16854
rect 3150 16652 3274 16694
rect 3318 16652 3442 16694
rect 33390 16898 33514 17022
rect 33558 16898 33682 17022
rect 33390 16730 33514 16854
rect 33558 16730 33682 16854
rect 48510 16898 48634 17022
rect 48678 16898 48802 17022
rect 48510 16730 48634 16854
rect 48678 16730 48802 16854
rect 63630 16898 63754 17022
rect 63798 16898 63922 17022
rect 63630 16730 63754 16854
rect 63798 16730 63922 16854
rect 3150 16612 3152 16652
rect 3152 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3274 16652
rect 3318 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3440 16652
rect 3440 16612 3442 16652
rect 3150 16570 3274 16612
rect 3318 16570 3442 16612
rect 78750 16652 78874 16694
rect 78918 16652 79042 16694
rect 78750 16612 78752 16652
rect 78752 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78874 16652
rect 78918 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79040 16652
rect 79040 16612 79042 16652
rect 78750 16570 78874 16612
rect 78918 16570 79042 16612
rect 4390 15896 4514 15938
rect 4558 15896 4682 15938
rect 4390 15856 4392 15896
rect 4392 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4514 15896
rect 4558 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4680 15896
rect 4680 15856 4682 15896
rect 4390 15814 4514 15856
rect 4558 15814 4682 15856
rect 79990 15896 80114 15938
rect 80158 15896 80282 15938
rect 79990 15856 79992 15896
rect 79992 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80114 15896
rect 80158 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80280 15896
rect 80280 15856 80282 15896
rect 79990 15814 80114 15856
rect 80158 15814 80282 15856
rect 3150 15140 3274 15182
rect 3318 15140 3442 15182
rect 3150 15100 3152 15140
rect 3152 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3274 15140
rect 3318 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3440 15140
rect 3440 15100 3442 15140
rect 3150 15058 3274 15100
rect 3318 15058 3442 15100
rect 78750 15140 78874 15182
rect 78918 15140 79042 15182
rect 78750 15100 78752 15140
rect 78752 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78874 15140
rect 78918 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79040 15140
rect 79040 15100 79042 15140
rect 78750 15058 78874 15100
rect 78918 15058 79042 15100
rect 4390 14384 4514 14426
rect 4558 14384 4682 14426
rect 4390 14344 4392 14384
rect 4392 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4514 14384
rect 4558 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4680 14384
rect 4680 14344 4682 14384
rect 4390 14302 4514 14344
rect 4558 14302 4682 14344
rect 79990 14384 80114 14426
rect 80158 14384 80282 14426
rect 79990 14344 79992 14384
rect 79992 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80114 14384
rect 80158 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80280 14384
rect 80280 14344 80282 14384
rect 79990 14302 80114 14344
rect 80158 14302 80282 14344
rect 3150 13628 3274 13670
rect 3318 13628 3442 13670
rect 3150 13588 3152 13628
rect 3152 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3274 13628
rect 3318 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3440 13628
rect 3440 13588 3442 13628
rect 3150 13546 3274 13588
rect 3318 13546 3442 13588
rect 78750 13628 78874 13670
rect 78918 13628 79042 13670
rect 78750 13588 78752 13628
rect 78752 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78874 13628
rect 78918 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79040 13628
rect 79040 13588 79042 13628
rect 78750 13546 78874 13588
rect 78918 13546 79042 13588
rect 4390 12872 4514 12914
rect 4558 12872 4682 12914
rect 4390 12832 4392 12872
rect 4392 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4514 12872
rect 4558 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4680 12872
rect 4680 12832 4682 12872
rect 4390 12790 4514 12832
rect 4558 12790 4682 12832
rect 79990 12872 80114 12914
rect 80158 12872 80282 12914
rect 79990 12832 79992 12872
rect 79992 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80114 12872
rect 80158 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80280 12872
rect 80280 12832 80282 12872
rect 79990 12790 80114 12832
rect 80158 12790 80282 12832
rect 3150 12116 3274 12158
rect 3318 12116 3442 12158
rect 3150 12076 3152 12116
rect 3152 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3274 12116
rect 3318 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3440 12116
rect 3440 12076 3442 12116
rect 3150 12034 3274 12076
rect 3318 12034 3442 12076
rect 19510 12138 19634 12262
rect 19678 12138 19802 12262
rect 19510 11970 19634 12094
rect 19678 11970 19802 12094
rect 34630 12138 34754 12262
rect 34798 12138 34922 12262
rect 34630 11970 34754 12094
rect 34798 11970 34922 12094
rect 49750 12138 49874 12262
rect 49918 12138 50042 12262
rect 49750 11970 49874 12094
rect 49918 11970 50042 12094
rect 64870 12138 64994 12262
rect 65038 12138 65162 12262
rect 64870 11970 64994 12094
rect 65038 11970 65162 12094
rect 78750 12116 78874 12158
rect 78918 12116 79042 12158
rect 78750 12076 78752 12116
rect 78752 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78874 12116
rect 78918 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79040 12116
rect 79040 12076 79042 12116
rect 78750 12034 78874 12076
rect 78918 12034 79042 12076
rect 95110 12138 95234 12262
rect 95278 12138 95402 12262
rect 95110 11970 95234 12094
rect 95278 11970 95402 12094
rect 4390 11360 4514 11402
rect 4558 11360 4682 11402
rect 4390 11320 4392 11360
rect 4392 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4514 11360
rect 4558 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4680 11360
rect 4680 11320 4682 11360
rect 4390 11278 4514 11320
rect 4558 11278 4682 11320
rect 79990 11360 80114 11402
rect 80158 11360 80282 11402
rect 79990 11320 79992 11360
rect 79992 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80114 11360
rect 80158 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80280 11360
rect 80280 11320 80282 11360
rect 79990 11278 80114 11320
rect 80158 11278 80282 11320
rect 18270 10898 18394 11022
rect 18438 10898 18562 11022
rect 18270 10730 18394 10854
rect 18438 10730 18562 10854
rect 33390 10898 33514 11022
rect 33558 10898 33682 11022
rect 33390 10730 33514 10854
rect 33558 10730 33682 10854
rect 48510 10898 48634 11022
rect 48678 10898 48802 11022
rect 48510 10730 48634 10854
rect 48678 10730 48802 10854
rect 63630 10898 63754 11022
rect 63798 10898 63922 11022
rect 63630 10730 63754 10854
rect 63798 10730 63922 10854
rect 93870 10898 93994 11022
rect 94038 10898 94162 11022
rect 93870 10730 93994 10854
rect 94038 10730 94162 10854
rect 3150 10604 3274 10646
rect 3318 10604 3442 10646
rect 3150 10564 3152 10604
rect 3152 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3274 10604
rect 3318 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3440 10604
rect 3440 10564 3442 10604
rect 3150 10522 3274 10564
rect 3318 10522 3442 10564
rect 78750 10604 78874 10646
rect 78918 10604 79042 10646
rect 78750 10564 78752 10604
rect 78752 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78874 10604
rect 78918 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79040 10604
rect 79040 10564 79042 10604
rect 78750 10522 78874 10564
rect 78918 10522 79042 10564
rect 4390 9848 4514 9890
rect 4558 9848 4682 9890
rect 4390 9808 4392 9848
rect 4392 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4514 9848
rect 4558 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4680 9848
rect 4680 9808 4682 9848
rect 4390 9766 4514 9808
rect 4558 9766 4682 9808
rect 79990 9848 80114 9890
rect 80158 9848 80282 9890
rect 79990 9808 79992 9848
rect 79992 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80114 9848
rect 80158 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80280 9848
rect 80280 9808 80282 9848
rect 79990 9766 80114 9808
rect 80158 9766 80282 9808
rect 3150 9092 3274 9134
rect 3318 9092 3442 9134
rect 3150 9052 3152 9092
rect 3152 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3274 9092
rect 3318 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3440 9092
rect 3440 9052 3442 9092
rect 3150 9010 3274 9052
rect 3318 9010 3442 9052
rect 78750 9092 78874 9134
rect 78918 9092 79042 9134
rect 78750 9052 78752 9092
rect 78752 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78874 9092
rect 78918 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79040 9092
rect 79040 9052 79042 9092
rect 78750 9010 78874 9052
rect 78918 9010 79042 9052
rect 4390 8336 4514 8378
rect 4558 8336 4682 8378
rect 4390 8296 4392 8336
rect 4392 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4514 8336
rect 4558 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4680 8336
rect 4680 8296 4682 8336
rect 4390 8254 4514 8296
rect 4558 8254 4682 8296
rect 79990 8336 80114 8378
rect 80158 8336 80282 8378
rect 79990 8296 79992 8336
rect 79992 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80114 8336
rect 80158 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80280 8336
rect 80280 8296 80282 8336
rect 79990 8254 80114 8296
rect 80158 8254 80282 8296
rect 67298 7750 67422 7874
rect 3150 7580 3274 7622
rect 3318 7580 3442 7622
rect 3150 7540 3152 7580
rect 3152 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3274 7580
rect 3318 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3440 7580
rect 3440 7540 3442 7580
rect 3150 7498 3274 7540
rect 3318 7498 3442 7540
rect 78750 7580 78874 7622
rect 78918 7580 79042 7622
rect 78750 7540 78752 7580
rect 78752 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78874 7580
rect 78918 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79040 7580
rect 79040 7540 79042 7580
rect 78750 7498 78874 7540
rect 78918 7498 79042 7540
rect 4390 6824 4514 6866
rect 4558 6824 4682 6866
rect 4390 6784 4392 6824
rect 4392 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4514 6824
rect 4558 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4680 6824
rect 4680 6784 4682 6824
rect 4390 6742 4514 6784
rect 4558 6742 4682 6784
rect 79990 6824 80114 6866
rect 80158 6824 80282 6866
rect 79990 6784 79992 6824
rect 79992 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80114 6824
rect 80158 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80280 6824
rect 80280 6784 80282 6824
rect 79990 6742 80114 6784
rect 80158 6742 80282 6784
rect 95110 6138 95234 6262
rect 95278 6138 95402 6262
rect 3150 6068 3274 6110
rect 3318 6068 3442 6110
rect 3150 6028 3152 6068
rect 3152 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3274 6068
rect 3318 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3440 6068
rect 3440 6028 3442 6068
rect 3150 5986 3274 6028
rect 3318 5986 3442 6028
rect 78750 6068 78874 6110
rect 78918 6068 79042 6110
rect 78750 6028 78752 6068
rect 78752 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78874 6068
rect 78918 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79040 6068
rect 79040 6028 79042 6068
rect 78750 5986 78874 6028
rect 78918 5986 79042 6028
rect 95110 5970 95234 6094
rect 95278 5970 95402 6094
rect 66386 5734 66510 5858
rect 4390 5312 4514 5354
rect 4558 5312 4682 5354
rect 4390 5272 4392 5312
rect 4392 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4514 5312
rect 4558 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4680 5312
rect 4680 5272 4682 5312
rect 4390 5230 4514 5272
rect 4558 5230 4682 5272
rect 19510 5312 19634 5354
rect 19678 5312 19802 5354
rect 19510 5272 19512 5312
rect 19512 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19634 5312
rect 19678 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19800 5312
rect 19800 5272 19802 5312
rect 19510 5230 19634 5272
rect 19678 5230 19802 5272
rect 34630 5312 34754 5354
rect 34798 5312 34922 5354
rect 34630 5272 34632 5312
rect 34632 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34754 5312
rect 34798 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34920 5312
rect 34920 5272 34922 5312
rect 34630 5230 34754 5272
rect 34798 5230 34922 5272
rect 49750 5312 49874 5354
rect 49918 5312 50042 5354
rect 49750 5272 49752 5312
rect 49752 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49874 5312
rect 49918 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50040 5312
rect 50040 5272 50042 5312
rect 49750 5230 49874 5272
rect 49918 5230 50042 5272
rect 64870 5312 64994 5354
rect 65038 5312 65162 5354
rect 64870 5272 64872 5312
rect 64872 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64994 5312
rect 65038 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65160 5312
rect 65160 5272 65162 5312
rect 64870 5230 64994 5272
rect 65038 5230 65162 5272
rect 79990 5312 80114 5354
rect 80158 5312 80282 5354
rect 79990 5272 79992 5312
rect 79992 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80114 5312
rect 80158 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80280 5312
rect 80280 5272 80282 5312
rect 79990 5230 80114 5272
rect 80158 5230 80282 5272
rect 93870 4898 93994 5022
rect 94038 4898 94162 5022
rect 93870 4730 93994 4854
rect 94038 4730 94162 4854
rect 3150 4556 3274 4598
rect 3318 4556 3442 4598
rect 3150 4516 3152 4556
rect 3152 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3274 4556
rect 3318 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3440 4556
rect 3440 4516 3442 4556
rect 3150 4474 3274 4516
rect 3318 4474 3442 4516
rect 18270 4556 18394 4598
rect 18438 4556 18562 4598
rect 18270 4516 18272 4556
rect 18272 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18394 4556
rect 18438 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18560 4556
rect 18560 4516 18562 4556
rect 18270 4474 18394 4516
rect 18438 4474 18562 4516
rect 33390 4556 33514 4598
rect 33558 4556 33682 4598
rect 33390 4516 33392 4556
rect 33392 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33514 4556
rect 33558 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33680 4556
rect 33680 4516 33682 4556
rect 33390 4474 33514 4516
rect 33558 4474 33682 4516
rect 48510 4556 48634 4598
rect 48678 4556 48802 4598
rect 48510 4516 48512 4556
rect 48512 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48634 4556
rect 48678 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48800 4556
rect 48800 4516 48802 4556
rect 48510 4474 48634 4516
rect 48678 4474 48802 4516
rect 63630 4556 63754 4598
rect 63798 4556 63922 4598
rect 63630 4516 63632 4556
rect 63632 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63754 4556
rect 63798 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63920 4556
rect 63920 4516 63922 4556
rect 63630 4474 63754 4516
rect 63798 4474 63922 4516
rect 78750 4556 78874 4598
rect 78918 4556 79042 4598
rect 78750 4516 78752 4556
rect 78752 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78874 4556
rect 78918 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79040 4556
rect 79040 4516 79042 4556
rect 78750 4474 78874 4516
rect 78918 4474 79042 4516
rect 4390 3800 4514 3842
rect 4558 3800 4682 3842
rect 4390 3760 4392 3800
rect 4392 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4514 3800
rect 4558 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4680 3800
rect 4680 3760 4682 3800
rect 4390 3718 4514 3760
rect 4558 3718 4682 3760
rect 19510 3800 19634 3842
rect 19678 3800 19802 3842
rect 19510 3760 19512 3800
rect 19512 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19634 3800
rect 19678 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19800 3800
rect 19800 3760 19802 3800
rect 19510 3718 19634 3760
rect 19678 3718 19802 3760
rect 34630 3800 34754 3842
rect 34798 3800 34922 3842
rect 34630 3760 34632 3800
rect 34632 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34754 3800
rect 34798 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34920 3800
rect 34920 3760 34922 3800
rect 34630 3718 34754 3760
rect 34798 3718 34922 3760
rect 49750 3800 49874 3842
rect 49918 3800 50042 3842
rect 49750 3760 49752 3800
rect 49752 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49874 3800
rect 49918 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50040 3800
rect 50040 3760 50042 3800
rect 49750 3718 49874 3760
rect 49918 3718 50042 3760
rect 64870 3800 64994 3842
rect 65038 3800 65162 3842
rect 64870 3760 64872 3800
rect 64872 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64994 3800
rect 65038 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65160 3800
rect 65160 3760 65162 3800
rect 64870 3718 64994 3760
rect 65038 3718 65162 3760
rect 79990 3800 80114 3842
rect 80158 3800 80282 3842
rect 79990 3760 79992 3800
rect 79992 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80114 3800
rect 80158 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80280 3800
rect 80280 3760 80282 3800
rect 79990 3718 80114 3760
rect 80158 3718 80282 3760
rect 3150 3044 3274 3086
rect 3318 3044 3442 3086
rect 3150 3004 3152 3044
rect 3152 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3274 3044
rect 3318 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3440 3044
rect 3440 3004 3442 3044
rect 3150 2962 3274 3004
rect 3318 2962 3442 3004
rect 18270 3044 18394 3086
rect 18438 3044 18562 3086
rect 18270 3004 18272 3044
rect 18272 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18394 3044
rect 18438 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18560 3044
rect 18560 3004 18562 3044
rect 18270 2962 18394 3004
rect 18438 2962 18562 3004
rect 33390 3044 33514 3086
rect 33558 3044 33682 3086
rect 33390 3004 33392 3044
rect 33392 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33514 3044
rect 33558 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33680 3044
rect 33680 3004 33682 3044
rect 33390 2962 33514 3004
rect 33558 2962 33682 3004
rect 48510 3044 48634 3086
rect 48678 3044 48802 3086
rect 48510 3004 48512 3044
rect 48512 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48634 3044
rect 48678 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48800 3044
rect 48800 3004 48802 3044
rect 48510 2962 48634 3004
rect 48678 2962 48802 3004
rect 63630 3044 63754 3086
rect 63798 3044 63922 3086
rect 63630 3004 63632 3044
rect 63632 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63754 3044
rect 63798 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63920 3044
rect 63920 3004 63922 3044
rect 63630 2962 63754 3004
rect 63798 2962 63922 3004
rect 78750 3044 78874 3086
rect 78918 3044 79042 3086
rect 78750 3004 78752 3044
rect 78752 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78874 3044
rect 78918 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79040 3044
rect 79040 3004 79042 3044
rect 78750 2962 78874 3004
rect 78918 2962 79042 3004
rect 4390 2288 4514 2330
rect 4558 2288 4682 2330
rect 4390 2248 4392 2288
rect 4392 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4514 2288
rect 4558 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4680 2288
rect 4680 2248 4682 2288
rect 4390 2206 4514 2248
rect 4558 2206 4682 2248
rect 19510 2288 19634 2330
rect 19678 2288 19802 2330
rect 19510 2248 19512 2288
rect 19512 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19634 2288
rect 19678 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19800 2288
rect 19800 2248 19802 2288
rect 19510 2206 19634 2248
rect 19678 2206 19802 2248
rect 34630 2288 34754 2330
rect 34798 2288 34922 2330
rect 34630 2248 34632 2288
rect 34632 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34754 2288
rect 34798 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34920 2288
rect 34920 2248 34922 2288
rect 34630 2206 34754 2248
rect 34798 2206 34922 2248
rect 49750 2288 49874 2330
rect 49918 2288 50042 2330
rect 49750 2248 49752 2288
rect 49752 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49874 2288
rect 49918 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50040 2288
rect 50040 2248 50042 2288
rect 49750 2206 49874 2248
rect 49918 2206 50042 2248
rect 64870 2288 64994 2330
rect 65038 2288 65162 2330
rect 64870 2248 64872 2288
rect 64872 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64994 2288
rect 65038 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65160 2288
rect 65160 2248 65162 2288
rect 64870 2206 64994 2248
rect 65038 2206 65162 2248
rect 79990 2288 80114 2330
rect 80158 2288 80282 2330
rect 79990 2248 79992 2288
rect 79992 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80114 2288
rect 80158 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80280 2288
rect 80280 2248 80282 2288
rect 79990 2206 80114 2248
rect 80158 2206 80282 2248
rect 3150 1532 3274 1574
rect 3318 1532 3442 1574
rect 3150 1492 3152 1532
rect 3152 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3274 1532
rect 3318 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3440 1532
rect 3440 1492 3442 1532
rect 3150 1450 3274 1492
rect 3318 1450 3442 1492
rect 18270 1532 18394 1574
rect 18438 1532 18562 1574
rect 18270 1492 18272 1532
rect 18272 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18394 1532
rect 18438 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18560 1532
rect 18560 1492 18562 1532
rect 18270 1450 18394 1492
rect 18438 1450 18562 1492
rect 33390 1532 33514 1574
rect 33558 1532 33682 1574
rect 33390 1492 33392 1532
rect 33392 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33514 1532
rect 33558 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33680 1532
rect 33680 1492 33682 1532
rect 33390 1450 33514 1492
rect 33558 1450 33682 1492
rect 48510 1532 48634 1574
rect 48678 1532 48802 1574
rect 48510 1492 48512 1532
rect 48512 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48634 1532
rect 48678 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48800 1532
rect 48800 1492 48802 1532
rect 48510 1450 48634 1492
rect 48678 1450 48802 1492
rect 63630 1532 63754 1574
rect 63798 1532 63922 1574
rect 63630 1492 63632 1532
rect 63632 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63754 1532
rect 63798 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63920 1532
rect 63920 1492 63922 1532
rect 63630 1450 63754 1492
rect 63798 1450 63922 1492
rect 78750 1532 78874 1574
rect 78918 1532 79042 1574
rect 78750 1492 78752 1532
rect 78752 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78874 1532
rect 78918 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79040 1532
rect 79040 1492 79042 1532
rect 78750 1450 78874 1492
rect 78918 1450 79042 1492
rect 4390 776 4514 818
rect 4558 776 4682 818
rect 4390 736 4392 776
rect 4392 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4514 776
rect 4558 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4680 776
rect 4680 736 4682 776
rect 4390 694 4514 736
rect 4558 694 4682 736
rect 19510 776 19634 818
rect 19678 776 19802 818
rect 19510 736 19512 776
rect 19512 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19634 776
rect 19678 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19800 776
rect 19800 736 19802 776
rect 19510 694 19634 736
rect 19678 694 19802 736
rect 34630 776 34754 818
rect 34798 776 34922 818
rect 34630 736 34632 776
rect 34632 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34754 776
rect 34798 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34920 776
rect 34920 736 34922 776
rect 34630 694 34754 736
rect 34798 694 34922 736
rect 49750 776 49874 818
rect 49918 776 50042 818
rect 49750 736 49752 776
rect 49752 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49874 776
rect 49918 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50040 776
rect 50040 736 50042 776
rect 49750 694 49874 736
rect 49918 694 50042 736
rect 64870 776 64994 818
rect 65038 776 65162 818
rect 64870 736 64872 776
rect 64872 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64994 776
rect 65038 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65160 776
rect 65160 736 65162 776
rect 64870 694 64994 736
rect 65038 694 65162 736
rect 79990 776 80114 818
rect 80158 776 80282 818
rect 79990 736 79992 776
rect 79992 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80114 776
rect 80158 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80280 776
rect 80280 736 80282 776
rect 79990 694 80114 736
rect 80158 694 80282 736
<< metal6 >>
rect 4316 38618 4756 38682
rect 3076 37862 3516 38600
rect 3076 37738 3150 37862
rect 3274 37738 3318 37862
rect 3442 37738 3516 37862
rect 3076 36350 3516 37738
rect 3076 36226 3150 36350
rect 3274 36226 3318 36350
rect 3442 36226 3516 36350
rect 3076 34838 3516 36226
rect 3076 34714 3150 34838
rect 3274 34714 3318 34838
rect 3442 34714 3516 34838
rect 3076 33326 3516 34714
rect 3076 33202 3150 33326
rect 3274 33202 3318 33326
rect 3442 33202 3516 33326
rect 3076 31814 3516 33202
rect 3076 31690 3150 31814
rect 3274 31690 3318 31814
rect 3442 31690 3516 31814
rect 3076 30302 3516 31690
rect 3076 30178 3150 30302
rect 3274 30178 3318 30302
rect 3442 30178 3516 30302
rect 3076 28790 3516 30178
rect 3076 28666 3150 28790
rect 3274 28666 3318 28790
rect 3442 28666 3516 28790
rect 3076 27278 3516 28666
rect 3076 27154 3150 27278
rect 3274 27154 3318 27278
rect 3442 27154 3516 27278
rect 3076 25766 3516 27154
rect 3076 25642 3150 25766
rect 3274 25642 3318 25766
rect 3442 25642 3516 25766
rect 3076 24254 3516 25642
rect 3076 24130 3150 24254
rect 3274 24130 3318 24254
rect 3442 24130 3516 24254
rect 3076 22742 3516 24130
rect 3076 22618 3150 22742
rect 3274 22618 3318 22742
rect 3442 22618 3516 22742
rect 3076 21230 3516 22618
rect 3076 21106 3150 21230
rect 3274 21106 3318 21230
rect 3442 21106 3516 21230
rect 3076 19718 3516 21106
rect 3076 19594 3150 19718
rect 3274 19594 3318 19718
rect 3442 19594 3516 19718
rect 3076 18206 3516 19594
rect 3076 18082 3150 18206
rect 3274 18082 3318 18206
rect 3442 18082 3516 18206
rect 3076 16694 3516 18082
rect 3076 16570 3150 16694
rect 3274 16570 3318 16694
rect 3442 16570 3516 16694
rect 3076 15182 3516 16570
rect 3076 15058 3150 15182
rect 3274 15058 3318 15182
rect 3442 15058 3516 15182
rect 3076 13670 3516 15058
rect 3076 13546 3150 13670
rect 3274 13546 3318 13670
rect 3442 13546 3516 13670
rect 3076 12158 3516 13546
rect 3076 12034 3150 12158
rect 3274 12034 3318 12158
rect 3442 12034 3516 12158
rect 3076 10646 3516 12034
rect 3076 10522 3150 10646
rect 3274 10522 3318 10646
rect 3442 10522 3516 10646
rect 3076 9134 3516 10522
rect 3076 9010 3150 9134
rect 3274 9010 3318 9134
rect 3442 9010 3516 9134
rect 3076 7622 3516 9010
rect 3076 7498 3150 7622
rect 3274 7498 3318 7622
rect 3442 7498 3516 7622
rect 3076 6110 3516 7498
rect 3076 5986 3150 6110
rect 3274 5986 3318 6110
rect 3442 5986 3516 6110
rect 3076 4598 3516 5986
rect 3076 4474 3150 4598
rect 3274 4474 3318 4598
rect 3442 4474 3516 4598
rect 3076 3086 3516 4474
rect 3076 2962 3150 3086
rect 3274 2962 3318 3086
rect 3442 2962 3516 3086
rect 3076 1574 3516 2962
rect 3076 1450 3150 1574
rect 3274 1450 3318 1574
rect 3442 1450 3516 1574
rect 3076 712 3516 1450
rect 4316 38494 4390 38618
rect 4514 38494 4558 38618
rect 4682 38494 4756 38618
rect 19436 38618 19876 38682
rect 4316 37106 4756 38494
rect 4316 36982 4390 37106
rect 4514 36982 4558 37106
rect 4682 36982 4756 37106
rect 4316 35594 4756 36982
rect 4316 35470 4390 35594
rect 4514 35470 4558 35594
rect 4682 35470 4756 35594
rect 4316 34082 4756 35470
rect 4316 33958 4390 34082
rect 4514 33958 4558 34082
rect 4682 33958 4756 34082
rect 4316 32570 4756 33958
rect 4316 32446 4390 32570
rect 4514 32446 4558 32570
rect 4682 32446 4756 32570
rect 4316 31058 4756 32446
rect 4316 30934 4390 31058
rect 4514 30934 4558 31058
rect 4682 30934 4756 31058
rect 4316 29546 4756 30934
rect 4316 29422 4390 29546
rect 4514 29422 4558 29546
rect 4682 29422 4756 29546
rect 4316 28034 4756 29422
rect 4316 27910 4390 28034
rect 4514 27910 4558 28034
rect 4682 27910 4756 28034
rect 4316 26522 4756 27910
rect 4316 26398 4390 26522
rect 4514 26398 4558 26522
rect 4682 26398 4756 26522
rect 4316 25010 4756 26398
rect 4316 24886 4390 25010
rect 4514 24886 4558 25010
rect 4682 24886 4756 25010
rect 4316 23498 4756 24886
rect 4316 23374 4390 23498
rect 4514 23374 4558 23498
rect 4682 23374 4756 23498
rect 4316 21986 4756 23374
rect 4316 21862 4390 21986
rect 4514 21862 4558 21986
rect 4682 21862 4756 21986
rect 4316 20474 4756 21862
rect 4316 20350 4390 20474
rect 4514 20350 4558 20474
rect 4682 20350 4756 20474
rect 4316 18962 4756 20350
rect 4316 18838 4390 18962
rect 4514 18838 4558 18962
rect 4682 18838 4756 18962
rect 4316 17450 4756 18838
rect 4316 17326 4390 17450
rect 4514 17326 4558 17450
rect 4682 17326 4756 17450
rect 4316 15938 4756 17326
rect 4316 15814 4390 15938
rect 4514 15814 4558 15938
rect 4682 15814 4756 15938
rect 4316 14426 4756 15814
rect 4316 14302 4390 14426
rect 4514 14302 4558 14426
rect 4682 14302 4756 14426
rect 4316 12914 4756 14302
rect 4316 12790 4390 12914
rect 4514 12790 4558 12914
rect 4682 12790 4756 12914
rect 4316 11402 4756 12790
rect 4316 11278 4390 11402
rect 4514 11278 4558 11402
rect 4682 11278 4756 11402
rect 4316 9890 4756 11278
rect 4316 9766 4390 9890
rect 4514 9766 4558 9890
rect 4682 9766 4756 9890
rect 4316 8378 4756 9766
rect 4316 8254 4390 8378
rect 4514 8254 4558 8378
rect 4682 8254 4756 8378
rect 4316 6866 4756 8254
rect 4316 6742 4390 6866
rect 4514 6742 4558 6866
rect 4682 6742 4756 6866
rect 4316 5354 4756 6742
rect 4316 5230 4390 5354
rect 4514 5230 4558 5354
rect 4682 5230 4756 5354
rect 4316 3842 4756 5230
rect 4316 3718 4390 3842
rect 4514 3718 4558 3842
rect 4682 3718 4756 3842
rect 4316 2330 4756 3718
rect 4316 2206 4390 2330
rect 4514 2206 4558 2330
rect 4682 2206 4756 2330
rect 4316 818 4756 2206
rect 4316 694 4390 818
rect 4514 694 4558 818
rect 4682 694 4756 818
rect 18196 37862 18636 38600
rect 18196 37738 18270 37862
rect 18394 37738 18438 37862
rect 18562 37738 18636 37862
rect 18196 36350 18636 37738
rect 18196 36226 18270 36350
rect 18394 36226 18438 36350
rect 18562 36226 18636 36350
rect 18196 34838 18636 36226
rect 18196 34714 18270 34838
rect 18394 34714 18438 34838
rect 18562 34714 18636 34838
rect 18196 29022 18636 34714
rect 18196 28898 18270 29022
rect 18394 28898 18438 29022
rect 18562 28898 18636 29022
rect 18196 28854 18636 28898
rect 18196 28730 18270 28854
rect 18394 28730 18438 28854
rect 18562 28730 18636 28854
rect 18196 23022 18636 28730
rect 18196 22898 18270 23022
rect 18394 22898 18438 23022
rect 18562 22898 18636 23022
rect 18196 22854 18636 22898
rect 18196 22730 18270 22854
rect 18394 22730 18438 22854
rect 18562 22730 18636 22854
rect 18196 17022 18636 22730
rect 18196 16898 18270 17022
rect 18394 16898 18438 17022
rect 18562 16898 18636 17022
rect 18196 16854 18636 16898
rect 18196 16730 18270 16854
rect 18394 16730 18438 16854
rect 18562 16730 18636 16854
rect 18196 11022 18636 16730
rect 18196 10898 18270 11022
rect 18394 10898 18438 11022
rect 18562 10898 18636 11022
rect 18196 10854 18636 10898
rect 18196 10730 18270 10854
rect 18394 10730 18438 10854
rect 18562 10730 18636 10854
rect 18196 4598 18636 10730
rect 18196 4474 18270 4598
rect 18394 4474 18438 4598
rect 18562 4474 18636 4598
rect 18196 3086 18636 4474
rect 18196 2962 18270 3086
rect 18394 2962 18438 3086
rect 18562 2962 18636 3086
rect 18196 1574 18636 2962
rect 18196 1450 18270 1574
rect 18394 1450 18438 1574
rect 18562 1450 18636 1574
rect 18196 712 18636 1450
rect 19436 38494 19510 38618
rect 19634 38494 19678 38618
rect 19802 38494 19876 38618
rect 34556 38618 34996 38682
rect 19436 37106 19876 38494
rect 19436 36982 19510 37106
rect 19634 36982 19678 37106
rect 19802 36982 19876 37106
rect 19436 35594 19876 36982
rect 19436 35470 19510 35594
rect 19634 35470 19678 35594
rect 19802 35470 19876 35594
rect 19436 34082 19876 35470
rect 19436 33958 19510 34082
rect 19634 33958 19678 34082
rect 19802 33958 19876 34082
rect 19436 24262 19876 33958
rect 19436 24138 19510 24262
rect 19634 24138 19678 24262
rect 19802 24138 19876 24262
rect 19436 24094 19876 24138
rect 19436 23970 19510 24094
rect 19634 23970 19678 24094
rect 19802 23970 19876 24094
rect 19436 18262 19876 23970
rect 19436 18138 19510 18262
rect 19634 18138 19678 18262
rect 19802 18138 19876 18262
rect 19436 18094 19876 18138
rect 19436 17970 19510 18094
rect 19634 17970 19678 18094
rect 19802 17970 19876 18094
rect 19436 12262 19876 17970
rect 19436 12138 19510 12262
rect 19634 12138 19678 12262
rect 19802 12138 19876 12262
rect 19436 12094 19876 12138
rect 19436 11970 19510 12094
rect 19634 11970 19678 12094
rect 19802 11970 19876 12094
rect 19436 5354 19876 11970
rect 19436 5230 19510 5354
rect 19634 5230 19678 5354
rect 19802 5230 19876 5354
rect 19436 3842 19876 5230
rect 19436 3718 19510 3842
rect 19634 3718 19678 3842
rect 19802 3718 19876 3842
rect 19436 2330 19876 3718
rect 19436 2206 19510 2330
rect 19634 2206 19678 2330
rect 19802 2206 19876 2330
rect 19436 818 19876 2206
rect 4316 630 4756 694
rect 19436 694 19510 818
rect 19634 694 19678 818
rect 19802 694 19876 818
rect 33316 37862 33756 38600
rect 33316 37738 33390 37862
rect 33514 37738 33558 37862
rect 33682 37738 33756 37862
rect 33316 36350 33756 37738
rect 33316 36226 33390 36350
rect 33514 36226 33558 36350
rect 33682 36226 33756 36350
rect 33316 34838 33756 36226
rect 33316 34714 33390 34838
rect 33514 34714 33558 34838
rect 33682 34714 33756 34838
rect 33316 29022 33756 34714
rect 33316 28898 33390 29022
rect 33514 28898 33558 29022
rect 33682 28898 33756 29022
rect 33316 28854 33756 28898
rect 33316 28730 33390 28854
rect 33514 28730 33558 28854
rect 33682 28730 33756 28854
rect 33316 23022 33756 28730
rect 33316 22898 33390 23022
rect 33514 22898 33558 23022
rect 33682 22898 33756 23022
rect 33316 22854 33756 22898
rect 33316 22730 33390 22854
rect 33514 22730 33558 22854
rect 33682 22730 33756 22854
rect 33316 17022 33756 22730
rect 33316 16898 33390 17022
rect 33514 16898 33558 17022
rect 33682 16898 33756 17022
rect 33316 16854 33756 16898
rect 33316 16730 33390 16854
rect 33514 16730 33558 16854
rect 33682 16730 33756 16854
rect 33316 11022 33756 16730
rect 33316 10898 33390 11022
rect 33514 10898 33558 11022
rect 33682 10898 33756 11022
rect 33316 10854 33756 10898
rect 33316 10730 33390 10854
rect 33514 10730 33558 10854
rect 33682 10730 33756 10854
rect 33316 4598 33756 10730
rect 33316 4474 33390 4598
rect 33514 4474 33558 4598
rect 33682 4474 33756 4598
rect 33316 3086 33756 4474
rect 33316 2962 33390 3086
rect 33514 2962 33558 3086
rect 33682 2962 33756 3086
rect 33316 1574 33756 2962
rect 33316 1450 33390 1574
rect 33514 1450 33558 1574
rect 33682 1450 33756 1574
rect 33316 712 33756 1450
rect 34556 38494 34630 38618
rect 34754 38494 34798 38618
rect 34922 38494 34996 38618
rect 49676 38618 50116 38682
rect 34556 37106 34996 38494
rect 34556 36982 34630 37106
rect 34754 36982 34798 37106
rect 34922 36982 34996 37106
rect 34556 35594 34996 36982
rect 34556 35470 34630 35594
rect 34754 35470 34798 35594
rect 34922 35470 34996 35594
rect 34556 34082 34996 35470
rect 34556 33958 34630 34082
rect 34754 33958 34798 34082
rect 34922 33958 34996 34082
rect 34556 24262 34996 33958
rect 34556 24138 34630 24262
rect 34754 24138 34798 24262
rect 34922 24138 34996 24262
rect 34556 24094 34996 24138
rect 34556 23970 34630 24094
rect 34754 23970 34798 24094
rect 34922 23970 34996 24094
rect 34556 18262 34996 23970
rect 34556 18138 34630 18262
rect 34754 18138 34798 18262
rect 34922 18138 34996 18262
rect 34556 18094 34996 18138
rect 34556 17970 34630 18094
rect 34754 17970 34798 18094
rect 34922 17970 34996 18094
rect 34556 12262 34996 17970
rect 34556 12138 34630 12262
rect 34754 12138 34798 12262
rect 34922 12138 34996 12262
rect 34556 12094 34996 12138
rect 34556 11970 34630 12094
rect 34754 11970 34798 12094
rect 34922 11970 34996 12094
rect 34556 5354 34996 11970
rect 34556 5230 34630 5354
rect 34754 5230 34798 5354
rect 34922 5230 34996 5354
rect 34556 3842 34996 5230
rect 34556 3718 34630 3842
rect 34754 3718 34798 3842
rect 34922 3718 34996 3842
rect 34556 2330 34996 3718
rect 34556 2206 34630 2330
rect 34754 2206 34798 2330
rect 34922 2206 34996 2330
rect 34556 818 34996 2206
rect 19436 630 19876 694
rect 34556 694 34630 818
rect 34754 694 34798 818
rect 34922 694 34996 818
rect 48436 37862 48876 38600
rect 48436 37738 48510 37862
rect 48634 37738 48678 37862
rect 48802 37738 48876 37862
rect 48436 36350 48876 37738
rect 48436 36226 48510 36350
rect 48634 36226 48678 36350
rect 48802 36226 48876 36350
rect 48436 34838 48876 36226
rect 48436 34714 48510 34838
rect 48634 34714 48678 34838
rect 48802 34714 48876 34838
rect 48436 29022 48876 34714
rect 48436 28898 48510 29022
rect 48634 28898 48678 29022
rect 48802 28898 48876 29022
rect 48436 28854 48876 28898
rect 48436 28730 48510 28854
rect 48634 28730 48678 28854
rect 48802 28730 48876 28854
rect 48436 23022 48876 28730
rect 48436 22898 48510 23022
rect 48634 22898 48678 23022
rect 48802 22898 48876 23022
rect 48436 22854 48876 22898
rect 48436 22730 48510 22854
rect 48634 22730 48678 22854
rect 48802 22730 48876 22854
rect 48436 17022 48876 22730
rect 48436 16898 48510 17022
rect 48634 16898 48678 17022
rect 48802 16898 48876 17022
rect 48436 16854 48876 16898
rect 48436 16730 48510 16854
rect 48634 16730 48678 16854
rect 48802 16730 48876 16854
rect 48436 11022 48876 16730
rect 48436 10898 48510 11022
rect 48634 10898 48678 11022
rect 48802 10898 48876 11022
rect 48436 10854 48876 10898
rect 48436 10730 48510 10854
rect 48634 10730 48678 10854
rect 48802 10730 48876 10854
rect 48436 4598 48876 10730
rect 48436 4474 48510 4598
rect 48634 4474 48678 4598
rect 48802 4474 48876 4598
rect 48436 3086 48876 4474
rect 48436 2962 48510 3086
rect 48634 2962 48678 3086
rect 48802 2962 48876 3086
rect 48436 1574 48876 2962
rect 48436 1450 48510 1574
rect 48634 1450 48678 1574
rect 48802 1450 48876 1574
rect 48436 712 48876 1450
rect 49676 38494 49750 38618
rect 49874 38494 49918 38618
rect 50042 38494 50116 38618
rect 64796 38618 65236 38682
rect 49676 37106 50116 38494
rect 49676 36982 49750 37106
rect 49874 36982 49918 37106
rect 50042 36982 50116 37106
rect 49676 35594 50116 36982
rect 49676 35470 49750 35594
rect 49874 35470 49918 35594
rect 50042 35470 50116 35594
rect 49676 34082 50116 35470
rect 49676 33958 49750 34082
rect 49874 33958 49918 34082
rect 50042 33958 50116 34082
rect 49676 24262 50116 33958
rect 49676 24138 49750 24262
rect 49874 24138 49918 24262
rect 50042 24138 50116 24262
rect 49676 24094 50116 24138
rect 49676 23970 49750 24094
rect 49874 23970 49918 24094
rect 50042 23970 50116 24094
rect 49676 18262 50116 23970
rect 49676 18138 49750 18262
rect 49874 18138 49918 18262
rect 50042 18138 50116 18262
rect 49676 18094 50116 18138
rect 49676 17970 49750 18094
rect 49874 17970 49918 18094
rect 50042 17970 50116 18094
rect 49676 12262 50116 17970
rect 49676 12138 49750 12262
rect 49874 12138 49918 12262
rect 50042 12138 50116 12262
rect 49676 12094 50116 12138
rect 49676 11970 49750 12094
rect 49874 11970 49918 12094
rect 50042 11970 50116 12094
rect 49676 5354 50116 11970
rect 49676 5230 49750 5354
rect 49874 5230 49918 5354
rect 50042 5230 50116 5354
rect 49676 3842 50116 5230
rect 49676 3718 49750 3842
rect 49874 3718 49918 3842
rect 50042 3718 50116 3842
rect 49676 2330 50116 3718
rect 49676 2206 49750 2330
rect 49874 2206 49918 2330
rect 50042 2206 50116 2330
rect 49676 818 50116 2206
rect 34556 630 34996 694
rect 49676 694 49750 818
rect 49874 694 49918 818
rect 50042 694 50116 818
rect 63556 37862 63996 38600
rect 63556 37738 63630 37862
rect 63754 37738 63798 37862
rect 63922 37738 63996 37862
rect 63556 36350 63996 37738
rect 63556 36226 63630 36350
rect 63754 36226 63798 36350
rect 63922 36226 63996 36350
rect 63556 34838 63996 36226
rect 63556 34714 63630 34838
rect 63754 34714 63798 34838
rect 63922 34714 63996 34838
rect 63556 29022 63996 34714
rect 63556 28898 63630 29022
rect 63754 28898 63798 29022
rect 63922 28898 63996 29022
rect 63556 28854 63996 28898
rect 63556 28730 63630 28854
rect 63754 28730 63798 28854
rect 63922 28730 63996 28854
rect 63556 23022 63996 28730
rect 63556 22898 63630 23022
rect 63754 22898 63798 23022
rect 63922 22898 63996 23022
rect 63556 22854 63996 22898
rect 63556 22730 63630 22854
rect 63754 22730 63798 22854
rect 63922 22730 63996 22854
rect 63556 17022 63996 22730
rect 63556 16898 63630 17022
rect 63754 16898 63798 17022
rect 63922 16898 63996 17022
rect 63556 16854 63996 16898
rect 63556 16730 63630 16854
rect 63754 16730 63798 16854
rect 63922 16730 63996 16854
rect 63556 11022 63996 16730
rect 63556 10898 63630 11022
rect 63754 10898 63798 11022
rect 63922 10898 63996 11022
rect 63556 10854 63996 10898
rect 63556 10730 63630 10854
rect 63754 10730 63798 10854
rect 63922 10730 63996 10854
rect 63556 4598 63996 10730
rect 63556 4474 63630 4598
rect 63754 4474 63798 4598
rect 63922 4474 63996 4598
rect 63556 3086 63996 4474
rect 63556 2962 63630 3086
rect 63754 2962 63798 3086
rect 63922 2962 63996 3086
rect 63556 1574 63996 2962
rect 63556 1450 63630 1574
rect 63754 1450 63798 1574
rect 63922 1450 63996 1574
rect 63556 712 63996 1450
rect 64796 38494 64870 38618
rect 64994 38494 65038 38618
rect 65162 38494 65236 38618
rect 79916 38618 80356 38682
rect 64796 37106 65236 38494
rect 64796 36982 64870 37106
rect 64994 36982 65038 37106
rect 65162 36982 65236 37106
rect 64796 35594 65236 36982
rect 64796 35470 64870 35594
rect 64994 35470 65038 35594
rect 65162 35470 65236 35594
rect 64796 34082 65236 35470
rect 64796 33958 64870 34082
rect 64994 33958 65038 34082
rect 65162 33958 65236 34082
rect 64796 24262 65236 33958
rect 78676 37862 79116 38600
rect 78676 37738 78750 37862
rect 78874 37738 78918 37862
rect 79042 37738 79116 37862
rect 78676 36350 79116 37738
rect 78676 36226 78750 36350
rect 78874 36226 78918 36350
rect 79042 36226 79116 36350
rect 78676 34838 79116 36226
rect 78676 34714 78750 34838
rect 78874 34714 78918 34838
rect 79042 34714 79116 34838
rect 78676 33326 79116 34714
rect 78676 33202 78750 33326
rect 78874 33202 78918 33326
rect 79042 33202 79116 33326
rect 67196 32486 67524 32588
rect 67196 32362 67298 32486
rect 67422 32362 67524 32486
rect 64796 24138 64870 24262
rect 64994 24138 65038 24262
rect 65162 24138 65236 24262
rect 64796 24094 65236 24138
rect 64796 23970 64870 24094
rect 64994 23970 65038 24094
rect 65162 23970 65236 24094
rect 64796 18262 65236 23970
rect 64796 18138 64870 18262
rect 64994 18138 65038 18262
rect 65162 18138 65236 18262
rect 64796 18094 65236 18138
rect 64796 17970 64870 18094
rect 64994 17970 65038 18094
rect 65162 17970 65236 18094
rect 64796 12262 65236 17970
rect 64796 12138 64870 12262
rect 64994 12138 65038 12262
rect 65162 12138 65236 12262
rect 64796 12094 65236 12138
rect 64796 11970 64870 12094
rect 64994 11970 65038 12094
rect 65162 11970 65236 12094
rect 64796 5354 65236 11970
rect 66284 30974 66612 31076
rect 66284 30850 66386 30974
rect 66510 30850 66612 30974
rect 66284 5858 66612 30850
rect 67196 7874 67524 32362
rect 67196 7750 67298 7874
rect 67422 7750 67524 7874
rect 67196 7648 67524 7750
rect 78676 31814 79116 33202
rect 78676 31690 78750 31814
rect 78874 31690 78918 31814
rect 79042 31690 79116 31814
rect 78676 30302 79116 31690
rect 78676 30178 78750 30302
rect 78874 30178 78918 30302
rect 79042 30178 79116 30302
rect 78676 28790 79116 30178
rect 78676 28666 78750 28790
rect 78874 28666 78918 28790
rect 79042 28666 79116 28790
rect 78676 27278 79116 28666
rect 78676 27154 78750 27278
rect 78874 27154 78918 27278
rect 79042 27154 79116 27278
rect 78676 25766 79116 27154
rect 78676 25642 78750 25766
rect 78874 25642 78918 25766
rect 79042 25642 79116 25766
rect 78676 24254 79116 25642
rect 78676 24130 78750 24254
rect 78874 24130 78918 24254
rect 79042 24130 79116 24254
rect 78676 22742 79116 24130
rect 78676 22618 78750 22742
rect 78874 22618 78918 22742
rect 79042 22618 79116 22742
rect 78676 21230 79116 22618
rect 78676 21106 78750 21230
rect 78874 21106 78918 21230
rect 79042 21106 79116 21230
rect 78676 19718 79116 21106
rect 78676 19594 78750 19718
rect 78874 19594 78918 19718
rect 79042 19594 79116 19718
rect 78676 18206 79116 19594
rect 78676 18082 78750 18206
rect 78874 18082 78918 18206
rect 79042 18082 79116 18206
rect 78676 16694 79116 18082
rect 78676 16570 78750 16694
rect 78874 16570 78918 16694
rect 79042 16570 79116 16694
rect 78676 15182 79116 16570
rect 78676 15058 78750 15182
rect 78874 15058 78918 15182
rect 79042 15058 79116 15182
rect 78676 13670 79116 15058
rect 78676 13546 78750 13670
rect 78874 13546 78918 13670
rect 79042 13546 79116 13670
rect 78676 12158 79116 13546
rect 78676 12034 78750 12158
rect 78874 12034 78918 12158
rect 79042 12034 79116 12158
rect 78676 10646 79116 12034
rect 78676 10522 78750 10646
rect 78874 10522 78918 10646
rect 79042 10522 79116 10646
rect 78676 9134 79116 10522
rect 78676 9010 78750 9134
rect 78874 9010 78918 9134
rect 79042 9010 79116 9134
rect 66284 5734 66386 5858
rect 66510 5734 66612 5858
rect 66284 5632 66612 5734
rect 78676 7622 79116 9010
rect 78676 7498 78750 7622
rect 78874 7498 78918 7622
rect 79042 7498 79116 7622
rect 78676 6110 79116 7498
rect 78676 5986 78750 6110
rect 78874 5986 78918 6110
rect 79042 5986 79116 6110
rect 64796 5230 64870 5354
rect 64994 5230 65038 5354
rect 65162 5230 65236 5354
rect 64796 3842 65236 5230
rect 64796 3718 64870 3842
rect 64994 3718 65038 3842
rect 65162 3718 65236 3842
rect 64796 2330 65236 3718
rect 64796 2206 64870 2330
rect 64994 2206 65038 2330
rect 65162 2206 65236 2330
rect 64796 818 65236 2206
rect 49676 630 50116 694
rect 64796 694 64870 818
rect 64994 694 65038 818
rect 65162 694 65236 818
rect 78676 4598 79116 5986
rect 78676 4474 78750 4598
rect 78874 4474 78918 4598
rect 79042 4474 79116 4598
rect 78676 3086 79116 4474
rect 78676 2962 78750 3086
rect 78874 2962 78918 3086
rect 79042 2962 79116 3086
rect 78676 1574 79116 2962
rect 78676 1450 78750 1574
rect 78874 1450 78918 1574
rect 79042 1450 79116 1574
rect 78676 712 79116 1450
rect 79916 38494 79990 38618
rect 80114 38494 80158 38618
rect 80282 38494 80356 38618
rect 79916 37106 80356 38494
rect 79916 36982 79990 37106
rect 80114 36982 80158 37106
rect 80282 36982 80356 37106
rect 79916 35594 80356 36982
rect 79916 35470 79990 35594
rect 80114 35470 80158 35594
rect 80282 35470 80356 35594
rect 79916 34082 80356 35470
rect 79916 33958 79990 34082
rect 80114 33958 80158 34082
rect 80282 33958 80356 34082
rect 79916 32570 80356 33958
rect 79916 32446 79990 32570
rect 80114 32446 80158 32570
rect 80282 32446 80356 32570
rect 79916 31058 80356 32446
rect 79916 30934 79990 31058
rect 80114 30934 80158 31058
rect 80282 30934 80356 31058
rect 79916 29546 80356 30934
rect 79916 29422 79990 29546
rect 80114 29422 80158 29546
rect 80282 29422 80356 29546
rect 79916 28034 80356 29422
rect 79916 27910 79990 28034
rect 80114 27910 80158 28034
rect 80282 27910 80356 28034
rect 79916 26522 80356 27910
rect 79916 26398 79990 26522
rect 80114 26398 80158 26522
rect 80282 26398 80356 26522
rect 79916 25010 80356 26398
rect 79916 24886 79990 25010
rect 80114 24886 80158 25010
rect 80282 24886 80356 25010
rect 79916 23498 80356 24886
rect 79916 23374 79990 23498
rect 80114 23374 80158 23498
rect 80282 23374 80356 23498
rect 79916 21986 80356 23374
rect 79916 21862 79990 21986
rect 80114 21862 80158 21986
rect 80282 21862 80356 21986
rect 79916 20474 80356 21862
rect 79916 20350 79990 20474
rect 80114 20350 80158 20474
rect 80282 20350 80356 20474
rect 79916 18962 80356 20350
rect 79916 18838 79990 18962
rect 80114 18838 80158 18962
rect 80282 18838 80356 18962
rect 79916 17450 80356 18838
rect 79916 17326 79990 17450
rect 80114 17326 80158 17450
rect 80282 17326 80356 17450
rect 79916 15938 80356 17326
rect 79916 15814 79990 15938
rect 80114 15814 80158 15938
rect 80282 15814 80356 15938
rect 79916 14426 80356 15814
rect 79916 14302 79990 14426
rect 80114 14302 80158 14426
rect 80282 14302 80356 14426
rect 79916 12914 80356 14302
rect 79916 12790 79990 12914
rect 80114 12790 80158 12914
rect 80282 12790 80356 12914
rect 79916 11402 80356 12790
rect 79916 11278 79990 11402
rect 80114 11278 80158 11402
rect 80282 11278 80356 11402
rect 79916 9890 80356 11278
rect 79916 9766 79990 9890
rect 80114 9766 80158 9890
rect 80282 9766 80356 9890
rect 79916 8378 80356 9766
rect 79916 8254 79990 8378
rect 80114 8254 80158 8378
rect 80282 8254 80356 8378
rect 79916 6866 80356 8254
rect 79916 6742 79990 6866
rect 80114 6742 80158 6866
rect 80282 6742 80356 6866
rect 79916 5354 80356 6742
rect 79916 5230 79990 5354
rect 80114 5230 80158 5354
rect 80282 5230 80356 5354
rect 79916 3842 80356 5230
rect 79916 3718 79990 3842
rect 80114 3718 80158 3842
rect 80282 3718 80356 3842
rect 79916 2330 80356 3718
rect 79916 2206 79990 2330
rect 80114 2206 80158 2330
rect 80282 2206 80356 2330
rect 79916 818 80356 2206
rect 64796 630 65236 694
rect 79916 694 79990 818
rect 80114 694 80158 818
rect 80282 694 80356 818
rect 93796 34222 94236 38600
rect 93796 34098 93870 34222
rect 93994 34098 94038 34222
rect 94162 34098 94236 34222
rect 93796 34054 94236 34098
rect 93796 33930 93870 34054
rect 93994 33930 94038 34054
rect 94162 33930 94236 34054
rect 93796 28222 94236 33930
rect 93796 28098 93870 28222
rect 93994 28098 94038 28222
rect 94162 28098 94236 28222
rect 93796 28054 94236 28098
rect 93796 27930 93870 28054
rect 93994 27930 94038 28054
rect 94162 27930 94236 28054
rect 93796 21230 94236 27930
rect 93796 21106 93870 21230
rect 93994 21106 94038 21230
rect 94162 21106 94236 21230
rect 93796 19718 94236 21106
rect 93796 19594 93870 19718
rect 93994 19594 94038 19718
rect 94162 19594 94236 19718
rect 93796 11022 94236 19594
rect 93796 10898 93870 11022
rect 93994 10898 94038 11022
rect 94162 10898 94236 11022
rect 93796 10854 94236 10898
rect 93796 10730 93870 10854
rect 93994 10730 94038 10854
rect 94162 10730 94236 10854
rect 93796 5022 94236 10730
rect 93796 4898 93870 5022
rect 93994 4898 94038 5022
rect 94162 4898 94236 5022
rect 93796 4854 94236 4898
rect 93796 4730 93870 4854
rect 93994 4730 94038 4854
rect 94162 4730 94236 4854
rect 93796 712 94236 4730
rect 95036 29462 95476 38600
rect 95036 29338 95110 29462
rect 95234 29338 95278 29462
rect 95402 29338 95476 29462
rect 95036 29294 95476 29338
rect 95036 29170 95110 29294
rect 95234 29170 95278 29294
rect 95402 29170 95476 29294
rect 95036 21986 95476 29170
rect 95036 21862 95110 21986
rect 95234 21862 95278 21986
rect 95402 21862 95476 21986
rect 95036 20474 95476 21862
rect 95036 20350 95110 20474
rect 95234 20350 95278 20474
rect 95402 20350 95476 20474
rect 95036 12262 95476 20350
rect 95036 12138 95110 12262
rect 95234 12138 95278 12262
rect 95402 12138 95476 12262
rect 95036 12094 95476 12138
rect 95036 11970 95110 12094
rect 95234 11970 95278 12094
rect 95402 11970 95476 12094
rect 95036 6262 95476 11970
rect 95036 6138 95110 6262
rect 95234 6138 95278 6262
rect 95402 6138 95476 6262
rect 95036 6094 95476 6138
rect 95036 5970 95110 6094
rect 95234 5970 95278 6094
rect 95402 5970 95476 6094
rect 95036 712 95476 5970
rect 79916 630 80356 694
use sg13g2_inv_1  _128_
timestamp 1676382929
transform 1 0 25920 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_1  _129_
timestamp 1676382929
transform -1 0 35520 0 1 35532
box -48 -56 336 834
use sg13g2_mux2_1  _130_
timestamp 1677247768
transform -1 0 37344 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _131_
timestamp 1677247768
transform 1 0 39744 0 1 35532
box -48 -56 1008 834
use sg13g2_nor2_1  _132_
timestamp 1676627187
transform 1 0 35520 0 1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _133_
timestamp 1683973020
transform 1 0 35904 0 1 3780
box -48 -56 528 834
use sg13g2_nor2b_1  _134_
timestamp 1685181386
transform 1 0 38784 0 1 3780
box -54 -56 528 834
use sg13g2_and2_1  _135_
timestamp 1676901763
transform -1 0 50112 0 -1 5292
box -48 -56 528 834
use sg13g2_and2_1  _136_
timestamp 1676901763
transform -1 0 49920 0 -1 3780
box -48 -56 528 834
use sg13g2_and2_1  _137_
timestamp 1676901763
transform -1 0 49440 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _138_
timestamp 1676627187
transform 1 0 35520 0 1 35532
box -48 -56 432 834
use sg13g2_and2_1  _139_
timestamp 1676901763
transform -1 0 32832 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _140_
timestamp 1685175443
transform -1 0 35040 0 1 3780
box -48 -56 538 834
use sg13g2_nor2_1  _141_
timestamp 1676627187
transform -1 0 37824 0 1 3780
box -48 -56 432 834
use sg13g2_a22oi_1  _142_
timestamp 1685173987
transform 1 0 36672 0 1 3780
box -48 -56 624 834
use sg13g2_o21ai_1  _143_
timestamp 1685175443
transform -1 0 35808 0 -1 5292
box -48 -56 538 834
use sg13g2_nand2_1  _144_
timestamp 1676557249
transform 1 0 38976 0 -1 3780
box -48 -56 432 834
use sg13g2_a22oi_1  _145_
timestamp 1685173987
transform 1 0 31584 0 1 3780
box -48 -56 624 834
use sg13g2_nand2_1  _146_
timestamp 1676557249
transform -1 0 31968 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2_1  _147_
timestamp 1676557249
transform 1 0 49248 0 -1 5292
box -48 -56 432 834
use sg13g2_a22oi_1  _148_
timestamp 1685173987
transform 1 0 33024 0 -1 5292
box -48 -56 624 834
use sg13g2_nand2_1  _149_
timestamp 1676557249
transform -1 0 33024 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2b_1  _150_
timestamp 1676567195
transform -1 0 36288 0 -1 5292
box -48 -56 528 834
use sg13g2_a22oi_1  _151_
timestamp 1685173987
transform 1 0 37536 0 -1 5292
box -48 -56 624 834
use sg13g2_nand2_1  _152_
timestamp 1676557249
transform -1 0 35328 0 -1 5292
box -48 -56 432 834
use sg13g2_mux4_1  _153_
timestamp 1677257233
transform -1 0 41376 0 -1 5292
box -48 -56 2064 834
use sg13g2_nor2b_1  _154_
timestamp 1685181386
transform 1 0 21120 0 1 35532
box -54 -56 528 834
use sg13g2_nand2b_1  _155_
timestamp 1676567195
transform -1 0 20832 0 1 37044
box -48 -56 528 834
use sg13g2_and2_1  _156_
timestamp 1676901763
transform 1 0 24768 0 -1 37044
box -48 -56 528 834
use sg13g2_nor3_1  _157_
timestamp 1676639442
transform 1 0 27456 0 1 35532
box -48 -56 528 834
use sg13g2_nand4_1  _158_
timestamp 1685201930
transform -1 0 27936 0 -1 38556
box -48 -56 624 834
use sg13g2_inv_1  _159_
timestamp 1676382929
transform -1 0 21504 0 -1 37044
box -48 -56 336 834
use sg13g2_nand3_1  _160_
timestamp 1683988354
transform 1 0 21600 0 1 35532
box -48 -56 528 834
use sg13g2_a21o_1  _161_
timestamp 1677175127
transform 1 0 21984 0 -1 37044
box -48 -56 720 834
use sg13g2_and2_1  _162_
timestamp 1676901763
transform -1 0 22176 0 -1 38556
box -48 -56 528 834
use sg13g2_nand3_1  _163_
timestamp 1683988354
transform 1 0 23808 0 -1 37044
box -48 -56 528 834
use sg13g2_xnor2_1  _164_
timestamp 1677516600
transform 1 0 22752 0 -1 37044
box -48 -56 816 834
use sg13g2_and3_1  _165_
timestamp 1676971669
transform -1 0 25920 0 -1 37044
box -48 -56 720 834
use sg13g2_a21oi_1  _166_
timestamp 1683973020
transform -1 0 24768 0 -1 37044
box -48 -56 528 834
use sg13g2_xor2_1  _167_
timestamp 1677577977
transform -1 0 26880 0 -1 37044
box -48 -56 816 834
use sg13g2_and2_1  _168_
timestamp 1676901763
transform -1 0 28224 0 -1 37044
box -48 -56 528 834
use sg13g2_and4_1  _169_
timestamp 1676985977
transform 1 0 26976 0 -1 37044
box -48 -56 816 834
use sg13g2_a21oi_1  _170_
timestamp 1683973020
transform -1 0 26784 0 1 37044
box -48 -56 528 834
use sg13g2_nor2_1  _171_
timestamp 1676627187
transform -1 0 26784 0 -1 38556
box -48 -56 432 834
use sg13g2_nand2_1  _172_
timestamp 1676557249
transform 1 0 29664 0 -1 38556
box -48 -56 432 834
use sg13g2_xor2_1  _173_
timestamp 1677577977
transform 1 0 28896 0 -1 38556
box -48 -56 816 834
use sg13g2_xnor2_1  _174_
timestamp 1677516600
transform 1 0 29376 0 1 37044
box -48 -56 816 834
use sg13g2_mux2_1  _175_
timestamp 1677247768
transform 1 0 22080 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _176_
timestamp 1677247768
transform 1 0 26592 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _177_
timestamp 1677247768
transform -1 0 31104 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _178_
timestamp 1677247768
transform 1 0 31104 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _179_
timestamp 1677247768
transform 1 0 36096 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _180_
timestamp 1677247768
transform 1 0 42912 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _181_
timestamp 1677247768
transform 1 0 48768 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _182_
timestamp 1677247768
transform 1 0 51456 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _183_
timestamp 1677247768
transform 1 0 50496 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _184_
timestamp 1677247768
transform -1 0 47424 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _185_
timestamp 1677247768
transform 1 0 45408 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _186_
timestamp 1677247768
transform 1 0 31392 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _187_
timestamp 1677247768
transform 1 0 33120 0 -1 38556
box -48 -56 1008 834
use sg13g2_mux2_1  _188_
timestamp 1677247768
transform 1 0 33312 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _189_
timestamp 1677247768
transform 1 0 35328 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _190_
timestamp 1677247768
transform -1 0 46944 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _191_
timestamp 1677247768
transform 1 0 47808 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _192_
timestamp 1677247768
transform 1 0 50304 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _193_
timestamp 1677247768
transform 1 0 52032 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _194_
timestamp 1677247768
transform 1 0 47616 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _195_
timestamp 1677247768
transform 1 0 46752 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _196_
timestamp 1677247768
transform 1 0 44352 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _197_
timestamp 1677247768
transform 1 0 43392 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _198_
timestamp 1677247768
transform 1 0 40800 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _199_
timestamp 1677247768
transform 1 0 39648 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _200_
timestamp 1677247768
transform 1 0 38016 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _201_
timestamp 1677247768
transform 1 0 34752 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _202_
timestamp 1677247768
transform -1 0 32928 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _203_
timestamp 1677247768
transform 1 0 27840 0 1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _204_
timestamp 1677247768
transform -1 0 27552 0 1 756
box -48 -56 1008 834
use sg13g2_mux2_1  _205_
timestamp 1677247768
transform -1 0 24864 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _206_
timestamp 1677247768
transform -1 0 21216 0 -1 2268
box -48 -56 1008 834
use sg13g2_mux2_1  _207_
timestamp 1677247768
transform 1 0 21024 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _208_
timestamp 1677247768
transform 1 0 22752 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _209_
timestamp 1677247768
transform -1 0 25248 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _210_
timestamp 1677247768
transform -1 0 27840 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _211_
timestamp 1677247768
transform 1 0 39456 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _212_
timestamp 1677247768
transform 1 0 41760 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _213_
timestamp 1677247768
transform 1 0 43680 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _214_
timestamp 1677247768
transform -1 0 3936 0 -1 21924
box -48 -56 1008 834
use sg13g2_mux2_1  _215_
timestamp 1677247768
transform -1 0 4128 0 -1 23436
box -48 -56 1008 834
use sg13g2_mux2_1  _216_
timestamp 1677247768
transform -1 0 5088 0 -1 23436
box -48 -56 1008 834
use sg13g2_mux2_1  _217_
timestamp 1677247768
transform -1 0 5088 0 -1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  _218_
timestamp 1677247768
transform 1 0 9792 0 1 34020
box -48 -56 1008 834
use sg13g2_mux2_1  _219_
timestamp 1677247768
transform -1 0 13824 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _220_
timestamp 1677247768
transform 1 0 13920 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _221_
timestamp 1677247768
transform 1 0 4320 0 1 27972
box -48 -56 1008 834
use sg13g2_mux2_1  _222_
timestamp 1677247768
transform -1 0 4800 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  _223_
timestamp 1677247768
transform -1 0 3168 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  _224_
timestamp 1677247768
transform -1 0 2304 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _225_
timestamp 1677247768
transform -1 0 2208 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _226_
timestamp 1677247768
transform -1 0 2400 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _227_
timestamp 1677247768
transform 1 0 2112 0 -1 17388
box -48 -56 1008 834
use sg13g2_mux2_1  _228_
timestamp 1677247768
transform 1 0 2400 0 -1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  _229_
timestamp 1677247768
transform -1 0 4512 0 1 18900
box -48 -56 1008 834
use sg13g2_mux2_1  _230_
timestamp 1677247768
transform -1 0 5088 0 1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  _231_
timestamp 1677247768
transform 1 0 16032 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _232_
timestamp 1677247768
transform 1 0 19488 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _233_
timestamp 1677247768
transform 1 0 18336 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _234_
timestamp 1677247768
transform -1 0 18144 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _235_
timestamp 1677247768
transform 1 0 18144 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _236_
timestamp 1677247768
transform -1 0 5184 0 1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _237_
timestamp 1677247768
transform 1 0 2400 0 1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  _238_
timestamp 1677247768
transform -1 0 4416 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _239_
timestamp 1677247768
transform -1 0 4416 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_1  _240_
timestamp 1677247768
transform -1 0 5088 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _241_
timestamp 1677247768
transform -1 0 79008 0 1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _242_
timestamp 1677247768
transform 1 0 80928 0 1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  _243_
timestamp 1677247768
transform 1 0 79776 0 1 27972
box -48 -56 1008 834
use sg13g2_mux2_1  _244_
timestamp 1677247768
transform -1 0 80736 0 1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  _245_
timestamp 1677247768
transform 1 0 79968 0 -1 27972
box -48 -56 1008 834
use sg13g2_mux2_1  _246_
timestamp 1677247768
transform -1 0 80256 0 -1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  _247_
timestamp 1677247768
transform 1 0 79488 0 -1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  _248_
timestamp 1677247768
transform -1 0 81120 0 1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  _249_
timestamp 1677247768
transform -1 0 82080 0 1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  _250_
timestamp 1677247768
transform -1 0 82272 0 1 29484
box -48 -56 1008 834
use sg13g2_mux2_1  _251_
timestamp 1677247768
transform -1 0 81600 0 1 30996
box -48 -56 1008 834
use sg13g2_mux2_1  _252_
timestamp 1677247768
transform -1 0 81408 0 1 32508
box -48 -56 1008 834
use sg13g2_mux2_1  _253_
timestamp 1677247768
transform 1 0 39840 0 -1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _254_
timestamp 1677247768
transform 1 0 40800 0 1 35532
box -48 -56 1008 834
use sg13g2_mux2_1  _255_
timestamp 1677247768
transform 1 0 39456 0 -1 37044
box -48 -56 1008 834
use sg13g2_mux2_1  _256_
timestamp 1677247768
transform -1 0 37152 0 1 37044
box -48 -56 1008 834
use sg13g2_mux2_1  _257_
timestamp 1677247768
transform -1 0 38016 0 -1 38556
box -48 -56 1008 834
use sg13g2_nor2_1  _258_
timestamp 1676627187
transform -1 0 36000 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _259_
timestamp 1683973020
transform 1 0 35904 0 1 35532
box -48 -56 528 834
use sg13g2_nor2_1  _260_
timestamp 1676627187
transform -1 0 35616 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _261_
timestamp 1683973020
transform -1 0 35232 0 1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _262_
timestamp 1677247768
transform -1 0 30912 0 1 2268
box -48 -56 1008 834
use sg13g2_a21o_1  _263_
timestamp 1677175127
transform 1 0 20448 0 1 35532
box -48 -56 720 834
use sg13g2_dfrbpq_1  _264_
timestamp 1746535128
transform 1 0 20928 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _265_
timestamp 1746535128
transform 1 0 23520 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _266_
timestamp 1746535128
transform 1 0 23232 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _267_
timestamp 1746535128
transform 1 0 26016 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _268_
timestamp 1746535128
transform 1 0 26784 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _269_
timestamp 1746535128
transform 1 0 29568 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _270_
timestamp 1746535128
transform 1 0 30144 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _271_
timestamp 1746535128
transform 1 0 23040 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _272_
timestamp 1746535128
transform 1 0 27552 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _273_
timestamp 1746535128
transform 1 0 29952 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _274_
timestamp 1746535128
transform 1 0 32064 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _275_
timestamp 1746535128
transform 1 0 38688 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _276_
timestamp 1746535128
transform 1 0 43872 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _277_
timestamp 1746535128
transform 1 0 49440 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _278_
timestamp 1746535128
transform 1 0 52032 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _279_
timestamp 1746535128
transform 1 0 52704 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _280_
timestamp 1746535128
transform 1 0 46848 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _281_
timestamp 1746535128
transform -1 0 46848 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _282_
timestamp 1746535128
transform 1 0 32640 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _283_
timestamp 1746535128
transform -1 0 35808 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _284_
timestamp 1746535128
transform 1 0 33504 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _285_
timestamp 1746535128
transform 1 0 36576 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _286_
timestamp 1746535128
transform 1 0 45888 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _287_
timestamp 1746535128
transform 1 0 48480 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _288_
timestamp 1746535128
transform 1 0 51072 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _289_
timestamp 1746535128
transform 1 0 52608 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _290_
timestamp 1746535128
transform -1 0 50976 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _291_
timestamp 1746535128
transform -1 0 50304 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _292_
timestamp 1746535128
transform -1 0 47616 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _293_
timestamp 1746535128
transform -1 0 46656 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _294_
timestamp 1746535128
transform 1 0 41760 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _295_
timestamp 1746535128
transform -1 0 42720 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _296_
timestamp 1746535128
transform -1 0 40224 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _297_
timestamp 1746535128
transform -1 0 37440 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _298_
timestamp 1746535128
transform 1 0 32160 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _299_
timestamp 1746535128
transform 1 0 28320 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _300_
timestamp 1746535128
transform 1 0 26784 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _301_
timestamp 1746535128
transform -1 0 26016 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _302_
timestamp 1746535128
transform 1 0 20256 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _303_
timestamp 1746535128
transform 1 0 21216 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _304_
timestamp 1746535128
transform 1 0 23232 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _305_
timestamp 1746535128
transform 1 0 24672 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _306_
timestamp 1746535128
transform 1 0 27264 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _307_
timestamp 1746535128
transform 1 0 40416 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _308_
timestamp 1746535128
transform 1 0 42720 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _309_
timestamp 1746535128
transform -1 0 47232 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _310_
timestamp 1746535128
transform 1 0 2880 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _311_
timestamp 1746535128
transform 1 0 3360 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _312_
timestamp 1746535128
transform 1 0 3360 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _313_
timestamp 1746535128
transform 1 0 3360 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _314_
timestamp 1746535128
transform 1 0 10752 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _315_
timestamp 1746535128
transform 1 0 13344 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _316_
timestamp 1746535128
transform 1 0 14880 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _317_
timestamp 1746535128
transform -1 0 5952 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _318_
timestamp 1746535128
transform 1 0 3360 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _319_
timestamp 1746535128
transform 1 0 2400 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _320_
timestamp 1746535128
transform 1 0 768 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _321_
timestamp 1746535128
transform 1 0 768 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _322_
timestamp 1746535128
transform 1 0 768 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _323_
timestamp 1746535128
transform 1 0 2592 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _324_
timestamp 1746535128
transform 1 0 3360 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _325_
timestamp 1746535128
transform 1 0 3360 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _326_
timestamp 1746535128
transform 1 0 3360 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _327_
timestamp 1746535128
transform 1 0 16800 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _328_
timestamp 1746535128
transform 1 0 20640 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _329_
timestamp 1746535128
transform -1 0 20064 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _330_
timestamp 1746535128
transform 1 0 16800 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _331_
timestamp 1746535128
transform 1 0 19104 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _332_
timestamp 1746535128
transform 1 0 3360 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _333_
timestamp 1746535128
transform 1 0 3360 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _334_
timestamp 1746535128
transform 1 0 3360 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _335_
timestamp 1746535128
transform 1 0 3360 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _336_
timestamp 1746535128
transform 1 0 3360 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _337_
timestamp 1746535128
transform 1 0 78144 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _338_
timestamp 1746535128
transform 1 0 81984 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _339_
timestamp 1746535128
transform 1 0 80736 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _340_
timestamp 1746535128
transform 1 0 80160 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _341_
timestamp 1746535128
transform 1 0 80736 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _342_
timestamp 1746535128
transform 1 0 78720 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _343_
timestamp 1746535128
transform 1 0 80448 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _344_
timestamp 1746535128
transform 1 0 80160 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _345_
timestamp 1746535128
transform 1 0 80736 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _346_
timestamp 1746535128
transform 1 0 80736 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _347_
timestamp 1746535128
transform 1 0 80736 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _348_
timestamp 1746535128
transform 1 0 80736 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _349_
timestamp 1746535128
transform 1 0 40800 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _350_
timestamp 1746535128
transform 1 0 41472 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _351_
timestamp 1746535128
transform -1 0 42432 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _352_
timestamp 1746535128
transform 1 0 36000 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _353_
timestamp 1746535128
transform 1 0 37248 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _354_
timestamp 1746535128
transform 1 0 35904 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _355_
timestamp 1746535128
transform -1 0 35904 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _356_
timestamp 1746535128
transform 1 0 29568 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _357_
timestamp 1746535128
transform 1 0 18624 0 -1 37044
box -48 -56 2640 834
use sg13g2_dlhq_1  _358_
timestamp 1678805552
transform 1 0 29856 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _359_
timestamp 1678805552
transform 1 0 31200 0 -1 3780
box -50 -56 1692 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform -1 0 39360 0 -1 5292
box -48 -56 336 834
use sg13g2_buf_16  clkbuf_0_clk
timestamp 1676553496
transform -1 0 64992 0 1 34020
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_0_clk_regs
timestamp 1676553496
transform 1 0 41472 0 1 34020
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_0__f_clk
timestamp 1676553496
transform 1 0 47424 0 1 34020
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_1__f_clk
timestamp 1676553496
transform -1 0 76416 0 1 27972
box -48 -56 2448 834
use sg13g2_buf_8  clkbuf_4_0_0_clk_regs
timestamp 1676451365
transform -1 0 35904 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_1_0_clk_regs
timestamp 1676451365
transform -1 0 38304 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_2_0_clk_regs
timestamp 1676451365
transform 1 0 24768 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_3_0_clk_regs
timestamp 1676451365
transform -1 0 27264 0 1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_4_0_clk_regs
timestamp 1676451365
transform -1 0 5952 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_5_0_clk_regs
timestamp 1676451365
transform -1 0 8064 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_6_0_clk_regs
timestamp 1676451365
transform 1 0 19392 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_7_0_clk_regs
timestamp 1676451365
transform 1 0 21120 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_8_0_clk_regs
timestamp 1676451365
transform -1 0 51072 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_9_0_clk_regs
timestamp 1676451365
transform -1 0 52704 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_10_0_clk_regs
timestamp 1676451365
transform -1 0 64896 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_11_0_clk_regs
timestamp 1676451365
transform 1 0 61344 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_12_0_clk_regs
timestamp 1676451365
transform -1 0 70464 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_13_0_clk_regs
timestamp 1676451365
transform -1 0 66624 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_14_0_clk_regs
timestamp 1676451365
transform -1 0 69216 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_15_0_clk_regs
timestamp 1676451365
transform 1 0 70464 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_16  clkbuf_regs_0_clk
timestamp 1676553496
transform -1 0 45120 0 -1 5292
box -48 -56 2448 834
use sg13g2_inv_1  clkload0
timestamp 1676382929
transform -1 0 21120 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1676382929
transform 1 0 70080 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_16  delaybuf_0_clk
timestamp 1676553496
transform -1 0 34752 0 1 35532
box -48 -56 2448 834
use sg13g2_buf_1  fanout14
timestamp 1676381911
transform -1 0 2400 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout15
timestamp 1676381911
transform -1 0 3552 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout16
timestamp 1676381911
transform 1 0 20832 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout17
timestamp 1676381911
transform -1 0 10752 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout18
timestamp 1676381911
transform -1 0 20448 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout19
timestamp 1676381911
transform 1 0 22368 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout20
timestamp 1676381911
transform 1 0 32160 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  fanout21
timestamp 1676381911
transform -1 0 32640 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout22
timestamp 1676381911
transform 1 0 26208 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout23
timestamp 1676381911
transform -1 0 19872 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform -1 0 42528 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform -1 0 43776 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform -1 0 80448 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform 1 0 80064 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform 1 0 43872 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform -1 0 22848 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout30
timestamp 1676381911
transform -1 0 2592 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform 1 0 3168 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout32
timestamp 1676381911
transform 1 0 2784 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform 1 0 4320 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform 1 0 13824 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform -1 0 26016 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform -1 0 26400 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform -1 0 24384 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform 1 0 32832 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform -1 0 24768 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform 1 0 23616 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform -1 0 5664 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform 1 0 45120 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout43
timestamp 1676381911
transform 1 0 43872 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform 1 0 79104 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform -1 0 82176 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout46
timestamp 1676381911
transform 1 0 44448 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_266
timestamp 1679577901
transform 1 0 26112 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_270
timestamp 1677579658
transform 1 0 26496 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_281
timestamp 1679581782
transform 1 0 27552 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_288
timestamp 1677579658
transform 1 0 28224 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_316
timestamp 1679581782
transform 1 0 30912 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_323
timestamp 1679577901
transform 1 0 31584 0 1 756
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_337
timestamp 1679581782
transform 1 0 32928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_344
timestamp 1679581782
transform 1 0 33600 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_351
timestamp 1679577901
transform 1 0 34272 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_355
timestamp 1677579658
transform 1 0 34656 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_366
timestamp 1679581782
transform 1 0 35712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_373
timestamp 1679581782
transform 1 0 36384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_380
timestamp 1679581782
transform 1 0 37056 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_387
timestamp 1677580104
transform 1 0 37728 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_389
timestamp 1677579658
transform 1 0 37920 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_400
timestamp 1679581782
transform 1 0 38976 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_407
timestamp 1679577901
transform 1 0 39648 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_411
timestamp 1677579658
transform 1 0 40032 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_439
timestamp 1679581782
transform 1 0 42720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_446
timestamp 1679581782
transform 1 0 43392 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_480
timestamp 1677579658
transform 1 0 46656 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679581782
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679581782
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679581782
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679581782
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679581782
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679581782
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679581782
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679581782
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679581782
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679581782
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679581782
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679581782
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679581782
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679581782
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679581782
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679581782
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679581782
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679581782
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679581782
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679581782
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679581782
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679581782
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679581782
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679581782
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679581782
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679581782
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679581782
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679581782
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679581782
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679581782
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679581782
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679581782
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_833
timestamp 1677580104
transform 1 0 80544 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_203
timestamp 1677580104
transform 1 0 20064 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_215
timestamp 1679581782
transform 1 0 21216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_222
timestamp 1679581782
transform 1 0 21888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_229
timestamp 1679581782
transform 1 0 22560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_236
timestamp 1679581782
transform 1 0 23232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_253
timestamp 1679581782
transform 1 0 24864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_260
timestamp 1679581782
transform 1 0 25536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_267
timestamp 1679577901
transform 1 0 26208 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_271
timestamp 1677580104
transform 1 0 26592 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_300
timestamp 1677580104
transform 1 0 29376 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_356
timestamp 1677579658
transform 1 0 34752 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_384
timestamp 1677580104
transform 1 0 37440 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_413
timestamp 1679577901
transform 1 0 40224 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_417
timestamp 1677580104
transform 1 0 40608 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_456
timestamp 1679581782
transform 1 0 44352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_497
timestamp 1677579658
transform 1 0 48288 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_833
timestamp 1677580104
transform 1 0 80544 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_200
timestamp 1679577901
transform 1 0 19776 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_204
timestamp 1677579658
transform 1 0 20160 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_232
timestamp 1679577901
transform 1 0 22848 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_236
timestamp 1677580104
transform 1 0 23232 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_265
timestamp 1679581782
transform 1 0 26016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_272
timestamp 1679581782
transform 1 0 26688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_279
timestamp 1679577901
transform 1 0 27360 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_283
timestamp 1677579658
transform 1 0 27744 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_294
timestamp 1679581782
transform 1 0 28800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_301
timestamp 1679577901
transform 1 0 29472 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_305
timestamp 1677579658
transform 1 0 29856 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_316
timestamp 1679581782
transform 1 0 30912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_323
timestamp 1679577901
transform 1 0 31584 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_327
timestamp 1677580104
transform 1 0 31968 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_333
timestamp 1679581782
transform 1 0 32544 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_340
timestamp 1677580104
transform 1 0 33216 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_342
timestamp 1677579658
transform 1 0 33408 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_370
timestamp 1679577901
transform 1 0 36096 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_374
timestamp 1677579658
transform 1 0 36480 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_402
timestamp 1679577901
transform 1 0 39168 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_406
timestamp 1677579658
transform 1 0 39552 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_417
timestamp 1679581782
transform 1 0 40608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_424
timestamp 1679581782
transform 1 0 41280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_431
timestamp 1679581782
transform 1 0 41952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_445
timestamp 1677579658
transform 1 0 43296 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_473
timestamp 1679581782
transform 1 0 45984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_487
timestamp 1677580104
transform 1 0 47328 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_489
timestamp 1677579658
transform 1 0 47520 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_500
timestamp 1679581782
transform 1 0 48576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_507
timestamp 1679581782
transform 1 0 49248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_514
timestamp 1679581782
transform 1 0 49920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_521
timestamp 1679581782
transform 1 0 50592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_528
timestamp 1679581782
transform 1 0 51264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_535
timestamp 1679581782
transform 1 0 51936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_542
timestamp 1679581782
transform 1 0 52608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_549
timestamp 1679581782
transform 1 0 53280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_556
timestamp 1679581782
transform 1 0 53952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_563
timestamp 1679581782
transform 1 0 54624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_570
timestamp 1679581782
transform 1 0 55296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_577
timestamp 1679581782
transform 1 0 55968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_584
timestamp 1679581782
transform 1 0 56640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_591
timestamp 1679581782
transform 1 0 57312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_598
timestamp 1679581782
transform 1 0 57984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_605
timestamp 1679581782
transform 1 0 58656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_612
timestamp 1679581782
transform 1 0 59328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_619
timestamp 1679581782
transform 1 0 60000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_626
timestamp 1679581782
transform 1 0 60672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_633
timestamp 1679581782
transform 1 0 61344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_640
timestamp 1679581782
transform 1 0 62016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_647
timestamp 1679581782
transform 1 0 62688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_654
timestamp 1679581782
transform 1 0 63360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_661
timestamp 1679581782
transform 1 0 64032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_668
timestamp 1679581782
transform 1 0 64704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_675
timestamp 1679581782
transform 1 0 65376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_682
timestamp 1679581782
transform 1 0 66048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_689
timestamp 1679581782
transform 1 0 66720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_696
timestamp 1679581782
transform 1 0 67392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_703
timestamp 1679581782
transform 1 0 68064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_710
timestamp 1679581782
transform 1 0 68736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_717
timestamp 1679581782
transform 1 0 69408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_724
timestamp 1679581782
transform 1 0 70080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_731
timestamp 1679581782
transform 1 0 70752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_738
timestamp 1679581782
transform 1 0 71424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_745
timestamp 1679581782
transform 1 0 72096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_752
timestamp 1679581782
transform 1 0 72768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_759
timestamp 1679581782
transform 1 0 73440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_766
timestamp 1679581782
transform 1 0 74112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_773
timestamp 1679581782
transform 1 0 74784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_780
timestamp 1679581782
transform 1 0 75456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_787
timestamp 1679581782
transform 1 0 76128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_794
timestamp 1679581782
transform 1 0 76800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_801
timestamp 1679581782
transform 1 0 77472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_808
timestamp 1679581782
transform 1 0 78144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_815
timestamp 1679581782
transform 1 0 78816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_822
timestamp 1679581782
transform 1 0 79488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_829
timestamp 1679577901
transform 1 0 80160 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_833
timestamp 1677580104
transform 1 0 80544 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 13728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 15744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679581782
transform 1 0 16416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679581782
transform 1 0 17088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 17760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679581782
transform 1 0 18432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679581782
transform 1 0 19104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_200
timestamp 1679581782
transform 1 0 19776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_207
timestamp 1679577901
transform 1 0 20448 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_211
timestamp 1677580104
transform 1 0 20832 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_223
timestamp 1679581782
transform 1 0 21984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_230
timestamp 1679577901
transform 1 0 22656 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_234
timestamp 1677580104
transform 1 0 23040 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_263
timestamp 1679581782
transform 1 0 25824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_270
timestamp 1679577901
transform 1 0 26496 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_284
timestamp 1679581782
transform 1 0 27840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_291
timestamp 1679581782
transform 1 0 28512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679581782
transform 1 0 29184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679581782
transform 1 0 29856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_312
timestamp 1679581782
transform 1 0 30528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_336
timestamp 1679577901
transform 1 0 32832 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_340
timestamp 1677579658
transform 1 0 33216 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_351
timestamp 1679581782
transform 1 0 34272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_358
timestamp 1679577901
transform 1 0 34944 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_372
timestamp 1679581782
transform 1 0 36288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_379
timestamp 1679581782
transform 1 0 36960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_386
timestamp 1679581782
transform 1 0 37632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_393
timestamp 1679581782
transform 1 0 38304 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_404
timestamp 1677579658
transform 1 0 39360 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_442
timestamp 1679581782
transform 1 0 43008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_486
timestamp 1679577901
transform 1 0 47232 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_490
timestamp 1677580104
transform 1 0 47616 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_502
timestamp 1677580104
transform 1 0 48768 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_514
timestamp 1679577901
transform 1 0 49920 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_528
timestamp 1679581782
transform 1 0 51264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_535
timestamp 1679581782
transform 1 0 51936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_569
timestamp 1679581782
transform 1 0 55200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_576
timestamp 1679581782
transform 1 0 55872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_583
timestamp 1679581782
transform 1 0 56544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_590
timestamp 1679581782
transform 1 0 57216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_597
timestamp 1679581782
transform 1 0 57888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_604
timestamp 1679581782
transform 1 0 58560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_611
timestamp 1679581782
transform 1 0 59232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_618
timestamp 1679581782
transform 1 0 59904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_625
timestamp 1679581782
transform 1 0 60576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_632
timestamp 1679581782
transform 1 0 61248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_639
timestamp 1679581782
transform 1 0 61920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_646
timestamp 1679581782
transform 1 0 62592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_653
timestamp 1679581782
transform 1 0 63264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_660
timestamp 1679581782
transform 1 0 63936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_667
timestamp 1679581782
transform 1 0 64608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_674
timestamp 1679581782
transform 1 0 65280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_681
timestamp 1679581782
transform 1 0 65952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_688
timestamp 1679581782
transform 1 0 66624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_695
timestamp 1679581782
transform 1 0 67296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_702
timestamp 1679581782
transform 1 0 67968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_709
timestamp 1679581782
transform 1 0 68640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_716
timestamp 1679581782
transform 1 0 69312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_723
timestamp 1679581782
transform 1 0 69984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_730
timestamp 1679581782
transform 1 0 70656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_737
timestamp 1679581782
transform 1 0 71328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_744
timestamp 1679581782
transform 1 0 72000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_751
timestamp 1679581782
transform 1 0 72672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_758
timestamp 1679581782
transform 1 0 73344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_765
timestamp 1679581782
transform 1 0 74016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_772
timestamp 1679581782
transform 1 0 74688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_779
timestamp 1679581782
transform 1 0 75360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_786
timestamp 1679581782
transform 1 0 76032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_793
timestamp 1679581782
transform 1 0 76704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_800
timestamp 1679581782
transform 1 0 77376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_807
timestamp 1679581782
transform 1 0 78048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_814
timestamp 1679581782
transform 1 0 78720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_821
timestamp 1679581782
transform 1 0 79392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_828
timestamp 1679581782
transform 1 0 80064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_109
timestamp 1679581782
transform 1 0 11040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_116
timestamp 1679581782
transform 1 0 11712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_123
timestamp 1679581782
transform 1 0 12384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679581782
transform 1 0 13056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 15744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_165
timestamp 1679577901
transform 1 0 16416 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_196
timestamp 1679581782
transform 1 0 19392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_203
timestamp 1679581782
transform 1 0 20064 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_210
timestamp 1677579658
transform 1 0 20736 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_242
timestamp 1679581782
transform 1 0 23808 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_249
timestamp 1677580104
transform 1 0 24480 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_322
timestamp 1677579658
transform 1 0 31488 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_329
timestamp 1677580104
transform 1 0 32160 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_336
timestamp 1679581782
transform 1 0 32832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_343
timestamp 1679581782
transform 1 0 33504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_350
timestamp 1679577901
transform 1 0 34176 0 1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_4_359
timestamp 1679577901
transform 1 0 35040 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_363
timestamp 1677579658
transform 1 0 35424 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_373
timestamp 1677580104
transform 1 0 36384 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_375
timestamp 1677579658
transform 1 0 36576 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_382
timestamp 1677580104
transform 1 0 37248 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_388
timestamp 1679581782
transform 1 0 37824 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_395
timestamp 1677580104
transform 1 0 38496 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_397
timestamp 1677579658
transform 1 0 38688 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_403
timestamp 1679581782
transform 1 0 39264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_410
timestamp 1679581782
transform 1 0 39936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_417
timestamp 1679581782
transform 1 0 40608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_424
timestamp 1679577901
transform 1 0 41280 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_428
timestamp 1677579658
transform 1 0 41664 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_466
timestamp 1679577901
transform 1 0 45312 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_470
timestamp 1677580104
transform 1 0 45696 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_553
timestamp 1679581782
transform 1 0 53664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_560
timestamp 1679581782
transform 1 0 54336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_567
timestamp 1679581782
transform 1 0 55008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_574
timestamp 1679581782
transform 1 0 55680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_581
timestamp 1679581782
transform 1 0 56352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_588
timestamp 1679581782
transform 1 0 57024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_595
timestamp 1679581782
transform 1 0 57696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_602
timestamp 1679581782
transform 1 0 58368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_609
timestamp 1679581782
transform 1 0 59040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_616
timestamp 1679581782
transform 1 0 59712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_623
timestamp 1679581782
transform 1 0 60384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_630
timestamp 1679581782
transform 1 0 61056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_637
timestamp 1679581782
transform 1 0 61728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_644
timestamp 1679581782
transform 1 0 62400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_651
timestamp 1679581782
transform 1 0 63072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_658
timestamp 1679581782
transform 1 0 63744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_665
timestamp 1679581782
transform 1 0 64416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_672
timestamp 1679581782
transform 1 0 65088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_679
timestamp 1679581782
transform 1 0 65760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_686
timestamp 1679581782
transform 1 0 66432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_693
timestamp 1679581782
transform 1 0 67104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_700
timestamp 1679581782
transform 1 0 67776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_707
timestamp 1679581782
transform 1 0 68448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_714
timestamp 1679581782
transform 1 0 69120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_721
timestamp 1679581782
transform 1 0 69792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_728
timestamp 1679581782
transform 1 0 70464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_735
timestamp 1679581782
transform 1 0 71136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_742
timestamp 1679581782
transform 1 0 71808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_749
timestamp 1679581782
transform 1 0 72480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_756
timestamp 1679581782
transform 1 0 73152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_763
timestamp 1679581782
transform 1 0 73824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_770
timestamp 1679581782
transform 1 0 74496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_777
timestamp 1679581782
transform 1 0 75168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_784
timestamp 1679581782
transform 1 0 75840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_791
timestamp 1679581782
transform 1 0 76512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_798
timestamp 1679581782
transform 1 0 77184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_805
timestamp 1679581782
transform 1 0 77856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_812
timestamp 1679581782
transform 1 0 78528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_819
timestamp 1679581782
transform 1 0 79200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_826
timestamp 1679581782
transform 1 0 79872 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_833
timestamp 1677580104
transform 1 0 80544 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_158
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_165
timestamp 1679581782
transform 1 0 16416 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_172
timestamp 1677579658
transform 1 0 17088 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_220
timestamp 1679581782
transform 1 0 21696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_241
timestamp 1679577901
transform 1 0 23712 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_245
timestamp 1677580104
transform 1 0 24096 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_257
timestamp 1679577901
transform 1 0 25248 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_269
timestamp 1679581782
transform 1 0 26400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_276
timestamp 1679581782
transform 1 0 27072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_283
timestamp 1679581782
transform 1 0 27744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_290
timestamp 1679581782
transform 1 0 28416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_297
timestamp 1679581782
transform 1 0 29088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_304
timestamp 1679581782
transform 1 0 29760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_311
timestamp 1679581782
transform 1 0 30432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_318
timestamp 1679577901
transform 1 0 31104 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_322
timestamp 1677579658
transform 1 0 31488 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_327
timestamp 1679581782
transform 1 0 31968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_344
timestamp 1679581782
transform 1 0 33600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_351
timestamp 1679581782
transform 1 0 34272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_372
timestamp 1679581782
transform 1 0 36288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_379
timestamp 1679577901
transform 1 0 36960 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_383
timestamp 1677580104
transform 1 0 37344 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_391
timestamp 1679581782
transform 1 0 38112 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_398
timestamp 1677580104
transform 1 0 38784 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_400
timestamp 1677579658
transform 1 0 38976 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_425
timestamp 1679581782
transform 1 0 41376 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_432
timestamp 1677579658
transform 1 0 42048 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_437
timestamp 1677580104
transform 1 0 42528 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_468
timestamp 1679577901
transform 1 0 45504 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_472
timestamp 1677579658
transform 1 0 45888 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_483
timestamp 1679581782
transform 1 0 46944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_490
timestamp 1679581782
transform 1 0 47616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_497
timestamp 1679581782
transform 1 0 48288 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_504
timestamp 1677580104
transform 1 0 48960 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_506
timestamp 1677579658
transform 1 0 49152 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_516
timestamp 1679581782
transform 1 0 50112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_523
timestamp 1679581782
transform 1 0 50784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_530
timestamp 1679577901
transform 1 0 51456 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_534
timestamp 1677580104
transform 1 0 51840 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_546
timestamp 1679581782
transform 1 0 52992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_553
timestamp 1679581782
transform 1 0 53664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_560
timestamp 1679581782
transform 1 0 54336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_567
timestamp 1679581782
transform 1 0 55008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_574
timestamp 1679581782
transform 1 0 55680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_581
timestamp 1679581782
transform 1 0 56352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_588
timestamp 1679581782
transform 1 0 57024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_595
timestamp 1679581782
transform 1 0 57696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_602
timestamp 1679581782
transform 1 0 58368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_609
timestamp 1679581782
transform 1 0 59040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_616
timestamp 1679581782
transform 1 0 59712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_623
timestamp 1679581782
transform 1 0 60384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_630
timestamp 1679581782
transform 1 0 61056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_637
timestamp 1679581782
transform 1 0 61728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_644
timestamp 1679581782
transform 1 0 62400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_651
timestamp 1679581782
transform 1 0 63072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_658
timestamp 1679581782
transform 1 0 63744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_665
timestamp 1679581782
transform 1 0 64416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_672
timestamp 1679581782
transform 1 0 65088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_679
timestamp 1679581782
transform 1 0 65760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_686
timestamp 1679581782
transform 1 0 66432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_693
timestamp 1679581782
transform 1 0 67104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_700
timestamp 1679581782
transform 1 0 67776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_707
timestamp 1679581782
transform 1 0 68448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_714
timestamp 1679581782
transform 1 0 69120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_721
timestamp 1679581782
transform 1 0 69792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_728
timestamp 1679581782
transform 1 0 70464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_735
timestamp 1679581782
transform 1 0 71136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_742
timestamp 1679581782
transform 1 0 71808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_749
timestamp 1679581782
transform 1 0 72480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_756
timestamp 1679581782
transform 1 0 73152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_763
timestamp 1679581782
transform 1 0 73824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_770
timestamp 1679581782
transform 1 0 74496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_777
timestamp 1679581782
transform 1 0 75168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_784
timestamp 1679581782
transform 1 0 75840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_791
timestamp 1679581782
transform 1 0 76512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_798
timestamp 1679581782
transform 1 0 77184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_805
timestamp 1679581782
transform 1 0 77856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_812
timestamp 1679581782
transform 1 0 78528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_819
timestamp 1679581782
transform 1 0 79200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_826
timestamp 1679581782
transform 1 0 79872 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_833
timestamp 1677580104
transform 1 0 80544 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679581782
transform 1 0 3648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679581782
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679581782
transform 1 0 4992 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_53
timestamp 1677580104
transform 1 0 5664 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_55
timestamp 1677579658
transform 1 0 5856 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_765
timestamp 1679581782
transform 1 0 74016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_772
timestamp 1679581782
transform 1 0 74688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_779
timestamp 1679581782
transform 1 0 75360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_786
timestamp 1679581782
transform 1 0 76032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_793
timestamp 1679581782
transform 1 0 76704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_800
timestamp 1679581782
transform 1 0 77376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_807
timestamp 1679581782
transform 1 0 78048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_814
timestamp 1679581782
transform 1 0 78720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_821
timestamp 1679581782
transform 1 0 79392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_828
timestamp 1679581782
transform 1 0 80064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_765
timestamp 1679581782
transform 1 0 74016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_772
timestamp 1679581782
transform 1 0 74688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_779
timestamp 1679581782
transform 1 0 75360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_786
timestamp 1679581782
transform 1 0 76032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_793
timestamp 1679581782
transform 1 0 76704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_800
timestamp 1679581782
transform 1 0 77376 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_807
timestamp 1677580104
transform 1 0 78048 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_809
timestamp 1677579658
transform 1 0 78240 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_32
timestamp 1679577901
transform 1 0 3648 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_36
timestamp 1677580104
transform 1 0 4032 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_48
timestamp 1679581782
transform 1 0 5184 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_55
timestamp 1677579658
transform 1 0 5856 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_765
timestamp 1679581782
transform 1 0 74016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_772
timestamp 1679581782
transform 1 0 74688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_779
timestamp 1679581782
transform 1 0 75360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_786
timestamp 1679581782
transform 1 0 76032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_793
timestamp 1679581782
transform 1 0 76704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_800
timestamp 1679581782
transform 1 0 77376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_807
timestamp 1679581782
transform 1 0 78048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_814
timestamp 1679581782
transform 1 0 78720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_821
timestamp 1679581782
transform 1 0 79392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_828
timestamp 1679581782
transform 1 0 80064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_25
timestamp 1679577901
transform 1 0 2976 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_765
timestamp 1679581782
transform 1 0 74016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_772
timestamp 1679581782
transform 1 0 74688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_779
timestamp 1679581782
transform 1 0 75360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_786
timestamp 1679581782
transform 1 0 76032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_793
timestamp 1679581782
transform 1 0 76704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_800
timestamp 1679581782
transform 1 0 77376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_807
timestamp 1679581782
transform 1 0 78048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_814
timestamp 1679581782
transform 1 0 78720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_821
timestamp 1679581782
transform 1 0 79392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_828
timestamp 1679581782
transform 1 0 80064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679581782
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679581782
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679581782
transform 1 0 2976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679581782
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679581782
transform 1 0 4320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_46
timestamp 1679581782
transform 1 0 4992 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_53
timestamp 1677580104
transform 1 0 5664 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_55
timestamp 1677579658
transform 1 0 5856 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_765
timestamp 1679581782
transform 1 0 74016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_772
timestamp 1679581782
transform 1 0 74688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_779
timestamp 1679581782
transform 1 0 75360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_786
timestamp 1679581782
transform 1 0 76032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_793
timestamp 1679581782
transform 1 0 76704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_800
timestamp 1679581782
transform 1 0 77376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_807
timestamp 1679581782
transform 1 0 78048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_814
timestamp 1679581782
transform 1 0 78720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_821
timestamp 1679581782
transform 1 0 79392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_828
timestamp 1679581782
transform 1 0 80064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_25
timestamp 1679577901
transform 1 0 2976 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_765
timestamp 1679581782
transform 1 0 74016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_772
timestamp 1679581782
transform 1 0 74688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_779
timestamp 1679581782
transform 1 0 75360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_786
timestamp 1679581782
transform 1 0 76032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_793
timestamp 1679581782
transform 1 0 76704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_800
timestamp 1679581782
transform 1 0 77376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_807
timestamp 1679581782
transform 1 0 78048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_814
timestamp 1679581782
transform 1 0 78720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_821
timestamp 1679581782
transform 1 0 79392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_828
timestamp 1679581782
transform 1 0 80064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679581782
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_11
timestamp 1679577901
transform 1 0 1632 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_15
timestamp 1677580104
transform 1 0 2016 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_27
timestamp 1679581782
transform 1 0 3168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_44
timestamp 1679581782
transform 1 0 4800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_51
timestamp 1679577901
transform 1 0 5472 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_55
timestamp 1677579658
transform 1 0 5856 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_765
timestamp 1679581782
transform 1 0 74016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_772
timestamp 1679581782
transform 1 0 74688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_779
timestamp 1679581782
transform 1 0 75360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_786
timestamp 1679581782
transform 1 0 76032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_793
timestamp 1679581782
transform 1 0 76704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_800
timestamp 1679581782
transform 1 0 77376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_807
timestamp 1679581782
transform 1 0 78048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_814
timestamp 1679581782
transform 1 0 78720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_821
timestamp 1679581782
transform 1 0 79392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_828
timestamp 1679581782
transform 1 0 80064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679581782
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_18
timestamp 1677579658
transform 1 0 2304 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679581782
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_53
timestamp 1677580104
transform 1 0 5664 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_55
timestamp 1677579658
transform 1 0 5856 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_765
timestamp 1679581782
transform 1 0 74016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_772
timestamp 1679581782
transform 1 0 74688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_779
timestamp 1679581782
transform 1 0 75360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_786
timestamp 1679581782
transform 1 0 76032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_793
timestamp 1679581782
transform 1 0 76704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_800
timestamp 1679581782
transform 1 0 77376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_807
timestamp 1679581782
transform 1 0 78048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_814
timestamp 1679581782
transform 1 0 78720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_821
timestamp 1679581782
transform 1 0 79392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_828
timestamp 1679581782
transform 1 0 80064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679581782
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_18
timestamp 1677579658
transform 1 0 2304 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_765
timestamp 1679581782
transform 1 0 74016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_772
timestamp 1679581782
transform 1 0 74688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_779
timestamp 1679581782
transform 1 0 75360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_786
timestamp 1679581782
transform 1 0 76032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_793
timestamp 1679581782
transform 1 0 76704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_800
timestamp 1679581782
transform 1 0 77376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_807
timestamp 1679581782
transform 1 0 78048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_814
timestamp 1679581782
transform 1 0 78720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_821
timestamp 1679581782
transform 1 0 79392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_828
timestamp 1679581782
transform 1 0 80064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679581782
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_25
timestamp 1679577901
transform 1 0 2976 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_29
timestamp 1677579658
transform 1 0 3360 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_40
timestamp 1679581782
transform 1 0 4416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_47
timestamp 1679581782
transform 1 0 5088 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_54
timestamp 1677580104
transform 1 0 5760 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_765
timestamp 1679581782
transform 1 0 74016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_772
timestamp 1679581782
transform 1 0 74688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_779
timestamp 1679581782
transform 1 0 75360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_786
timestamp 1679581782
transform 1 0 76032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_793
timestamp 1679581782
transform 1 0 76704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_800
timestamp 1679581782
transform 1 0 77376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_807
timestamp 1679581782
transform 1 0 78048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_814
timestamp 1679581782
transform 1 0 78720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_821
timestamp 1679581782
transform 1 0 79392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_828
timestamp 1679581782
transform 1 0 80064 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_0
timestamp 1677580104
transform 1 0 576 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_765
timestamp 1679581782
transform 1 0 74016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_772
timestamp 1679581782
transform 1 0 74688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_779
timestamp 1679581782
transform 1 0 75360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_786
timestamp 1679581782
transform 1 0 76032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_793
timestamp 1679581782
transform 1 0 76704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_800
timestamp 1679581782
transform 1 0 77376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_807
timestamp 1679581782
transform 1 0 78048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_814
timestamp 1679581782
transform 1 0 78720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_821
timestamp 1679581782
transform 1 0 79392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_828
timestamp 1679581782
transform 1 0 80064 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_4
timestamp 1677580104
transform 1 0 960 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_6
timestamp 1677579658
transform 1 0 1152 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_17
timestamp 1679581782
transform 1 0 2208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_24
timestamp 1679577901
transform 1 0 2880 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_28
timestamp 1677580104
transform 1 0 3264 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_40
timestamp 1679581782
transform 1 0 4416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_47
timestamp 1679581782
transform 1 0 5088 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_54
timestamp 1677580104
transform 1 0 5760 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_765
timestamp 1679581782
transform 1 0 74016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_772
timestamp 1679581782
transform 1 0 74688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_779
timestamp 1679581782
transform 1 0 75360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_786
timestamp 1679581782
transform 1 0 76032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_793
timestamp 1679581782
transform 1 0 76704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_800
timestamp 1679581782
transform 1 0 77376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_807
timestamp 1679581782
transform 1 0 78048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_814
timestamp 1679581782
transform 1 0 78720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_821
timestamp 1679581782
transform 1 0 79392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_828
timestamp 1679581782
transform 1 0 80064 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_0
timestamp 1677580104
transform 1 0 576 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_765
timestamp 1679581782
transform 1 0 74016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_772
timestamp 1679581782
transform 1 0 74688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_779
timestamp 1679581782
transform 1 0 75360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_786
timestamp 1679581782
transform 1 0 76032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_793
timestamp 1679581782
transform 1 0 76704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_800
timestamp 1679581782
transform 1 0 77376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_807
timestamp 1679581782
transform 1 0 78048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_814
timestamp 1679581782
transform 1 0 78720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_821
timestamp 1679581782
transform 1 0 79392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_828
timestamp 1679581782
transform 1 0 80064 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_8
timestamp 1677579658
transform 1 0 1344 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_19
timestamp 1679581782
transform 1 0 2400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_26
timestamp 1679581782
transform 1 0 3072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_33
timestamp 1679577901
transform 1 0 3744 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_47
timestamp 1679581782
transform 1 0 5088 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_54
timestamp 1677580104
transform 1 0 5760 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_765
timestamp 1679581782
transform 1 0 74016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_772
timestamp 1679581782
transform 1 0 74688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_779
timestamp 1679581782
transform 1 0 75360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_786
timestamp 1679581782
transform 1 0 76032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_793
timestamp 1679581782
transform 1 0 76704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_800
timestamp 1679581782
transform 1 0 77376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_807
timestamp 1679581782
transform 1 0 78048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_814
timestamp 1679581782
transform 1 0 78720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_821
timestamp 1679581782
transform 1 0 79392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_828
timestamp 1679581782
transform 1 0 80064 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_0
timestamp 1677580104
transform 1 0 576 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_765
timestamp 1679581782
transform 1 0 74016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_772
timestamp 1679581782
transform 1 0 74688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_779
timestamp 1679581782
transform 1 0 75360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_786
timestamp 1679581782
transform 1 0 76032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_793
timestamp 1679581782
transform 1 0 76704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_800
timestamp 1679581782
transform 1 0 77376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_817
timestamp 1679581782
transform 1 0 79008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_824
timestamp 1679581782
transform 1 0 79680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_831
timestamp 1679577901
transform 1 0 80352 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_11
timestamp 1679577901
transform 1 0 1632 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_15
timestamp 1677579658
transform 1 0 2016 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_26
timestamp 1677579658
transform 1 0 3072 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_31
timestamp 1679581782
transform 1 0 3552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_38
timestamp 1679581782
transform 1 0 4224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_45
timestamp 1679581782
transform 1 0 4896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_52
timestamp 1679577901
transform 1 0 5568 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_765
timestamp 1679581782
transform 1 0 74016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_772
timestamp 1679581782
transform 1 0 74688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_779
timestamp 1679581782
transform 1 0 75360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_786
timestamp 1679581782
transform 1 0 76032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_793
timestamp 1679581782
transform 1 0 76704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_800
timestamp 1679581782
transform 1 0 77376 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_807
timestamp 1677579658
transform 1 0 78048 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679581782
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_11
timestamp 1679577901
transform 1 0 1632 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_15
timestamp 1677580104
transform 1 0 2016 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_48
timestamp 1679581782
transform 1 0 5184 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_55
timestamp 1677579658
transform 1 0 5856 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_765
timestamp 1679581782
transform 1 0 74016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_772
timestamp 1679581782
transform 1 0 74688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_779
timestamp 1679581782
transform 1 0 75360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_786
timestamp 1679581782
transform 1 0 76032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_793
timestamp 1679581782
transform 1 0 76704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_800
timestamp 1679581782
transform 1 0 77376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_807
timestamp 1679581782
transform 1 0 78048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_814
timestamp 1679581782
transform 1 0 78720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_821
timestamp 1679581782
transform 1 0 79392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_828
timestamp 1679581782
transform 1 0 80064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_11
timestamp 1679577901
transform 1 0 1632 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_765
timestamp 1679581782
transform 1 0 74016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_772
timestamp 1679581782
transform 1 0 74688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_779
timestamp 1679581782
transform 1 0 75360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_786
timestamp 1679581782
transform 1 0 76032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_793
timestamp 1679581782
transform 1 0 76704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_800
timestamp 1679581782
transform 1 0 77376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_807
timestamp 1679581782
transform 1 0 78048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_814
timestamp 1679581782
transform 1 0 78720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_821
timestamp 1679581782
transform 1 0 79392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_828
timestamp 1679581782
transform 1 0 80064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_18
timestamp 1679577901
transform 1 0 2304 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_22
timestamp 1677579658
transform 1 0 2688 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_41
timestamp 1679581782
transform 1 0 4512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_48
timestamp 1679581782
transform 1 0 5184 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_55
timestamp 1677579658
transform 1 0 5856 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_765
timestamp 1679581782
transform 1 0 74016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_772
timestamp 1679581782
transform 1 0 74688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_779
timestamp 1679581782
transform 1 0 75360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_786
timestamp 1679581782
transform 1 0 76032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_793
timestamp 1679581782
transform 1 0 76704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_800
timestamp 1679581782
transform 1 0 77376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_807
timestamp 1679581782
transform 1 0 78048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_814
timestamp 1679581782
transform 1 0 78720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_821
timestamp 1679581782
transform 1 0 79392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_828
timestamp 1679581782
transform 1 0 80064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_25
timestamp 1679577901
transform 1 0 2976 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_765
timestamp 1679581782
transform 1 0 74016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_772
timestamp 1679581782
transform 1 0 74688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_779
timestamp 1679581782
transform 1 0 75360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_786
timestamp 1679581782
transform 1 0 76032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_793
timestamp 1679581782
transform 1 0 76704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_800
timestamp 1679581782
transform 1 0 77376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_807
timestamp 1679581782
transform 1 0 78048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_814
timestamp 1679581782
transform 1 0 78720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_821
timestamp 1679581782
transform 1 0 79392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_828
timestamp 1679581782
transform 1 0 80064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_835
timestamp 1679581782
transform 1 0 80736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_842
timestamp 1679581782
transform 1 0 81408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_849
timestamp 1679581782
transform 1 0 82080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_856
timestamp 1679581782
transform 1 0 82752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_863
timestamp 1679581782
transform 1 0 83424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_870
timestamp 1679581782
transform 1 0 84096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_877
timestamp 1679581782
transform 1 0 84768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_884
timestamp 1679581782
transform 1 0 85440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_891
timestamp 1679581782
transform 1 0 86112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_898
timestamp 1679581782
transform 1 0 86784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_905
timestamp 1679581782
transform 1 0 87456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_912
timestamp 1679581782
transform 1 0 88128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_919
timestamp 1679581782
transform 1 0 88800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_926
timestamp 1679581782
transform 1 0 89472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_933
timestamp 1679581782
transform 1 0 90144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_940
timestamp 1679581782
transform 1 0 90816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_947
timestamp 1679581782
transform 1 0 91488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_954
timestamp 1679581782
transform 1 0 92160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_961
timestamp 1679581782
transform 1 0 92832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_968
timestamp 1679581782
transform 1 0 93504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_975
timestamp 1679581782
transform 1 0 94176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_982
timestamp 1679581782
transform 1 0 94848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_989
timestamp 1679581782
transform 1 0 95520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_996
timestamp 1679577901
transform 1 0 96192 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_1025
timestamp 1679577901
transform 1 0 98976 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_18
timestamp 1679577901
transform 1 0 2304 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_22
timestamp 1677580104
transform 1 0 2688 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_51
timestamp 1679577901
transform 1 0 5472 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_55
timestamp 1677579658
transform 1 0 5856 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_765
timestamp 1679581782
transform 1 0 74016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_772
timestamp 1679581782
transform 1 0 74688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_779
timestamp 1679581782
transform 1 0 75360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_786
timestamp 1679581782
transform 1 0 76032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_793
timestamp 1679581782
transform 1 0 76704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_800
timestamp 1679581782
transform 1 0 77376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_807
timestamp 1679581782
transform 1 0 78048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_814
timestamp 1679581782
transform 1 0 78720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_821
timestamp 1679581782
transform 1 0 79392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_828
timestamp 1679581782
transform 1 0 80064 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_835
timestamp 1677580104
transform 1 0 80736 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_847
timestamp 1677579658
transform 1 0 81888 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_875
timestamp 1679581782
transform 1 0 84576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_882
timestamp 1679581782
transform 1 0 85248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_889
timestamp 1679581782
transform 1 0 85920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_896
timestamp 1679581782
transform 1 0 86592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_903
timestamp 1679581782
transform 1 0 87264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_910
timestamp 1679581782
transform 1 0 87936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_917
timestamp 1679581782
transform 1 0 88608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_924
timestamp 1679581782
transform 1 0 89280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_931
timestamp 1679581782
transform 1 0 89952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_938
timestamp 1679581782
transform 1 0 90624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_945
timestamp 1679581782
transform 1 0 91296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_952
timestamp 1679581782
transform 1 0 91968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_959
timestamp 1679581782
transform 1 0 92640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_966
timestamp 1679581782
transform 1 0 93312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_973
timestamp 1679581782
transform 1 0 93984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_980
timestamp 1679581782
transform 1 0 94656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_987
timestamp 1679581782
transform 1 0 95328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_994
timestamp 1679581782
transform 1 0 96000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1001
timestamp 1679581782
transform 1 0 96672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1008
timestamp 1679581782
transform 1 0 97344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1015
timestamp 1679581782
transform 1 0 98016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1022
timestamp 1679581782
transform 1 0 98688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_21
timestamp 1679577901
transform 1 0 2592 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679581782
transform 1 0 3936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_42
timestamp 1679581782
transform 1 0 4608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_49
timestamp 1679581782
transform 1 0 5280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_765
timestamp 1679581782
transform 1 0 74016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_772
timestamp 1679581782
transform 1 0 74688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_779
timestamp 1679581782
transform 1 0 75360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_786
timestamp 1679581782
transform 1 0 76032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_793
timestamp 1679581782
transform 1 0 76704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_800
timestamp 1679581782
transform 1 0 77376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_807
timestamp 1679581782
transform 1 0 78048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_814
timestamp 1679581782
transform 1 0 78720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_821
timestamp 1679581782
transform 1 0 79392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_828
timestamp 1679581782
transform 1 0 80064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_835
timestamp 1679581782
transform 1 0 80736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_842
timestamp 1679581782
transform 1 0 81408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_849
timestamp 1679581782
transform 1 0 82080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_856
timestamp 1679581782
transform 1 0 82752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_863
timestamp 1679581782
transform 1 0 83424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_870
timestamp 1679581782
transform 1 0 84096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_877
timestamp 1679581782
transform 1 0 84768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_884
timestamp 1679581782
transform 1 0 85440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_891
timestamp 1679581782
transform 1 0 86112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_898
timestamp 1679581782
transform 1 0 86784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_905
timestamp 1679581782
transform 1 0 87456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_912
timestamp 1679581782
transform 1 0 88128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_919
timestamp 1679581782
transform 1 0 88800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_926
timestamp 1679581782
transform 1 0 89472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_933
timestamp 1679581782
transform 1 0 90144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_940
timestamp 1679581782
transform 1 0 90816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_947
timestamp 1679581782
transform 1 0 91488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_954
timestamp 1679581782
transform 1 0 92160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_961
timestamp 1679581782
transform 1 0 92832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_968
timestamp 1679581782
transform 1 0 93504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_975
timestamp 1679581782
transform 1 0 94176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_982
timestamp 1679581782
transform 1 0 94848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_989
timestamp 1679581782
transform 1 0 95520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_996
timestamp 1679581782
transform 1 0 96192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1003
timestamp 1679581782
transform 1 0 96864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1010
timestamp 1679581782
transform 1 0 97536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1017
timestamp 1679581782
transform 1 0 98208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_1024
timestamp 1679577901
transform 1 0 98880 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_1028
timestamp 1677579658
transform 1 0 99264 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_25
timestamp 1679577901
transform 1 0 2976 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_765
timestamp 1679581782
transform 1 0 74016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_772
timestamp 1679581782
transform 1 0 74688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_779
timestamp 1679581782
transform 1 0 75360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_786
timestamp 1679581782
transform 1 0 76032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_793
timestamp 1679581782
transform 1 0 76704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_800
timestamp 1679581782
transform 1 0 77376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_807
timestamp 1679581782
transform 1 0 78048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_814
timestamp 1679581782
transform 1 0 78720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_821
timestamp 1679581782
transform 1 0 79392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_828
timestamp 1679581782
transform 1 0 80064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_835
timestamp 1679581782
transform 1 0 80736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_842
timestamp 1679581782
transform 1 0 81408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_849
timestamp 1679581782
transform 1 0 82080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_856
timestamp 1679577901
transform 1 0 82752 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_860
timestamp 1677580104
transform 1 0 83136 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_4
timestamp 1679581782
transform 1 0 960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_11
timestamp 1679581782
transform 1 0 1632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_18
timestamp 1679581782
transform 1 0 2304 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_25
timestamp 1677580104
transform 1 0 2976 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_47
timestamp 1679581782
transform 1 0 5088 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_54
timestamp 1677580104
transform 1 0 5760 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_765
timestamp 1679581782
transform 1 0 74016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_772
timestamp 1679581782
transform 1 0 74688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_779
timestamp 1679581782
transform 1 0 75360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_786
timestamp 1679581782
transform 1 0 76032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_793
timestamp 1679581782
transform 1 0 76704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_800
timestamp 1679581782
transform 1 0 77376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_807
timestamp 1679581782
transform 1 0 78048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_814
timestamp 1679581782
transform 1 0 78720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_821
timestamp 1679581782
transform 1 0 79392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_828
timestamp 1679581782
transform 1 0 80064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_835
timestamp 1679581782
transform 1 0 80736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_842
timestamp 1679581782
transform 1 0 81408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_849
timestamp 1679581782
transform 1 0 82080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_856
timestamp 1679577901
transform 1 0 82752 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_860
timestamp 1677580104
transform 1 0 83136 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_4
timestamp 1679581782
transform 1 0 960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_11
timestamp 1679581782
transform 1 0 1632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_18
timestamp 1679581782
transform 1 0 2304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_25
timestamp 1679577901
transform 1 0 2976 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_765
timestamp 1679581782
transform 1 0 74016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_772
timestamp 1679581782
transform 1 0 74688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_779
timestamp 1679581782
transform 1 0 75360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_786
timestamp 1679581782
transform 1 0 76032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_793
timestamp 1679581782
transform 1 0 76704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_800
timestamp 1679581782
transform 1 0 77376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_807
timestamp 1679581782
transform 1 0 78048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_814
timestamp 1679581782
transform 1 0 78720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_821
timestamp 1679581782
transform 1 0 79392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_828
timestamp 1679581782
transform 1 0 80064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_4
timestamp 1679581782
transform 1 0 960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_11
timestamp 1679581782
transform 1 0 1632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_18
timestamp 1679581782
transform 1 0 2304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_25
timestamp 1679581782
transform 1 0 2976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_32
timestamp 1679581782
transform 1 0 3648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_39
timestamp 1679581782
transform 1 0 4320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_46
timestamp 1679581782
transform 1 0 4992 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_53
timestamp 1677580104
transform 1 0 5664 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_55
timestamp 1677579658
transform 1 0 5856 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_765
timestamp 1679581782
transform 1 0 74016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_772
timestamp 1679581782
transform 1 0 74688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_779
timestamp 1679581782
transform 1 0 75360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_786
timestamp 1679581782
transform 1 0 76032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_793
timestamp 1679581782
transform 1 0 76704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_800
timestamp 1679581782
transform 1 0 77376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_807
timestamp 1679581782
transform 1 0 78048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_814
timestamp 1679581782
transform 1 0 78720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_821
timestamp 1679581782
transform 1 0 79392 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_828
timestamp 1677579658
transform 1 0 80064 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_856
timestamp 1679577901
transform 1 0 82752 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_860
timestamp 1677580104
transform 1 0 83136 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_11
timestamp 1679581782
transform 1 0 1632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_18
timestamp 1679581782
transform 1 0 2304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_25
timestamp 1679581782
transform 1 0 2976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_32
timestamp 1679577901
transform 1 0 3648 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_36
timestamp 1677579658
transform 1 0 4032 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_47
timestamp 1679581782
transform 1 0 5088 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_54
timestamp 1677580104
transform 1 0 5760 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_765
timestamp 1679581782
transform 1 0 74016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_772
timestamp 1679581782
transform 1 0 74688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_779
timestamp 1679581782
transform 1 0 75360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_786
timestamp 1679581782
transform 1 0 76032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_793
timestamp 1679581782
transform 1 0 76704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_800
timestamp 1679581782
transform 1 0 77376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_807
timestamp 1679581782
transform 1 0 78048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_814
timestamp 1679581782
transform 1 0 78720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_821
timestamp 1679581782
transform 1 0 79392 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_828
timestamp 1677579658
transform 1 0 80064 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_849
timestamp 1679581782
transform 1 0 82080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_856
timestamp 1679577901
transform 1 0 82752 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_860
timestamp 1677580104
transform 1 0 83136 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679581782
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679581782
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679581782
transform 1 0 1920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679581782
transform 1 0 2592 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_28
timestamp 1677579658
transform 1 0 3264 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_765
timestamp 1679581782
transform 1 0 74016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_772
timestamp 1679581782
transform 1 0 74688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_779
timestamp 1679581782
transform 1 0 75360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_786
timestamp 1679581782
transform 1 0 76032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_793
timestamp 1679581782
transform 1 0 76704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_800
timestamp 1679581782
transform 1 0 77376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_807
timestamp 1679581782
transform 1 0 78048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_814
timestamp 1679581782
transform 1 0 78720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_821
timestamp 1679581782
transform 1 0 79392 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_828
timestamp 1677579658
transform 1 0 80064 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_856
timestamp 1679577901
transform 1 0 82752 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_860
timestamp 1677580104
transform 1 0 83136 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679581782
transform 1 0 3936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679581782
transform 1 0 4608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_765
timestamp 1679581782
transform 1 0 74016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_772
timestamp 1679581782
transform 1 0 74688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_779
timestamp 1679581782
transform 1 0 75360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_786
timestamp 1679581782
transform 1 0 76032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_793
timestamp 1679581782
transform 1 0 76704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_800
timestamp 1679581782
transform 1 0 77376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_807
timestamp 1679581782
transform 1 0 78048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_814
timestamp 1679581782
transform 1 0 78720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_821
timestamp 1679577901
transform 1 0 79392 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679581782
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_765
timestamp 1679581782
transform 1 0 74016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_772
timestamp 1679581782
transform 1 0 74688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_779
timestamp 1679581782
transform 1 0 75360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_786
timestamp 1679581782
transform 1 0 76032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_793
timestamp 1679581782
transform 1 0 76704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_800
timestamp 1679581782
transform 1 0 77376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_807
timestamp 1679581782
transform 1 0 78048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_814
timestamp 1679581782
transform 1 0 78720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_821
timestamp 1679577901
transform 1 0 79392 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_825
timestamp 1677580104
transform 1 0 79776 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_837
timestamp 1679581782
transform 1 0 80928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_844
timestamp 1679581782
transform 1 0 81600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_851
timestamp 1679581782
transform 1 0 82272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_858
timestamp 1679577901
transform 1 0 82944 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_35
timestamp 1679577901
transform 1 0 3936 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_790
timestamp 1679581782
transform 1 0 76416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_797
timestamp 1679581782
transform 1 0 77088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_804
timestamp 1679581782
transform 1 0 77760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_811
timestamp 1679581782
transform 1 0 78432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_818
timestamp 1679581782
transform 1 0 79104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_28
timestamp 1677579658
transform 1 0 3264 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_765
timestamp 1679581782
transform 1 0 74016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_772
timestamp 1679581782
transform 1 0 74688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_779
timestamp 1679581782
transform 1 0 75360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_786
timestamp 1679581782
transform 1 0 76032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_793
timestamp 1679581782
transform 1 0 76704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_800
timestamp 1679581782
transform 1 0 77376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_807
timestamp 1679581782
transform 1 0 78048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_814
timestamp 1679577901
transform 1 0 78720 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_818
timestamp 1677580104
transform 1 0 79104 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_830
timestamp 1679577901
transform 1 0 80256 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_834
timestamp 1677579658
transform 1 0 80640 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_765
timestamp 1679581782
transform 1 0 74016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_772
timestamp 1679581782
transform 1 0 74688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_779
timestamp 1679581782
transform 1 0 75360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_786
timestamp 1679581782
transform 1 0 76032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_793
timestamp 1679581782
transform 1 0 76704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_800
timestamp 1679581782
transform 1 0 77376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_807
timestamp 1679581782
transform 1 0 78048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_851
timestamp 1679581782
transform 1 0 82272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_858
timestamp 1679577901
transform 1 0 82944 0 1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_35
timestamp 1677580104
transform 1 0 3936 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_47
timestamp 1679581782
transform 1 0 5088 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_54
timestamp 1677580104
transform 1 0 5760 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_765
timestamp 1679581782
transform 1 0 74016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_772
timestamp 1679581782
transform 1 0 74688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_779
timestamp 1679581782
transform 1 0 75360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_786
timestamp 1679581782
transform 1 0 76032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_793
timestamp 1679581782
transform 1 0 76704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_800
timestamp 1679581782
transform 1 0 77376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_807
timestamp 1679581782
transform 1 0 78048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_814
timestamp 1679577901
transform 1 0 78720 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_859
timestamp 1677580104
transform 1 0 83040 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_861
timestamp 1677579658
transform 1 0 83232 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_28
timestamp 1677579658
transform 1 0 3264 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_765
timestamp 1679581782
transform 1 0 74016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_772
timestamp 1679581782
transform 1 0 74688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_779
timestamp 1679581782
transform 1 0 75360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_786
timestamp 1679581782
transform 1 0 76032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_793
timestamp 1679581782
transform 1 0 76704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_800
timestamp 1679581782
transform 1 0 77376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_807
timestamp 1679581782
transform 1 0 78048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_814
timestamp 1679581782
transform 1 0 78720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_821
timestamp 1679581782
transform 1 0 79392 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_832
timestamp 1677580104
transform 1 0 80448 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_844
timestamp 1679581782
transform 1 0 81600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_851
timestamp 1679581782
transform 1 0 82272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_858
timestamp 1679577901
transform 1 0 82944 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_35
timestamp 1679577901
transform 1 0 3936 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_765
timestamp 1679581782
transform 1 0 74016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_772
timestamp 1679581782
transform 1 0 74688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_779
timestamp 1679581782
transform 1 0 75360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_786
timestamp 1679581782
transform 1 0 76032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_793
timestamp 1679581782
transform 1 0 76704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_800
timestamp 1679581782
transform 1 0 77376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_807
timestamp 1679581782
transform 1 0 78048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_814
timestamp 1679581782
transform 1 0 78720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_821
timestamp 1679581782
transform 1 0 79392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_828
timestamp 1679581782
transform 1 0 80064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_53
timestamp 1677580104
transform 1 0 5664 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_55
timestamp 1677579658
transform 1 0 5856 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_765
timestamp 1679581782
transform 1 0 74016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_772
timestamp 1679581782
transform 1 0 74688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_779
timestamp 1679581782
transform 1 0 75360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_786
timestamp 1679581782
transform 1 0 76032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_793
timestamp 1679581782
transform 1 0 76704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_800
timestamp 1679581782
transform 1 0 77376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_807
timestamp 1679581782
transform 1 0 78048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_814
timestamp 1679581782
transform 1 0 78720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_821
timestamp 1679581782
transform 1 0 79392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_842
timestamp 1679577901
transform 1 0 81408 0 1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_42_850
timestamp 1679581782
transform 1 0 82176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_857
timestamp 1679577901
transform 1 0 82848 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_861
timestamp 1677579658
transform 1 0 83232 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_765
timestamp 1679581782
transform 1 0 74016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_772
timestamp 1679581782
transform 1 0 74688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_779
timestamp 1679581782
transform 1 0 75360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_786
timestamp 1679581782
transform 1 0 76032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_793
timestamp 1679581782
transform 1 0 76704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_800
timestamp 1679581782
transform 1 0 77376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_807
timestamp 1679581782
transform 1 0 78048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_814
timestamp 1679581782
transform 1 0 78720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_821
timestamp 1679581782
transform 1 0 79392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_828
timestamp 1679581782
transform 1 0 80064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_63
timestamp 1677580104
transform 1 0 6624 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_78
timestamp 1679581782
transform 1 0 8064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_85
timestamp 1679581782
transform 1 0 8736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_92
timestamp 1679577901
transform 1 0 9408 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_160
timestamp 1679581782
transform 1 0 15936 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_167
timestamp 1677580104
transform 1 0 16608 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_209
timestamp 1677580104
transform 1 0 20640 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_227
timestamp 1679581782
transform 1 0 22368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_261
timestamp 1679577901
transform 1 0 25632 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_265
timestamp 1677580104
transform 1 0 26016 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_368
timestamp 1677580104
transform 1 0 35904 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_393
timestamp 1679577901
transform 1 0 38304 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_424
timestamp 1677580104
transform 1 0 41280 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_526
timestamp 1679577901
transform 1 0 51072 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_570
timestamp 1679581782
transform 1 0 55296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_577
timestamp 1679581782
transform 1 0 55968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_584
timestamp 1679581782
transform 1 0 56640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_591
timestamp 1679581782
transform 1 0 57312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_598
timestamp 1679581782
transform 1 0 57984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_605
timestamp 1679581782
transform 1 0 58656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_612
timestamp 1679581782
transform 1 0 59328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_619
timestamp 1679581782
transform 1 0 60000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_626
timestamp 1679581782
transform 1 0 60672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_671
timestamp 1679577901
transform 1 0 64992 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_688
timestamp 1679581782
transform 1 0 66624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_695
timestamp 1679581782
transform 1 0 67296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_741
timestamp 1679581782
transform 1 0 71712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_748
timestamp 1679581782
transform 1 0 72384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_755
timestamp 1679581782
transform 1 0 73056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_762
timestamp 1679581782
transform 1 0 73728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_769
timestamp 1679581782
transform 1 0 74400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_776
timestamp 1679581782
transform 1 0 75072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_783
timestamp 1679581782
transform 1 0 75744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_790
timestamp 1679581782
transform 1 0 76416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_797
timestamp 1679581782
transform 1 0 77088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_804
timestamp 1679581782
transform 1 0 77760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_811
timestamp 1679581782
transform 1 0 78432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_818
timestamp 1679581782
transform 1 0 79104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_825
timestamp 1679581782
transform 1 0 79776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_832
timestamp 1679581782
transform 1 0 80448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_839
timestamp 1679581782
transform 1 0 81120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_846
timestamp 1679581782
transform 1 0 81792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_853
timestamp 1679581782
transform 1 0 82464 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_860
timestamp 1677580104
transform 1 0 83136 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_98
timestamp 1679577901
transform 1 0 9984 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_106
timestamp 1679581782
transform 1 0 10752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_113
timestamp 1679581782
transform 1 0 11424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_120
timestamp 1679581782
transform 1 0 12096 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_127
timestamp 1677579658
transform 1 0 12768 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_138
timestamp 1677579658
transform 1 0 13824 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_207
timestamp 1677580104
transform 1 0 20448 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_236
timestamp 1679581782
transform 1 0 23232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_243
timestamp 1679581782
transform 1 0 23904 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_250
timestamp 1677580104
transform 1 0 24576 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_292
timestamp 1679581782
transform 1 0 28608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_299
timestamp 1679581782
transform 1 0 29280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_333
timestamp 1679581782
transform 1 0 32544 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_340
timestamp 1677579658
transform 1 0 33216 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_395
timestamp 1679581782
transform 1 0 38496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_402
timestamp 1679581782
transform 1 0 39168 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_450
timestamp 1677579658
transform 1 0 43776 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_563
timestamp 1679581782
transform 1 0 54624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_570
timestamp 1679581782
transform 1 0 55296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_577
timestamp 1679581782
transform 1 0 55968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_584
timestamp 1679581782
transform 1 0 56640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_591
timestamp 1679581782
transform 1 0 57312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_598
timestamp 1679581782
transform 1 0 57984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_605
timestamp 1679581782
transform 1 0 58656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_612
timestamp 1679581782
transform 1 0 59328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_619
timestamp 1679581782
transform 1 0 60000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_626
timestamp 1679581782
transform 1 0 60672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_633
timestamp 1679581782
transform 1 0 61344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_640
timestamp 1679581782
transform 1 0 62016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_647
timestamp 1679581782
transform 1 0 62688 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_654
timestamp 1677580104
transform 1 0 63360 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_656
timestamp 1677579658
transform 1 0 63552 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_670
timestamp 1679581782
transform 1 0 64896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_677
timestamp 1679581782
transform 1 0 65568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_684
timestamp 1679581782
transform 1 0 66240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_691
timestamp 1679581782
transform 1 0 66912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_698
timestamp 1679581782
transform 1 0 67584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_705
timestamp 1679581782
transform 1 0 68256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_712
timestamp 1679581782
transform 1 0 68928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_719
timestamp 1679577901
transform 1 0 69600 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_723
timestamp 1677579658
transform 1 0 69984 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_727
timestamp 1679581782
transform 1 0 70368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_734
timestamp 1679581782
transform 1 0 71040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_741
timestamp 1679581782
transform 1 0 71712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_748
timestamp 1679581782
transform 1 0 72384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_755
timestamp 1679581782
transform 1 0 73056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_762
timestamp 1679581782
transform 1 0 73728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_769
timestamp 1679581782
transform 1 0 74400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_776
timestamp 1679581782
transform 1 0 75072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_783
timestamp 1679581782
transform 1 0 75744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_790
timestamp 1679581782
transform 1 0 76416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_797
timestamp 1679581782
transform 1 0 77088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_804
timestamp 1679581782
transform 1 0 77760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_811
timestamp 1679581782
transform 1 0 78432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_818
timestamp 1679581782
transform 1 0 79104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_825
timestamp 1679581782
transform 1 0 79776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_832
timestamp 1679581782
transform 1 0 80448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_839
timestamp 1679581782
transform 1 0 81120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_846
timestamp 1679581782
transform 1 0 81792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_853
timestamp 1679581782
transform 1 0 82464 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_860
timestamp 1677580104
transform 1 0 83136 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_133
timestamp 1679577901
transform 1 0 13344 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_137
timestamp 1677579658
transform 1 0 13728 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_142
timestamp 1679581782
transform 1 0 14208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_149
timestamp 1679581782
transform 1 0 14880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_156
timestamp 1679577901
transform 1 0 15552 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_160
timestamp 1677579658
transform 1 0 15936 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_171
timestamp 1679581782
transform 1 0 16992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_178
timestamp 1679581782
transform 1 0 17664 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_195
timestamp 1677580104
transform 1 0 19296 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_234
timestamp 1677580104
transform 1 0 23040 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_263
timestamp 1677580104
transform 1 0 25824 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_278
timestamp 1677580104
transform 1 0 27264 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_285
timestamp 1679581782
transform 1 0 27936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_292
timestamp 1679581782
transform 1 0 28608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_299
timestamp 1679581782
transform 1 0 29280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_306
timestamp 1679581782
transform 1 0 29952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_313
timestamp 1679581782
transform 1 0 30624 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_320
timestamp 1677579658
transform 1 0 31296 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_383
timestamp 1679581782
transform 1 0 37344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_390
timestamp 1679581782
transform 1 0 38016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_397
timestamp 1679581782
transform 1 0 38688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_404
timestamp 1679577901
transform 1 0 39360 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_418
timestamp 1677579658
transform 1 0 40704 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_429
timestamp 1679581782
transform 1 0 41760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_436
timestamp 1679577901
transform 1 0 42432 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_440
timestamp 1677579658
transform 1 0 42816 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_455
timestamp 1677580104
transform 1 0 44256 0 1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_46_461
timestamp 1679577901
transform 1 0 44832 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_465
timestamp 1677580104
transform 1 0 45216 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_477
timestamp 1679581782
transform 1 0 46368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_484
timestamp 1679581782
transform 1 0 47040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_491
timestamp 1679581782
transform 1 0 47712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_498
timestamp 1679577901
transform 1 0 48384 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_512
timestamp 1679581782
transform 1 0 49728 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_519
timestamp 1677579658
transform 1 0 50400 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_540
timestamp 1679581782
transform 1 0 52416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_547
timestamp 1679581782
transform 1 0 53088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_554
timestamp 1679581782
transform 1 0 53760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_561
timestamp 1679581782
transform 1 0 54432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_568
timestamp 1679581782
transform 1 0 55104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_575
timestamp 1679581782
transform 1 0 55776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_582
timestamp 1679581782
transform 1 0 56448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_589
timestamp 1679581782
transform 1 0 57120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_596
timestamp 1679581782
transform 1 0 57792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_603
timestamp 1679581782
transform 1 0 58464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_610
timestamp 1679581782
transform 1 0 59136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_617
timestamp 1679581782
transform 1 0 59808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_624
timestamp 1679581782
transform 1 0 60480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_631
timestamp 1679581782
transform 1 0 61152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_638
timestamp 1679581782
transform 1 0 61824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_645
timestamp 1679581782
transform 1 0 62496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_652
timestamp 1679581782
transform 1 0 63168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_659
timestamp 1679581782
transform 1 0 63840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_666
timestamp 1679581782
transform 1 0 64512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_673
timestamp 1679581782
transform 1 0 65184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_680
timestamp 1679581782
transform 1 0 65856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_687
timestamp 1679581782
transform 1 0 66528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_694
timestamp 1679581782
transform 1 0 67200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_701
timestamp 1679581782
transform 1 0 67872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_708
timestamp 1679581782
transform 1 0 68544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_715
timestamp 1679581782
transform 1 0 69216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_722
timestamp 1679581782
transform 1 0 69888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_729
timestamp 1679581782
transform 1 0 70560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_736
timestamp 1679581782
transform 1 0 71232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_743
timestamp 1679581782
transform 1 0 71904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_750
timestamp 1679581782
transform 1 0 72576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_757
timestamp 1679581782
transform 1 0 73248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_764
timestamp 1679581782
transform 1 0 73920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_771
timestamp 1679581782
transform 1 0 74592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_778
timestamp 1679581782
transform 1 0 75264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_785
timestamp 1679581782
transform 1 0 75936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_792
timestamp 1679581782
transform 1 0 76608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_799
timestamp 1679581782
transform 1 0 77280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_806
timestamp 1679581782
transform 1 0 77952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_813
timestamp 1679581782
transform 1 0 78624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_820
timestamp 1679581782
transform 1 0 79296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_827
timestamp 1679581782
transform 1 0 79968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_834
timestamp 1679581782
transform 1 0 80640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_841
timestamp 1679581782
transform 1 0 81312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_848
timestamp 1679581782
transform 1 0 81984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_855
timestamp 1679581782
transform 1 0 82656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_182
timestamp 1679577901
transform 1 0 18048 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_186
timestamp 1677580104
transform 1 0 18432 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_4  FILLER_47_218
timestamp 1679577901
transform 1 0 21504 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_222
timestamp 1677579658
transform 1 0 21888 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_230
timestamp 1677579658
transform 1 0 22656 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_239
timestamp 1677580104
transform 1 0 23520 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_241
timestamp 1677579658
transform 1 0 23712 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_264
timestamp 1677580104
transform 1 0 25920 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_274
timestamp 1677579658
transform 1 0 26880 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_288
timestamp 1679581782
transform 1 0 28224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_295
timestamp 1679581782
transform 1 0 28896 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_329
timestamp 1677579658
transform 1 0 32160 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_396
timestamp 1679581782
transform 1 0 38592 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_403
timestamp 1677580104
transform 1 0 39264 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_415
timestamp 1679581782
transform 1 0 40416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_422
timestamp 1679577901
transform 1 0 41088 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_47_453
timestamp 1679581782
transform 1 0 44064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_460
timestamp 1679581782
transform 1 0 44736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_467
timestamp 1679581782
transform 1 0 45408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_474
timestamp 1679581782
transform 1 0 46080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_481
timestamp 1679581782
transform 1 0 46752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_488
timestamp 1679581782
transform 1 0 47424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_495
timestamp 1679581782
transform 1 0 48096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_502
timestamp 1679581782
transform 1 0 48768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_509
timestamp 1679581782
transform 1 0 49440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_516
timestamp 1679581782
transform 1 0 50112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_523
timestamp 1679581782
transform 1 0 50784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_530
timestamp 1679581782
transform 1 0 51456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_537
timestamp 1679581782
transform 1 0 52128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_544
timestamp 1679581782
transform 1 0 52800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_551
timestamp 1679581782
transform 1 0 53472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_558
timestamp 1679581782
transform 1 0 54144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_565
timestamp 1679581782
transform 1 0 54816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_572
timestamp 1679581782
transform 1 0 55488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_579
timestamp 1679581782
transform 1 0 56160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_586
timestamp 1679581782
transform 1 0 56832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_593
timestamp 1679581782
transform 1 0 57504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_600
timestamp 1679581782
transform 1 0 58176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_607
timestamp 1679581782
transform 1 0 58848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_614
timestamp 1679581782
transform 1 0 59520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_621
timestamp 1679581782
transform 1 0 60192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_628
timestamp 1679581782
transform 1 0 60864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_635
timestamp 1679581782
transform 1 0 61536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_642
timestamp 1679581782
transform 1 0 62208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_649
timestamp 1679581782
transform 1 0 62880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_656
timestamp 1679581782
transform 1 0 63552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_663
timestamp 1679581782
transform 1 0 64224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_670
timestamp 1679581782
transform 1 0 64896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_677
timestamp 1679581782
transform 1 0 65568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_684
timestamp 1679581782
transform 1 0 66240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_691
timestamp 1679581782
transform 1 0 66912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_698
timestamp 1679581782
transform 1 0 67584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_705
timestamp 1679581782
transform 1 0 68256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_712
timestamp 1679581782
transform 1 0 68928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_719
timestamp 1679581782
transform 1 0 69600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_726
timestamp 1679581782
transform 1 0 70272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_733
timestamp 1679581782
transform 1 0 70944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_740
timestamp 1679581782
transform 1 0 71616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_747
timestamp 1679581782
transform 1 0 72288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_754
timestamp 1679581782
transform 1 0 72960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_761
timestamp 1679581782
transform 1 0 73632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_768
timestamp 1679581782
transform 1 0 74304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_775
timestamp 1679581782
transform 1 0 74976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_782
timestamp 1679581782
transform 1 0 75648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_789
timestamp 1679581782
transform 1 0 76320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_796
timestamp 1679581782
transform 1 0 76992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_803
timestamp 1679581782
transform 1 0 77664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_810
timestamp 1679581782
transform 1 0 78336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_817
timestamp 1679581782
transform 1 0 79008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_824
timestamp 1679581782
transform 1 0 79680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_831
timestamp 1679581782
transform 1 0 80352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_838
timestamp 1679581782
transform 1 0 81024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_845
timestamp 1679581782
transform 1 0 81696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_852
timestamp 1679581782
transform 1 0 82368 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_859
timestamp 1677580104
transform 1 0 83040 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_861
timestamp 1677579658
transform 1 0 83232 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_196
timestamp 1677579658
transform 1 0 19392 0 1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_48_201
timestamp 1679577901
transform 1 0 19872 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_205
timestamp 1677579658
transform 1 0 20256 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_211
timestamp 1677579658
transform 1 0 20832 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_266
timestamp 1677580104
transform 1 0 26112 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_335
timestamp 1677579658
transform 1 0 32736 0 1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_48_367
timestamp 1679577901
transform 1 0 35808 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_381
timestamp 1677579658
transform 1 0 37152 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_436
timestamp 1679581782
transform 1 0 42432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_443
timestamp 1679581782
transform 1 0 43104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_450
timestamp 1679581782
transform 1 0 43776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_457
timestamp 1679581782
transform 1 0 44448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_464
timestamp 1679581782
transform 1 0 45120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_471
timestamp 1679581782
transform 1 0 45792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_478
timestamp 1679581782
transform 1 0 46464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_485
timestamp 1679581782
transform 1 0 47136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_492
timestamp 1679581782
transform 1 0 47808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_499
timestamp 1679581782
transform 1 0 48480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_506
timestamp 1679581782
transform 1 0 49152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_513
timestamp 1679581782
transform 1 0 49824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_520
timestamp 1679581782
transform 1 0 50496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_527
timestamp 1679581782
transform 1 0 51168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_534
timestamp 1679581782
transform 1 0 51840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_541
timestamp 1679581782
transform 1 0 52512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_548
timestamp 1679581782
transform 1 0 53184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_555
timestamp 1679581782
transform 1 0 53856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_562
timestamp 1679581782
transform 1 0 54528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_569
timestamp 1679581782
transform 1 0 55200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_576
timestamp 1679581782
transform 1 0 55872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_583
timestamp 1679581782
transform 1 0 56544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_590
timestamp 1679581782
transform 1 0 57216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_597
timestamp 1679581782
transform 1 0 57888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_604
timestamp 1679581782
transform 1 0 58560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_611
timestamp 1679581782
transform 1 0 59232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_618
timestamp 1679581782
transform 1 0 59904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_625
timestamp 1679581782
transform 1 0 60576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_632
timestamp 1679581782
transform 1 0 61248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_639
timestamp 1679581782
transform 1 0 61920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_646
timestamp 1679581782
transform 1 0 62592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_653
timestamp 1679581782
transform 1 0 63264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_660
timestamp 1679581782
transform 1 0 63936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_667
timestamp 1679581782
transform 1 0 64608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_674
timestamp 1679581782
transform 1 0 65280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_681
timestamp 1679581782
transform 1 0 65952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_688
timestamp 1679581782
transform 1 0 66624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_695
timestamp 1679581782
transform 1 0 67296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_702
timestamp 1679581782
transform 1 0 67968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_709
timestamp 1679581782
transform 1 0 68640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_716
timestamp 1679581782
transform 1 0 69312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_723
timestamp 1679581782
transform 1 0 69984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_730
timestamp 1679581782
transform 1 0 70656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_737
timestamp 1679581782
transform 1 0 71328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_744
timestamp 1679581782
transform 1 0 72000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_751
timestamp 1679581782
transform 1 0 72672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_758
timestamp 1679581782
transform 1 0 73344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_765
timestamp 1679581782
transform 1 0 74016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_772
timestamp 1679581782
transform 1 0 74688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_779
timestamp 1679581782
transform 1 0 75360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_786
timestamp 1679581782
transform 1 0 76032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_793
timestamp 1679581782
transform 1 0 76704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_800
timestamp 1679581782
transform 1 0 77376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_807
timestamp 1679581782
transform 1 0 78048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_814
timestamp 1679581782
transform 1 0 78720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_821
timestamp 1679581782
transform 1 0 79392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_828
timestamp 1679581782
transform 1 0 80064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_835
timestamp 1679581782
transform 1 0 80736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_842
timestamp 1679581782
transform 1 0 81408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_849
timestamp 1679581782
transform 1 0 82080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_856
timestamp 1679577901
transform 1 0 82752 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_860
timestamp 1677580104
transform 1 0 83136 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679581782
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679581782
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679581782
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679581782
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679581782
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679581782
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679581782
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679581782
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679581782
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679581782
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679581782
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679581782
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679581782
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_214
timestamp 1679577901
transform 1 0 21120 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_218
timestamp 1677580104
transform 1 0 21504 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_225
timestamp 1677580104
transform 1 0 22176 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_227
timestamp 1677579658
transform 1 0 22368 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_232
timestamp 1679581782
transform 1 0 22848 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_239
timestamp 1677579658
transform 1 0 23520 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679581782
transform 1 0 24768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_259
timestamp 1679577901
transform 1 0 25440 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_263
timestamp 1677579658
transform 1 0 25824 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_267
timestamp 1677580104
transform 1 0 26208 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_4  FILLER_49_273
timestamp 1679577901
transform 1 0 26784 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_277
timestamp 1677580104
transform 1 0 27168 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_285
timestamp 1679581782
transform 1 0 27936 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_292
timestamp 1677580104
transform 1 0 28608 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_294
timestamp 1677579658
transform 1 0 28800 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_307
timestamp 1679581782
transform 1 0 30048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_314
timestamp 1679581782
transform 1 0 30720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_321
timestamp 1679581782
transform 1 0 31392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_328
timestamp 1679581782
transform 1 0 32064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_335
timestamp 1679577901
transform 1 0 32736 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_349
timestamp 1679581782
transform 1 0 34080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_356
timestamp 1679581782
transform 1 0 34752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_363
timestamp 1679581782
transform 1 0 35424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_370
timestamp 1679581782
transform 1 0 36096 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_377
timestamp 1677580104
transform 1 0 36768 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_379
timestamp 1677579658
transform 1 0 36960 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_390
timestamp 1679581782
transform 1 0 38016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_397
timestamp 1679581782
transform 1 0 38688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_404
timestamp 1679581782
transform 1 0 39360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_411
timestamp 1679581782
transform 1 0 40032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_418
timestamp 1679581782
transform 1 0 40704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_425
timestamp 1679581782
transform 1 0 41376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_432
timestamp 1679581782
transform 1 0 42048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_439
timestamp 1679581782
transform 1 0 42720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_446
timestamp 1679581782
transform 1 0 43392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_453
timestamp 1679581782
transform 1 0 44064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_460
timestamp 1679581782
transform 1 0 44736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_467
timestamp 1679581782
transform 1 0 45408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_474
timestamp 1679581782
transform 1 0 46080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_481
timestamp 1679581782
transform 1 0 46752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_488
timestamp 1679581782
transform 1 0 47424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_495
timestamp 1679581782
transform 1 0 48096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_502
timestamp 1679581782
transform 1 0 48768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_509
timestamp 1679581782
transform 1 0 49440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_516
timestamp 1679581782
transform 1 0 50112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_523
timestamp 1679581782
transform 1 0 50784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_530
timestamp 1679581782
transform 1 0 51456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_537
timestamp 1679581782
transform 1 0 52128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_544
timestamp 1679581782
transform 1 0 52800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_551
timestamp 1679581782
transform 1 0 53472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_558
timestamp 1679581782
transform 1 0 54144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_565
timestamp 1679581782
transform 1 0 54816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_572
timestamp 1679581782
transform 1 0 55488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_579
timestamp 1679581782
transform 1 0 56160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_586
timestamp 1679581782
transform 1 0 56832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_593
timestamp 1679581782
transform 1 0 57504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_600
timestamp 1679581782
transform 1 0 58176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_607
timestamp 1679581782
transform 1 0 58848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_614
timestamp 1679581782
transform 1 0 59520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_621
timestamp 1679581782
transform 1 0 60192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_628
timestamp 1679581782
transform 1 0 60864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_635
timestamp 1679581782
transform 1 0 61536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_642
timestamp 1679581782
transform 1 0 62208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_649
timestamp 1679581782
transform 1 0 62880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_656
timestamp 1679581782
transform 1 0 63552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_663
timestamp 1679581782
transform 1 0 64224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_670
timestamp 1679581782
transform 1 0 64896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_677
timestamp 1679581782
transform 1 0 65568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_684
timestamp 1679581782
transform 1 0 66240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_691
timestamp 1679581782
transform 1 0 66912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_698
timestamp 1679581782
transform 1 0 67584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_705
timestamp 1679581782
transform 1 0 68256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_712
timestamp 1679581782
transform 1 0 68928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_719
timestamp 1679581782
transform 1 0 69600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_726
timestamp 1679581782
transform 1 0 70272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_733
timestamp 1679581782
transform 1 0 70944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_740
timestamp 1679581782
transform 1 0 71616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_747
timestamp 1679581782
transform 1 0 72288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_754
timestamp 1679581782
transform 1 0 72960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_761
timestamp 1679581782
transform 1 0 73632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_768
timestamp 1679581782
transform 1 0 74304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_775
timestamp 1679581782
transform 1 0 74976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_782
timestamp 1679581782
transform 1 0 75648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_789
timestamp 1679581782
transform 1 0 76320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_796
timestamp 1679581782
transform 1 0 76992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_803
timestamp 1679581782
transform 1 0 77664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_810
timestamp 1679581782
transform 1 0 78336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_817
timestamp 1679581782
transform 1 0 79008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_824
timestamp 1679581782
transform 1 0 79680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_831
timestamp 1679581782
transform 1 0 80352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_838
timestamp 1679581782
transform 1 0 81024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_845
timestamp 1679581782
transform 1 0 81696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_852
timestamp 1679581782
transform 1 0 82368 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_859
timestamp 1677580104
transform 1 0 83040 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_861
timestamp 1677579658
transform 1 0 83232 0 -1 38556
box -48 -56 144 834
use sg13g2_tielo  heichips25_internal_47
timestamp 1680000637
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_48
timestamp 1680000637
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_49
timestamp 1680000637
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_50
timestamp 1680000637
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_51
timestamp 1680000637
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_52
timestamp 1680000637
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_53
timestamp 1680000637
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal
timestamp 1680000637
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_54
timestamp 1680000637
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_55
timestamp 1680000637
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_56
timestamp 1680000637
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_57
timestamp 1680000637
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_58
timestamp 1680000637
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_59
timestamp 1680000637
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_60
timestamp 1680000637
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  heichips25_internal_61
timestamp 1680000637
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform -1 0 1344 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform -1 0 960 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform -1 0 1344 0 -1 15876
box -48 -56 432 834
use adc  u_adc
timestamp 0
transform 1 0 82800 0 1 1400
box 0 0 1 1
use sg13g2_buf_16  u_clkbuf_analog_pin0.u_buf
timestamp 1676553496
transform -1 0 80736 0 -1 6804
box -48 -56 2448 834
use sg13g2_buf_16  u_clkbuf_analog_pin1.u_buf
timestamp 1676553496
transform -1 0 98976 0 -1 20412
box -48 -56 2448 834
use delay_line  u_delay_line
timestamp 0
transform 1 0 85400 0 1 24600
box 0 0 1 1
use multimode_dll  u_multimode_dll
timestamp 0
transform 1 0 8000 0 1 7400
box 0 0 1 1
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 712 95476 38600 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 99920 33140 100000 33220 0 FreeSans 320 0 0 0 analog_adc
port 2 nsew signal bidirectional
flabel metal3 s 99920 6596 100000 6676 0 FreeSans 320 0 0 0 analog_pin0
port 3 nsew signal bidirectional
flabel metal3 s 99920 19868 100000 19948 0 FreeSans 320 0 0 0 analog_pin1
port 4 nsew signal bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 5 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 6 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 7 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 8 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 9 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 10 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 11 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 12 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 13 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 14 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 15 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 16 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 17 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 18 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 19 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 20 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 21 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 22 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 23 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 24 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 25 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 26 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 27 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 28 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 29 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 30 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 31 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 32 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 33 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 34 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 35 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 36 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 37 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 38 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 39 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 40 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 41 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 42 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 43 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 44 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 45 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 46 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 47 nsew signal output
rlabel via5 65100 24200 65100 24200 0 VGND
rlabel via5 63860 28960 63860 28960 0 VPWR
rlabel metal2 29952 4074 29952 4074 0 _000_
rlabel metal3 21408 37380 21408 37380 0 _001_
rlabel metal2 23472 36876 23472 36876 0 _002_
rlabel metal2 23328 36162 23328 36162 0 _003_
rlabel metal2 26112 36036 26112 36036 0 _004_
rlabel metal2 26880 37884 26880 37884 0 _005_
rlabel metal2 29664 37548 29664 37548 0 _006_
rlabel metal2 30240 37254 30240 37254 0 _007_
rlabel metal2 22944 35196 22944 35196 0 _008_
rlabel metal2 27648 34440 27648 34440 0 _009_
rlabel metal2 30048 34902 30048 34902 0 _010_
rlabel metal2 32160 34440 32160 34440 0 _011_
rlabel metal2 38784 34104 38784 34104 0 _012_
rlabel metal2 43968 34650 43968 34650 0 _013_
rlabel metal2 49584 35280 49584 35280 0 _014_
rlabel metal2 52128 35448 52128 35448 0 _015_
rlabel metal2 52800 33978 52800 33978 0 _016_
rlabel metal2 46944 34902 46944 34902 0 _017_
rlabel metal2 46752 35448 46752 35448 0 _018_
rlabel metal2 32592 36792 32592 36792 0 _019_
rlabel metal3 34848 37968 34848 37968 0 _020_
rlabel metal2 33696 2604 33696 2604 0 _021_
rlabel metal2 36672 2898 36672 2898 0 _022_
rlabel metal2 46032 4116 46032 4116 0 _023_
rlabel metal2 48672 3654 48672 3654 0 _024_
rlabel metal2 51168 3654 51168 3654 0 _025_
rlabel metal2 52704 4116 52704 4116 0 _026_
rlabel metal3 49680 2016 49680 2016 0 _027_
rlabel metal3 48912 1092 48912 1092 0 _028_
rlabel metal2 45216 2394 45216 2394 0 _029_
rlabel metal3 45456 1092 45456 1092 0 _030_
rlabel metal2 41856 1848 41856 1848 0 _031_
rlabel metal3 41568 1092 41568 1092 0 _032_
rlabel metal2 40128 1638 40128 1638 0 _033_
rlabel metal2 37344 1638 37344 1638 0 _034_
rlabel metal2 32256 1638 32256 1638 0 _035_
rlabel metal2 28560 1092 28560 1092 0 _036_
rlabel metal2 26880 1638 26880 1638 0 _037_
rlabel metal3 24960 1764 24960 1764 0 _038_
rlabel metal2 20352 2142 20352 2142 0 _039_
rlabel metal3 21600 3276 21600 3276 0 _040_
rlabel metal2 23328 4116 23328 4116 0 _041_
rlabel metal2 24768 4410 24768 4410 0 _042_
rlabel metal2 26976 3486 26976 3486 0 _043_
rlabel metal2 40512 3360 40512 3360 0 _044_
rlabel metal2 42816 4200 42816 4200 0 _045_
rlabel metal3 45840 3444 45840 3444 0 _046_
rlabel metal2 2976 21042 2976 21042 0 _047_
rlabel metal2 3504 22260 3504 22260 0 _048_
rlabel metal2 4224 23499 4224 23499 0 _049_
rlabel metal3 3840 30492 3840 30492 0 _050_
rlabel metal2 10848 34440 10848 34440 0 _051_
rlabel metal2 13440 34440 13440 34440 0 _052_
rlabel metal2 14976 35112 14976 35112 0 _053_
rlabel metal3 5520 29148 5520 29148 0 _054_
rlabel metal2 3456 9954 3456 9954 0 _055_
rlabel metal2 2496 10710 2496 10710 0 _056_
rlabel metal3 1152 12600 1152 12600 0 _057_
rlabel metal2 1248 13860 1248 13860 0 _058_
rlabel metal3 1200 15372 1200 15372 0 _059_
rlabel metal2 2784 17640 2784 17640 0 _060_
rlabel metal2 3456 18480 3456 18480 0 _061_
rlabel metal2 3504 20076 3504 20076 0 _062_
rlabel metal3 3840 26124 3840 26124 0 _063_
rlabel metal2 16896 35196 16896 35196 0 _064_
rlabel metal2 20736 35448 20736 35448 0 _065_
rlabel metal2 19968 35490 19968 35490 0 _066_
rlabel metal2 16896 4242 16896 4242 0 _067_
rlabel metal2 19200 4872 19200 4872 0 _068_
rlabel metal3 3888 7980 3888 7980 0 _069_
rlabel metal2 3456 11760 3456 11760 0 _070_
rlabel metal2 3456 13032 3456 13032 0 _071_
rlabel metal2 3504 13860 3504 13860 0 _072_
rlabel metal2 4224 15414 4224 15414 0 _073_
rlabel metal2 78192 17052 78192 17052 0 _074_
rlabel metal2 81936 20664 81936 20664 0 _075_
rlabel metal2 80832 28392 80832 28392 0 _076_
rlabel metal2 80256 26250 80256 26250 0 _077_
rlabel metal2 80832 27090 80832 27090 0 _078_
rlabel metal3 79104 28980 79104 28980 0 _079_
rlabel metal2 80544 30576 80544 30576 0 _080_
rlabel metal2 80352 24696 80352 24696 0 _081_
rlabel metal2 80832 24612 80832 24612 0 _082_
rlabel metal3 81120 29232 81120 29232 0 _083_
rlabel metal2 80784 32172 80784 32172 0 _084_
rlabel metal2 80832 33516 80832 33516 0 _085_
rlabel metal2 40896 35112 40896 35112 0 _086_
rlabel metal2 41616 36708 41616 36708 0 _087_
rlabel metal3 41328 36540 41328 36540 0 _088_
rlabel metal2 36288 36981 36288 36981 0 _089_
rlabel metal2 37152 37704 37152 37704 0 _090_
rlabel metal2 36048 35280 36048 35280 0 _091_
rlabel metal3 35520 35280 35520 35280 0 _092_
rlabel metal2 29664 2394 29664 2394 0 _093_
rlabel metal3 19632 36708 19632 36708 0 _094_
rlabel metal2 24480 36834 24480 36834 0 _095_
rlabel metal2 35664 35868 35664 35868 0 _096_
rlabel metal2 36192 5754 36192 5754 0 _097_
rlabel metal2 40128 4326 40128 4326 0 _098_
rlabel metal2 36000 4200 36000 4200 0 _099_
rlabel metal2 39072 3864 39072 3864 0 _100_
rlabel metal3 19008 34734 19008 34734 0 _101_
rlabel metal2 34752 4032 34752 4032 0 _102_
rlabel metal2 34656 4284 34656 4284 0 _103_
rlabel metal2 37632 4326 37632 4326 0 _104_
rlabel metal2 35520 4872 35520 4872 0 _105_
rlabel metal2 32160 3906 32160 3906 0 _106_
rlabel metal2 31872 4620 31872 4620 0 _107_
rlabel metal2 32736 5166 32736 5166 0 _108_
rlabel metal2 32928 4872 32928 4872 0 _109_
rlabel metal2 35040 4872 35040 4872 0 _110_
rlabel metal3 37632 4788 37632 4788 0 _111_
rlabel metal2 21408 35364 21408 35364 0 _112_
rlabel metal3 20112 37464 20112 37464 0 _113_
rlabel metal2 27360 36834 27360 36834 0 _114_
rlabel metal2 27888 36036 27888 36036 0 _115_
rlabel metal2 22560 37115 22560 37115 0 _116_
rlabel via1 21024 35698 21024 35698 0 _117_
rlabel metal2 21984 38388 21984 38388 0 _118_
rlabel metal2 21984 37830 21984 37830 0 _119_
rlabel metal2 24288 36540 24288 36540 0 _120_
rlabel metal2 26400 37044 26400 37044 0 _121_
rlabel metal2 27456 36624 27456 36624 0 _122_
rlabel metal2 27696 36540 27696 36540 0 _123_
rlabel metal2 26640 37632 26640 37632 0 _124_
rlabel metal2 29856 37674 29856 37674 0 _125_
rlabel metal2 36000 36036 36000 36036 0 _126_
rlabel via1 35136 35873 35136 35873 0 _127_
rlabel metal4 98880 8376 98880 8376 0 adc_data\[0\]
rlabel metal2 80928 2688 80928 2688 0 adc_data\[1\]
rlabel metal2 80736 2562 80736 2562 0 adc_data\[2\]
rlabel metal4 36768 2898 36768 2898 0 adc_data\[3\]
rlabel metal2 39264 2520 39264 2520 0 adc_data\[4\]
rlabel metal4 98592 8568 98592 8568 0 adc_data\[5\]
rlabel metal2 37632 5796 37632 5796 0 adc_data\[6\]
rlabel metal2 40704 3024 40704 3024 0 adc_data\[7\]
rlabel metal4 82944 20568 82944 20568 0 analog_adc
rlabel metal3 81456 6636 81456 6636 0 analog_pin0
rlabel metal3 99266 19908 99266 19908 0 analog_pin1
rlabel metal3 3582 36708 3582 36708 0 clk
rlabel metal2 41088 5628 41088 5628 0 clk0_out
rlabel metal2 37920 5964 37920 5964 0 clk1_out
rlabel metal2 37632 7002 37632 7002 0 clk2_out
rlabel metal2 40608 5208 40608 5208 0 clk_delayed
rlabel metal2 44544 5292 44544 5292 0 clk_regs
rlabel metal3 63504 34356 63504 34356 0 clknet_0_clk
rlabel metal2 19584 34398 19584 34398 0 clknet_0_clk_regs
rlabel metal3 26376 7224 26376 7224 0 clknet_1_0__leaf_clk
rlabel metal3 98830 9399 98830 9399 0 clknet_1_1__leaf_clk
rlabel metal2 20448 4536 20448 4536 0 clknet_4_0_0_clk_regs
rlabel metal3 81408 20748 81408 20748 0 clknet_4_10_0_clk_regs
rlabel metal2 62496 34188 62496 34188 0 clknet_4_11_0_clk_regs
rlabel metal3 38592 37338 38592 37338 0 clknet_4_12_0_clk_regs
rlabel metal2 65472 34776 65472 34776 0 clknet_4_13_0_clk_regs
rlabel metal3 62592 34440 62592 34440 0 clknet_4_14_0_clk_regs
rlabel metal2 45504 35154 45504 35154 0 clknet_4_15_0_clk_regs
rlabel metal3 5568 14700 5568 14700 0 clknet_4_1_0_clk_regs
rlabel metal2 26016 3486 26016 3486 0 clknet_4_2_0_clk_regs
rlabel metal2 24672 3024 24672 3024 0 clknet_4_3_0_clk_regs
rlabel metal3 4608 20748 4608 20748 0 clknet_4_4_0_clk_regs
rlabel metal3 9840 34524 9840 34524 0 clknet_4_5_0_clk_regs
rlabel metal2 20544 34776 20544 34776 0 clknet_4_6_0_clk_regs
rlabel metal2 21024 34314 21024 34314 0 clknet_4_7_0_clk_regs
rlabel metal2 45312 1512 45312 1512 0 clknet_4_8_0_clk_regs
rlabel metal2 41760 3780 41760 3780 0 clknet_4_9_0_clk_regs
rlabel metal2 22560 35154 22560 35154 0 data\[0\]
rlabel metal2 44352 35406 44352 35406 0 data\[10\]
rlabel metal2 33696 37968 33696 37968 0 data\[11\]
rlabel metal2 33792 5250 33792 5250 0 data\[12\]
rlabel metal3 34128 3528 34128 3528 0 data\[13\]
rlabel metal2 39072 2940 39072 2940 0 data\[14\]
rlabel metal2 48384 4662 48384 4662 0 data\[15\]
rlabel metal2 47328 5364 47328 5364 0 data\[16\]
rlabel metal2 46944 5448 46944 5448 0 data\[17\]
rlabel metal2 47136 5784 47136 5784 0 data\[18\]
rlabel metal2 47232 1554 47232 1554 0 data\[19\]
rlabel metal2 29773 31573 29773 31573 0 data\[1\]
rlabel metal2 44832 2016 44832 2016 0 data\[20\]
rlabel metal2 43872 2646 43872 2646 0 data\[21\]
rlabel metal3 40944 1932 40944 1932 0 data\[22\]
rlabel metal3 39936 2604 39936 2604 0 data\[23\]
rlabel metal2 40224 2772 40224 2772 0 data\[24\]
rlabel metal3 38160 1680 38160 1680 0 data\[25\]
rlabel metal2 34992 2100 34992 2100 0 data\[26\]
rlabel metal3 35040 2100 35040 2100 0 data\[27\]
rlabel metal2 27072 1008 27072 1008 0 data\[28\]
rlabel metal2 26976 1512 26976 1512 0 data\[29\]
rlabel metal2 32070 31752 32070 31752 0 data\[2\]
rlabel metal2 20736 1890 20736 1890 0 data\[30\]
rlabel metal2 21504 3108 21504 3108 0 data\[31\]
rlabel metal3 22656 3948 22656 3948 0 data\[32\]
rlabel metal2 24816 4956 24816 4956 0 data\[33\]
rlabel metal2 24672 5166 24672 5166 0 data\[34\]
rlabel metal3 41520 3444 41520 3444 0 data\[35\]
rlabel metal2 42240 4074 42240 4074 0 data\[36\]
rlabel metal2 42336 4158 42336 4158 0 data\[37\]
rlabel metal3 4944 21588 4944 21588 0 data\[38\]
rlabel metal2 3360 22050 3360 22050 0 data\[39\]
rlabel metal2 31609 31752 31609 31752 0 data\[3\]
rlabel metal2 5904 22092 5904 22092 0 data\[40\]
rlabel metal3 6880 20916 6880 20916 0 data\[41\]
rlabel metal2 10272 34272 10272 34272 0 data\[42\]
rlabel metal2 18816 32970 18816 32970 0 data\[43\]
rlabel metal2 24006 31752 24006 31752 0 data\[44\]
rlabel metal2 17376 34860 17376 34860 0 data\[45\]
rlabel metal3 4800 11676 4800 11676 0 data\[46\]
rlabel metal2 23808 7086 23808 7086 0 data\[47\]
rlabel metal3 2160 12516 2160 12516 0 data\[48\]
rlabel metal2 1728 12390 1728 12390 0 data\[49\]
rlabel metal2 41184 34020 41184 34020 0 data\[4\]
rlabel metal2 1920 15204 1920 15204 0 data\[50\]
rlabel metal3 3600 16464 3600 16464 0 data\[51\]
rlabel metal2 2880 18228 2880 18228 0 data\[52\]
rlabel metal2 5856 18774 5856 18774 0 data\[53\]
rlabel metal3 5472 19992 5472 19992 0 data\[54\]
rlabel metal2 16333 31447 16333 31447 0 data\[55\]
rlabel metal2 19296 32970 19296 32970 0 data\[56\]
rlabel metal2 23814 31752 23814 31752 0 data\[57\]
rlabel metal2 17472 5838 17472 5838 0 data\[58\]
rlabel metal2 17568 5250 17568 5250 0 data\[59\]
rlabel metal2 46368 34104 46368 34104 0 data\[5\]
rlabel metal2 21600 5376 21600 5376 0 data\[60\]
rlabel metal2 2784 12432 2784 12432 0 data\[61\]
rlabel metal2 5856 12138 5856 12138 0 data\[62\]
rlabel metal3 6928 12684 6928 12684 0 data\[63\]
rlabel metal2 5904 14952 5904 14952 0 data\[64\]
rlabel metal2 5856 16590 5856 16590 0 data\[65\]
rlabel metal3 81936 9240 81936 9240 0 data\[66\]
rlabel metal2 81504 21798 81504 21798 0 data\[67\]
rlabel metal2 83232 28644 83232 28644 0 data\[68\]
rlabel metal2 82704 25956 82704 25956 0 data\[69\]
rlabel metal2 51936 34902 51936 34902 0 data\[6\]
rlabel metal2 83280 27048 83280 27048 0 data\[70\]
rlabel metal3 80928 29652 80928 29652 0 data\[71\]
rlabel metal2 80688 25284 80688 25284 0 data\[72\]
rlabel metal2 82656 24486 82656 24486 0 data\[73\]
rlabel metal2 81504 25368 81504 25368 0 data\[74\]
rlabel metal2 83280 29316 83280 29316 0 data\[75\]
rlabel metal2 83232 31500 83232 31500 0 data\[76\]
rlabel metal3 43968 33894 43968 33894 0 data\[77\]
rlabel metal2 41280 35826 41280 35826 0 data\[78\]
rlabel metal3 42624 35868 42624 35868 0 data\[79\]
rlabel metal3 54192 34944 54192 34944 0 data\[7\]
rlabel metal2 40032 37002 40032 37002 0 data\[80\]
rlabel metal2 38400 37128 38400 37128 0 data\[81\]
rlabel metal2 39744 36540 39744 36540 0 data\[82\]
rlabel metal2 38400 35490 38400 35490 0 data\[83\]
rlabel metal2 30432 2898 30432 2898 0 data\[84\]
rlabel metal3 32304 2100 32304 2100 0 data\[85\]
rlabel metal2 46944 34146 46944 34146 0 data\[8\]
rlabel metal2 46848 34440 46848 34440 0 data\[9\]
rlabel metal3 42528 34440 42528 34440 0 delaynet_0_clk
rlabel metal2 25680 7140 25680 7140 0 ena
rlabel metal3 366 15708 366 15708 0 net
rlabel metal3 3216 37968 3216 37968 0 net1
rlabel metal2 31776 5754 31776 5754 0 net10
rlabel metal2 32784 4788 32784 4788 0 net11
rlabel metal2 912 13944 912 13944 0 net12
rlabel metal4 1248 10248 1248 10248 0 net13
rlabel metal2 2160 18312 2160 18312 0 net14
rlabel metal2 3264 18858 3264 18858 0 net15
rlabel metal2 3984 18732 3984 18732 0 net16
rlabel metal2 3840 21588 3840 21588 0 net17
rlabel via2 19104 35868 19104 35868 0 net18
rlabel via2 27168 2016 27168 2016 0 net19
rlabel metal2 912 23268 912 23268 0 net2
rlabel metal2 38208 1050 38208 1050 0 net20
rlabel metal2 40992 36246 40992 36246 0 net21
rlabel metal2 36288 35280 36288 35280 0 net22
rlabel metal2 22464 4284 22464 4284 0 net23
rlabel metal2 43872 4200 43872 4200 0 net24
rlabel metal2 42432 4662 42432 4662 0 net25
rlabel metal2 80928 23016 80928 23016 0 net26
rlabel metal2 81408 30912 81408 30912 0 net27
rlabel metal2 45600 34272 45600 34272 0 net28
rlabel metal2 22560 37704 22560 37704 0 net29
rlabel metal4 864 29904 864 29904 0 net3
rlabel metal2 3792 13188 3792 13188 0 net30
rlabel metal3 3168 17808 3168 17808 0 net31
rlabel metal2 3024 18312 3024 18312 0 net32
rlabel metal2 3504 20748 3504 20748 0 net33
rlabel metal2 21120 35280 21120 35280 0 net34
rlabel metal2 25728 5166 25728 5166 0 net35
rlabel metal2 26112 3276 26112 3276 0 net36
rlabel metal3 30336 36708 30336 36708 0 net37
rlabel metal2 39168 35196 39168 35196 0 net38
rlabel metal2 41952 36582 41952 36582 0 net39
rlabel metal3 912 24780 912 24780 0 net4
rlabel metal2 26304 5124 26304 5124 0 net40
rlabel metal2 13920 34020 13920 34020 0 net41
rlabel metal2 46368 4158 46368 4158 0 net42
rlabel metal2 44160 34650 44160 34650 0 net43
rlabel metal2 81216 23730 81216 23730 0 net44
rlabel metal2 80928 29904 80928 29904 0 net45
rlabel metal2 43968 35406 43968 35406 0 net46
rlabel metal3 366 16548 366 16548 0 net47
rlabel metal3 366 17388 366 17388 0 net48
rlabel metal3 366 18228 366 18228 0 net49
rlabel metal2 816 25116 816 25116 0 net5
rlabel metal3 366 19068 366 19068 0 net50
rlabel metal3 366 19908 366 19908 0 net51
rlabel metal3 366 20748 366 20748 0 net52
rlabel metal3 366 21588 366 21588 0 net53
rlabel metal3 366 2268 366 2268 0 net54
rlabel metal3 366 3108 366 3108 0 net55
rlabel metal3 366 3948 366 3948 0 net56
rlabel metal3 366 4788 366 4788 0 net57
rlabel metal3 366 5628 366 5628 0 net58
rlabel metal3 366 6468 366 6468 0 net59
rlabel metal4 864 7056 864 7056 0 net6
rlabel metal3 366 7308 366 7308 0 net60
rlabel metal3 318 8148 318 8148 0 net61
rlabel metal3 37440 6426 37440 6426 0 net7
rlabel metal2 49056 5166 49056 5166 0 net8
rlabel metal2 35424 5208 35424 5208 0 net9
rlabel metal2 31968 5700 31968 5700 0 osc_out
rlabel metal3 366 37548 366 37548 0 rst_n
rlabel metal2 34608 5460 34608 5460 0 stable
rlabel metal2 31680 4074 31680 4074 0 u_custom_cells.u_latch0.D
rlabel metal2 33120 4284 33120 4284 0 u_custom_cells.u_latch0.Q
rlabel metal2 22272 36708 22272 36708 0 u_shift_reg.bit_count\[0\]
rlabel metal2 27168 36666 27168 36666 0 u_shift_reg.bit_count\[1\]
rlabel metal2 25728 36498 25728 36498 0 u_shift_reg.bit_count\[2\]
rlabel metal2 27744 36036 27744 36036 0 u_shift_reg.bit_count\[3\]
rlabel metal3 28656 36708 28656 36708 0 u_shift_reg.bit_count\[4\]
rlabel metal2 28992 37338 28992 37338 0 u_shift_reg.bit_count\[5\]
rlabel metal2 29760 37296 29760 37296 0 u_shift_reg.bit_count\[6\]
rlabel metal2 21120 36918 21120 36918 0 u_shift_reg.locked
rlabel metal3 366 22428 366 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 8988 366 8988 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 366 10668 366 10668 0 uio_out[2]
rlabel metal3 366 11508 366 11508 0 uio_out[3]
rlabel metal3 558 12348 558 12348 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 366 14028 366 14028 0 uio_out[6]
rlabel metal3 558 14868 558 14868 0 uio_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
