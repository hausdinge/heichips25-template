module heichips25_internal (analog_adc,
    analog_pin0,
    analog_pin1,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 inout analog_adc;
 inout analog_pin0;
 inout analog_pin1;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire \adc_data[0] ;
 wire \adc_data[1] ;
 wire \adc_data[2] ;
 wire \adc_data[3] ;
 wire \adc_data[4] ;
 wire \adc_data[5] ;
 wire \adc_data[6] ;
 wire \adc_data[7] ;
 wire adc_ready;
 wire clk0_out;
 wire clk1_out;
 wire clk2_out;
 wire clk_delayed;
 wire \data[0] ;
 wire \data[10] ;
 wire \data[11] ;
 wire \data[12] ;
 wire \data[13] ;
 wire \data[14] ;
 wire \data[15] ;
 wire \data[16] ;
 wire \data[17] ;
 wire \data[18] ;
 wire \data[19] ;
 wire \data[1] ;
 wire \data[20] ;
 wire \data[21] ;
 wire \data[22] ;
 wire \data[23] ;
 wire \data[24] ;
 wire \data[25] ;
 wire \data[26] ;
 wire \data[27] ;
 wire \data[28] ;
 wire \data[29] ;
 wire \data[2] ;
 wire \data[30] ;
 wire \data[31] ;
 wire \data[32] ;
 wire \data[33] ;
 wire \data[34] ;
 wire \data[35] ;
 wire \data[36] ;
 wire \data[37] ;
 wire \data[38] ;
 wire \data[39] ;
 wire \data[3] ;
 wire \data[40] ;
 wire \data[41] ;
 wire \data[42] ;
 wire \data[43] ;
 wire \data[44] ;
 wire \data[45] ;
 wire \data[46] ;
 wire \data[47] ;
 wire \data[48] ;
 wire \data[49] ;
 wire \data[4] ;
 wire \data[50] ;
 wire \data[51] ;
 wire \data[52] ;
 wire \data[53] ;
 wire \data[54] ;
 wire \data[55] ;
 wire \data[56] ;
 wire \data[57] ;
 wire \data[58] ;
 wire \data[59] ;
 wire \data[5] ;
 wire \data[60] ;
 wire \data[61] ;
 wire \data[62] ;
 wire \data[63] ;
 wire \data[64] ;
 wire \data[65] ;
 wire \data[66] ;
 wire \data[67] ;
 wire \data[68] ;
 wire \data[69] ;
 wire \data[6] ;
 wire \data[70] ;
 wire \data[71] ;
 wire \data[72] ;
 wire \data[73] ;
 wire \data[74] ;
 wire \data[75] ;
 wire \data[76] ;
 wire \data[77] ;
 wire \data[78] ;
 wire \data[79] ;
 wire \data[7] ;
 wire \data[80] ;
 wire \data[81] ;
 wire \data[82] ;
 wire \data[83] ;
 wire \data[84] ;
 wire \data[85] ;
 wire \data[8] ;
 wire \data[9] ;
 wire osc_out;
 wire net1;
 wire stable;
 wire \u_custom_cells.u_latch0.D ;
 wire \u_custom_cells.u_latch0.Q ;
 wire \u_shift_reg.bit_count[0] ;
 wire \u_shift_reg.bit_count[1] ;
 wire \u_shift_reg.bit_count[2] ;
 wire \u_shift_reg.bit_count[3] ;
 wire \u_shift_reg.bit_count[4] ;
 wire \u_shift_reg.bit_count[5] ;
 wire \u_shift_reg.bit_count[6] ;
 wire \u_shift_reg.locked ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire clk_regs;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;

 sg13g2_inv_1 _128_ (.Y(_095_),
    .A(\u_shift_reg.bit_count[2] ));
 sg13g2_inv_1 _129_ (.Y(_096_),
    .A(\data[83] ));
 sg13g2_mux2_1 _130_ (.A0(\data[80] ),
    .A1(\data[81] ),
    .S(\data[82] ),
    .X(_097_));
 sg13g2_mux2_1 _131_ (.A0(\data[78] ),
    .A1(\data[79] ),
    .S(\data[82] ),
    .X(_098_));
 sg13g2_nor2_1 _132_ (.A(\data[83] ),
    .B(_098_),
    .Y(_099_));
 sg13g2_a21oi_1 _133_ (.A1(\data[83] ),
    .A2(_097_),
    .Y(_000_),
    .B1(_099_));
 sg13g2_nor2b_1 _134_ (.A(net5),
    .B_N(net4),
    .Y(_100_));
 sg13g2_and2_1 _135_ (.A(\adc_data[0] ),
    .B(_100_),
    .X(net6));
 sg13g2_and2_1 _136_ (.A(\adc_data[1] ),
    .B(_100_),
    .X(net7));
 sg13g2_and2_1 _137_ (.A(\adc_data[2] ),
    .B(_100_),
    .X(net8));
 sg13g2_nor2_1 _138_ (.A(_096_),
    .B(_098_),
    .Y(_101_));
 sg13g2_and2_1 _139_ (.A(net5),
    .B(net4),
    .X(_102_));
 sg13g2_o21ai_1 _140_ (.B1(_102_),
    .Y(_103_),
    .A1(\data[83] ),
    .A2(\u_custom_cells.u_latch0.Q ));
 sg13g2_nor2_1 _141_ (.A(net5),
    .B(net4),
    .Y(_104_));
 sg13g2_a22oi_1 _142_ (.Y(_105_),
    .B1(_104_),
    .B2(stable),
    .A2(_100_),
    .A1(\adc_data[3] ));
 sg13g2_o21ai_1 _143_ (.B1(_105_),
    .Y(net9),
    .A1(_101_),
    .A2(_103_));
 sg13g2_nand2_1 _144_ (.Y(_106_),
    .A(\adc_data[4] ),
    .B(_100_));
 sg13g2_a22oi_1 _145_ (.Y(_107_),
    .B1(_104_),
    .B2(osc_out),
    .A2(_102_),
    .A1(\u_custom_cells.u_latch0.D ));
 sg13g2_nand2_1 _146_ (.Y(net10),
    .A(_106_),
    .B(_107_));
 sg13g2_nand2_1 _147_ (.Y(_108_),
    .A(\adc_data[5] ),
    .B(_100_));
 sg13g2_a22oi_1 _148_ (.Y(_109_),
    .B1(_104_),
    .B2(clk2_out),
    .A2(_102_),
    .A1(\u_custom_cells.u_latch0.Q ));
 sg13g2_nand2_1 _149_ (.Y(net11),
    .A(_108_),
    .B(_109_));
 sg13g2_nand2b_1 _150_ (.Y(_110_),
    .B(_102_),
    .A_N(_097_));
 sg13g2_a22oi_1 _151_ (.Y(_111_),
    .B1(_104_),
    .B2(clk1_out),
    .A2(_100_),
    .A1(\adc_data[6] ));
 sg13g2_nand2_1 _152_ (.Y(net12),
    .A(_110_),
    .B(_111_));
 sg13g2_mux4_1 _153_ (.S0(net4),
    .A0(clk0_out),
    .A1(\adc_data[7] ),
    .A2(clk_delayed),
    .A3(_098_),
    .S1(net5),
    .X(net13));
 sg13g2_nor2b_1 _154_ (.A(\u_shift_reg.locked ),
    .B_N(net2),
    .Y(_112_));
 sg13g2_nand2b_1 _155_ (.Y(_113_),
    .B(net2),
    .A_N(\u_shift_reg.locked ));
 sg13g2_and2_1 _156_ (.A(\u_shift_reg.bit_count[0] ),
    .B(\u_shift_reg.bit_count[2] ),
    .X(_114_));
 sg13g2_nor3_1 _157_ (.A(\u_shift_reg.bit_count[1] ),
    .B(\u_shift_reg.bit_count[3] ),
    .C(\u_shift_reg.bit_count[5] ),
    .Y(_115_));
 sg13g2_nand4_1 _158_ (.B(\u_shift_reg.bit_count[6] ),
    .C(_114_),
    .A(\u_shift_reg.bit_count[4] ),
    .Y(_116_),
    .D(_115_));
 sg13g2_inv_1 _159_ (.Y(_117_),
    .A(_116_));
 sg13g2_nand3_1 _160_ (.B(net29),
    .C(_116_),
    .A(\u_shift_reg.bit_count[0] ),
    .Y(_118_));
 sg13g2_a21o_1 _161_ (.A2(_116_),
    .A1(net29),
    .B1(\u_shift_reg.bit_count[0] ),
    .X(_119_));
 sg13g2_and2_1 _162_ (.A(_118_),
    .B(_119_),
    .X(_001_));
 sg13g2_nand3_1 _163_ (.B(\u_shift_reg.bit_count[1] ),
    .C(net29),
    .A(\u_shift_reg.bit_count[0] ),
    .Y(_120_));
 sg13g2_xnor2_1 _164_ (.Y(_002_),
    .A(\u_shift_reg.bit_count[1] ),
    .B(_118_));
 sg13g2_and3_1 _165_ (.X(_121_),
    .A(\u_shift_reg.bit_count[1] ),
    .B(net29),
    .C(_114_));
 sg13g2_a21oi_1 _166_ (.A1(_095_),
    .A2(_120_),
    .Y(_003_),
    .B1(_121_));
 sg13g2_xor2_1 _167_ (.B(_121_),
    .A(\u_shift_reg.bit_count[3] ),
    .X(_004_));
 sg13g2_and2_1 _168_ (.A(\u_shift_reg.bit_count[3] ),
    .B(\u_shift_reg.bit_count[4] ),
    .X(_122_));
 sg13g2_and4_1 _169_ (.A(\u_shift_reg.bit_count[1] ),
    .B(net29),
    .C(_114_),
    .D(_122_),
    .X(_123_));
 sg13g2_a21oi_1 _170_ (.A1(\u_shift_reg.bit_count[3] ),
    .A2(_121_),
    .Y(_124_),
    .B1(\u_shift_reg.bit_count[4] ));
 sg13g2_nor2_1 _171_ (.A(_123_),
    .B(_124_),
    .Y(_005_));
 sg13g2_nand2_1 _172_ (.Y(_125_),
    .A(\u_shift_reg.bit_count[5] ),
    .B(_123_));
 sg13g2_xor2_1 _173_ (.B(_123_),
    .A(\u_shift_reg.bit_count[5] ),
    .X(_006_));
 sg13g2_xnor2_1 _174_ (.Y(_007_),
    .A(\u_shift_reg.bit_count[6] ),
    .B(_125_));
 sg13g2_mux2_1 _175_ (.A0(\data[0] ),
    .A1(net3),
    .S(net29),
    .X(_008_));
 sg13g2_mux2_1 _176_ (.A0(\data[0] ),
    .A1(\data[1] ),
    .S(net22),
    .X(_009_));
 sg13g2_mux2_1 _177_ (.A0(\data[1] ),
    .A1(\data[2] ),
    .S(net22),
    .X(_010_));
 sg13g2_mux2_1 _178_ (.A0(\data[2] ),
    .A1(\data[3] ),
    .S(net21),
    .X(_011_));
 sg13g2_mux2_1 _179_ (.A0(\data[3] ),
    .A1(\data[4] ),
    .S(net21),
    .X(_012_));
 sg13g2_mux2_1 _180_ (.A0(\data[4] ),
    .A1(\data[5] ),
    .S(net25),
    .X(_013_));
 sg13g2_mux2_1 _181_ (.A0(\data[5] ),
    .A1(\data[6] ),
    .S(net25),
    .X(_014_));
 sg13g2_mux2_1 _182_ (.A0(\data[6] ),
    .A1(\data[7] ),
    .S(net25),
    .X(_015_));
 sg13g2_mux2_1 _183_ (.A0(\data[7] ),
    .A1(\data[8] ),
    .S(net25),
    .X(_016_));
 sg13g2_mux2_1 _184_ (.A0(\data[8] ),
    .A1(\data[9] ),
    .S(net25),
    .X(_017_));
 sg13g2_mux2_1 _185_ (.A0(\data[9] ),
    .A1(\data[10] ),
    .S(net28),
    .X(_018_));
 sg13g2_mux2_1 _186_ (.A0(\data[10] ),
    .A1(\data[11] ),
    .S(net21),
    .X(_019_));
 sg13g2_mux2_1 _187_ (.A0(\data[11] ),
    .A1(\data[12] ),
    .S(net21),
    .X(_020_));
 sg13g2_mux2_1 _188_ (.A0(\data[12] ),
    .A1(\data[13] ),
    .S(net19),
    .X(_021_));
 sg13g2_mux2_1 _189_ (.A0(\data[13] ),
    .A1(\data[14] ),
    .S(net20),
    .X(_022_));
 sg13g2_mux2_1 _190_ (.A0(\data[14] ),
    .A1(\data[15] ),
    .S(net24),
    .X(_023_));
 sg13g2_mux2_1 _191_ (.A0(\data[15] ),
    .A1(\data[16] ),
    .S(net24),
    .X(_024_));
 sg13g2_mux2_1 _192_ (.A0(\data[16] ),
    .A1(\data[17] ),
    .S(net24),
    .X(_025_));
 sg13g2_mux2_1 _193_ (.A0(\data[17] ),
    .A1(\data[18] ),
    .S(net25),
    .X(_026_));
 sg13g2_mux2_1 _194_ (.A0(\data[18] ),
    .A1(\data[19] ),
    .S(net24),
    .X(_027_));
 sg13g2_mux2_1 _195_ (.A0(\data[19] ),
    .A1(\data[20] ),
    .S(net25),
    .X(_028_));
 sg13g2_mux2_1 _196_ (.A0(\data[20] ),
    .A1(\data[21] ),
    .S(net24),
    .X(_029_));
 sg13g2_mux2_1 _197_ (.A0(\data[21] ),
    .A1(\data[22] ),
    .S(net24),
    .X(_030_));
 sg13g2_mux2_1 _198_ (.A0(\data[22] ),
    .A1(\data[23] ),
    .S(net20),
    .X(_031_));
 sg13g2_mux2_1 _199_ (.A0(\data[23] ),
    .A1(\data[24] ),
    .S(net20),
    .X(_032_));
 sg13g2_mux2_1 _200_ (.A0(\data[24] ),
    .A1(\data[25] ),
    .S(net20),
    .X(_033_));
 sg13g2_mux2_1 _201_ (.A0(\data[25] ),
    .A1(\data[26] ),
    .S(net20),
    .X(_034_));
 sg13g2_mux2_1 _202_ (.A0(\data[26] ),
    .A1(\data[27] ),
    .S(net20),
    .X(_035_));
 sg13g2_mux2_1 _203_ (.A0(\data[27] ),
    .A1(\data[28] ),
    .S(net19),
    .X(_036_));
 sg13g2_mux2_1 _204_ (.A0(\data[28] ),
    .A1(\data[29] ),
    .S(net19),
    .X(_037_));
 sg13g2_mux2_1 _205_ (.A0(\data[29] ),
    .A1(\data[30] ),
    .S(net19),
    .X(_038_));
 sg13g2_mux2_1 _206_ (.A0(\data[30] ),
    .A1(\data[31] ),
    .S(net16),
    .X(_039_));
 sg13g2_mux2_1 _207_ (.A0(\data[31] ),
    .A1(\data[32] ),
    .S(net16),
    .X(_040_));
 sg13g2_mux2_1 _208_ (.A0(\data[32] ),
    .A1(\data[33] ),
    .S(net19),
    .X(_041_));
 sg13g2_mux2_1 _209_ (.A0(\data[33] ),
    .A1(\data[34] ),
    .S(net19),
    .X(_042_));
 sg13g2_mux2_1 _210_ (.A0(\data[34] ),
    .A1(\data[35] ),
    .S(net19),
    .X(_043_));
 sg13g2_mux2_1 _211_ (.A0(\data[35] ),
    .A1(\data[36] ),
    .S(net20),
    .X(_044_));
 sg13g2_mux2_1 _212_ (.A0(\data[36] ),
    .A1(\data[37] ),
    .S(net24),
    .X(_045_));
 sg13g2_mux2_1 _213_ (.A0(\data[37] ),
    .A1(\data[38] ),
    .S(net24),
    .X(_046_));
 sg13g2_mux2_1 _214_ (.A0(\data[38] ),
    .A1(\data[39] ),
    .S(net17),
    .X(_047_));
 sg13g2_mux2_1 _215_ (.A0(\data[39] ),
    .A1(\data[40] ),
    .S(net17),
    .X(_048_));
 sg13g2_mux2_1 _216_ (.A0(\data[40] ),
    .A1(\data[41] ),
    .S(net17),
    .X(_049_));
 sg13g2_mux2_1 _217_ (.A0(\data[41] ),
    .A1(\data[42] ),
    .S(net17),
    .X(_050_));
 sg13g2_mux2_1 _218_ (.A0(\data[42] ),
    .A1(\data[43] ),
    .S(net17),
    .X(_051_));
 sg13g2_mux2_1 _219_ (.A0(\data[43] ),
    .A1(\data[44] ),
    .S(net18),
    .X(_052_));
 sg13g2_mux2_1 _220_ (.A0(\data[44] ),
    .A1(\data[45] ),
    .S(net18),
    .X(_053_));
 sg13g2_mux2_1 _221_ (.A0(\data[45] ),
    .A1(\data[46] ),
    .S(net17),
    .X(_054_));
 sg13g2_mux2_1 _222_ (.A0(\data[46] ),
    .A1(\data[47] ),
    .S(net15),
    .X(_055_));
 sg13g2_mux2_1 _223_ (.A0(\data[47] ),
    .A1(\data[48] ),
    .S(net15),
    .X(_056_));
 sg13g2_mux2_1 _224_ (.A0(\data[48] ),
    .A1(\data[49] ),
    .S(net14),
    .X(_057_));
 sg13g2_mux2_1 _225_ (.A0(\data[49] ),
    .A1(\data[50] ),
    .S(net14),
    .X(_058_));
 sg13g2_mux2_1 _226_ (.A0(\data[50] ),
    .A1(\data[51] ),
    .S(net14),
    .X(_059_));
 sg13g2_mux2_1 _227_ (.A0(\data[51] ),
    .A1(\data[52] ),
    .S(net14),
    .X(_060_));
 sg13g2_mux2_1 _228_ (.A0(\data[52] ),
    .A1(\data[53] ),
    .S(net14),
    .X(_061_));
 sg13g2_mux2_1 _229_ (.A0(\data[53] ),
    .A1(\data[54] ),
    .S(net17),
    .X(_062_));
 sg13g2_mux2_1 _230_ (.A0(\data[54] ),
    .A1(\data[55] ),
    .S(net17),
    .X(_063_));
 sg13g2_mux2_1 _231_ (.A0(\data[55] ),
    .A1(\data[56] ),
    .S(net18),
    .X(_064_));
 sg13g2_mux2_1 _232_ (.A0(\data[56] ),
    .A1(\data[57] ),
    .S(net18),
    .X(_065_));
 sg13g2_mux2_1 _233_ (.A0(\data[57] ),
    .A1(\data[58] ),
    .S(net18),
    .X(_066_));
 sg13g2_mux2_1 _234_ (.A0(\data[58] ),
    .A1(\data[59] ),
    .S(net16),
    .X(_067_));
 sg13g2_mux2_1 _235_ (.A0(\data[59] ),
    .A1(\data[60] ),
    .S(net16),
    .X(_068_));
 sg13g2_mux2_1 _236_ (.A0(\data[60] ),
    .A1(\data[61] ),
    .S(net15),
    .X(_069_));
 sg13g2_mux2_1 _237_ (.A0(\data[61] ),
    .A1(\data[62] ),
    .S(net14),
    .X(_070_));
 sg13g2_mux2_1 _238_ (.A0(\data[62] ),
    .A1(\data[63] ),
    .S(net14),
    .X(_071_));
 sg13g2_mux2_1 _239_ (.A0(\data[63] ),
    .A1(\data[64] ),
    .S(net14),
    .X(_072_));
 sg13g2_mux2_1 _240_ (.A0(\data[64] ),
    .A1(\data[65] ),
    .S(net15),
    .X(_073_));
 sg13g2_mux2_1 _241_ (.A0(\data[65] ),
    .A1(\data[66] ),
    .S(net28),
    .X(_074_));
 sg13g2_mux2_1 _242_ (.A0(\data[66] ),
    .A1(\data[67] ),
    .S(net26),
    .X(_075_));
 sg13g2_mux2_1 _243_ (.A0(\data[67] ),
    .A1(\data[68] ),
    .S(net26),
    .X(_076_));
 sg13g2_mux2_1 _244_ (.A0(\data[68] ),
    .A1(\data[69] ),
    .S(net26),
    .X(_077_));
 sg13g2_mux2_1 _245_ (.A0(\data[69] ),
    .A1(\data[70] ),
    .S(net26),
    .X(_078_));
 sg13g2_mux2_1 _246_ (.A0(\data[70] ),
    .A1(\data[71] ),
    .S(net26),
    .X(_079_));
 sg13g2_mux2_1 _247_ (.A0(\data[71] ),
    .A1(\data[72] ),
    .S(net26),
    .X(_080_));
 sg13g2_mux2_1 _248_ (.A0(\data[72] ),
    .A1(\data[73] ),
    .S(net26),
    .X(_081_));
 sg13g2_mux2_1 _249_ (.A0(\data[73] ),
    .A1(\data[74] ),
    .S(net26),
    .X(_082_));
 sg13g2_mux2_1 _250_ (.A0(\data[74] ),
    .A1(\data[75] ),
    .S(net27),
    .X(_083_));
 sg13g2_mux2_1 _251_ (.A0(\data[75] ),
    .A1(\data[76] ),
    .S(net27),
    .X(_084_));
 sg13g2_mux2_1 _252_ (.A0(\data[76] ),
    .A1(\data[77] ),
    .S(net27),
    .X(_085_));
 sg13g2_mux2_1 _253_ (.A0(\data[78] ),
    .A1(\data[77] ),
    .S(net29),
    .X(_086_));
 sg13g2_mux2_1 _254_ (.A0(\data[78] ),
    .A1(\data[79] ),
    .S(net21),
    .X(_087_));
 sg13g2_mux2_1 _255_ (.A0(\data[79] ),
    .A1(\data[80] ),
    .S(net21),
    .X(_088_));
 sg13g2_mux2_1 _256_ (.A0(\data[80] ),
    .A1(\data[81] ),
    .S(net21),
    .X(_089_));
 sg13g2_mux2_1 _257_ (.A0(\data[82] ),
    .A1(\data[81] ),
    .S(net29),
    .X(_090_));
 sg13g2_nor2_1 _258_ (.A(\data[82] ),
    .B(net21),
    .Y(_126_));
 sg13g2_a21oi_1 _259_ (.A1(_096_),
    .A2(net22),
    .Y(_091_),
    .B1(_126_));
 sg13g2_nor2_1 _260_ (.A(\data[84] ),
    .B(_112_),
    .Y(_127_));
 sg13g2_a21oi_1 _261_ (.A1(_096_),
    .A2(_112_),
    .Y(_092_),
    .B1(_127_));
 sg13g2_mux2_1 _262_ (.A0(\data[84] ),
    .A1(\data[85] ),
    .S(net19),
    .X(_093_));
 sg13g2_a21o_1 _263_ (.A2(_117_),
    .A1(net2),
    .B1(\u_shift_reg.locked ),
    .X(_094_));
 sg13g2_dfrbpq_1 _264_ (.RESET_B(net34),
    .D(_001_),
    .Q(\u_shift_reg.bit_count[0] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _265_ (.RESET_B(net37),
    .D(_002_),
    .Q(\u_shift_reg.bit_count[1] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _266_ (.RESET_B(net37),
    .D(_003_),
    .Q(\u_shift_reg.bit_count[2] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _267_ (.RESET_B(net37),
    .D(_004_),
    .Q(\u_shift_reg.bit_count[3] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _268_ (.RESET_B(net37),
    .D(_005_),
    .Q(\u_shift_reg.bit_count[4] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _269_ (.RESET_B(net37),
    .D(_006_),
    .Q(\u_shift_reg.bit_count[5] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _270_ (.RESET_B(net37),
    .D(_007_),
    .Q(\u_shift_reg.bit_count[6] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _271_ (.RESET_B(net37),
    .D(_008_),
    .Q(\data[0] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _272_ (.RESET_B(net37),
    .D(_009_),
    .Q(\data[1] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _273_ (.RESET_B(net39),
    .D(_010_),
    .Q(\data[2] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _274_ (.RESET_B(net39),
    .D(_011_),
    .Q(\data[3] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _275_ (.RESET_B(net38),
    .D(_012_),
    .Q(\data[4] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _276_ (.RESET_B(net43),
    .D(_013_),
    .Q(\data[5] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _277_ (.RESET_B(net43),
    .D(_014_),
    .Q(\data[6] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _278_ (.RESET_B(net43),
    .D(_015_),
    .Q(\data[7] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _279_ (.RESET_B(net43),
    .D(_016_),
    .Q(\data[8] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _280_ (.RESET_B(net43),
    .D(_017_),
    .Q(\data[9] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _281_ (.RESET_B(net43),
    .D(_018_),
    .Q(\data[10] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _282_ (.RESET_B(net38),
    .D(_019_),
    .Q(\data[11] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _283_ (.RESET_B(net38),
    .D(_020_),
    .Q(\data[12] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _284_ (.RESET_B(net36),
    .D(_021_),
    .Q(\data[13] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _285_ (.RESET_B(net36),
    .D(_022_),
    .Q(\data[14] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _286_ (.RESET_B(net42),
    .D(_023_),
    .Q(\data[15] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _287_ (.RESET_B(net42),
    .D(_024_),
    .Q(\data[16] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _288_ (.RESET_B(net42),
    .D(_025_),
    .Q(\data[17] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _289_ (.RESET_B(net42),
    .D(_026_),
    .Q(\data[18] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _290_ (.RESET_B(net43),
    .D(_027_),
    .Q(\data[19] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _291_ (.RESET_B(net42),
    .D(_028_),
    .Q(\data[20] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _292_ (.RESET_B(net42),
    .D(_029_),
    .Q(\data[21] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _293_ (.RESET_B(net42),
    .D(_030_),
    .Q(\data[22] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _294_ (.RESET_B(net36),
    .D(_031_),
    .Q(\data[23] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _295_ (.RESET_B(net36),
    .D(_032_),
    .Q(\data[24] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _296_ (.RESET_B(net36),
    .D(_033_),
    .Q(\data[25] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _297_ (.RESET_B(net36),
    .D(_034_),
    .Q(\data[26] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _298_ (.RESET_B(net35),
    .D(_035_),
    .Q(\data[27] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _299_ (.RESET_B(net35),
    .D(_036_),
    .Q(\data[28] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _300_ (.RESET_B(net35),
    .D(_037_),
    .Q(\data[29] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _301_ (.RESET_B(net35),
    .D(_038_),
    .Q(\data[30] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _302_ (.RESET_B(net32),
    .D(_039_),
    .Q(\data[31] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _303_ (.RESET_B(net32),
    .D(_040_),
    .Q(\data[32] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _304_ (.RESET_B(net35),
    .D(_041_),
    .Q(\data[33] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _305_ (.RESET_B(net35),
    .D(_042_),
    .Q(\data[34] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _306_ (.RESET_B(net35),
    .D(_043_),
    .Q(\data[35] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _307_ (.RESET_B(net40),
    .D(_044_),
    .Q(\data[36] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _308_ (.RESET_B(net40),
    .D(_045_),
    .Q(\data[37] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _309_ (.RESET_B(net42),
    .D(_046_),
    .Q(\data[38] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _310_ (.RESET_B(net33),
    .D(_047_),
    .Q(\data[39] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _311_ (.RESET_B(net33),
    .D(_048_),
    .Q(\data[40] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _312_ (.RESET_B(net33),
    .D(_049_),
    .Q(\data[41] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _313_ (.RESET_B(net33),
    .D(_050_),
    .Q(\data[42] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _314_ (.RESET_B(net33),
    .D(_051_),
    .Q(\data[43] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _315_ (.RESET_B(net34),
    .D(_052_),
    .Q(\data[44] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _316_ (.RESET_B(net34),
    .D(_053_),
    .Q(\data[45] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _317_ (.RESET_B(net33),
    .D(_054_),
    .Q(\data[46] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _318_ (.RESET_B(net31),
    .D(_055_),
    .Q(\data[47] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _319_ (.RESET_B(net30),
    .D(_056_),
    .Q(\data[48] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _320_ (.RESET_B(net30),
    .D(_057_),
    .Q(\data[49] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _321_ (.RESET_B(net30),
    .D(_058_),
    .Q(\data[50] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _322_ (.RESET_B(net30),
    .D(_059_),
    .Q(\data[51] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _323_ (.RESET_B(net30),
    .D(_060_),
    .Q(\data[52] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _324_ (.RESET_B(net31),
    .D(_061_),
    .Q(\data[53] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _325_ (.RESET_B(net33),
    .D(_062_),
    .Q(\data[54] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _326_ (.RESET_B(net33),
    .D(_063_),
    .Q(\data[55] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _327_ (.RESET_B(net34),
    .D(_064_),
    .Q(\data[56] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _328_ (.RESET_B(net34),
    .D(_065_),
    .Q(\data[57] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _329_ (.RESET_B(net34),
    .D(_066_),
    .Q(\data[58] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _330_ (.RESET_B(net32),
    .D(_067_),
    .Q(\data[59] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _331_ (.RESET_B(net32),
    .D(_068_),
    .Q(\data[60] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _332_ (.RESET_B(net31),
    .D(_069_),
    .Q(\data[61] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _333_ (.RESET_B(net30),
    .D(_070_),
    .Q(\data[62] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _334_ (.RESET_B(net30),
    .D(_071_),
    .Q(\data[63] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _335_ (.RESET_B(net30),
    .D(_072_),
    .Q(\data[64] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _336_ (.RESET_B(net31),
    .D(_073_),
    .Q(\data[65] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _337_ (.RESET_B(net46),
    .D(_074_),
    .Q(\data[66] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _338_ (.RESET_B(net44),
    .D(_075_),
    .Q(\data[67] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _339_ (.RESET_B(net44),
    .D(_076_),
    .Q(\data[68] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _340_ (.RESET_B(net44),
    .D(_077_),
    .Q(\data[69] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _341_ (.RESET_B(net44),
    .D(_078_),
    .Q(\data[70] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_1 _342_ (.RESET_B(net44),
    .D(_079_),
    .Q(\data[71] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _343_ (.RESET_B(net45),
    .D(_080_),
    .Q(\data[72] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _344_ (.RESET_B(net44),
    .D(_081_),
    .Q(\data[73] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _345_ (.RESET_B(net44),
    .D(_082_),
    .Q(\data[74] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _346_ (.RESET_B(net45),
    .D(_083_),
    .Q(\data[75] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _347_ (.RESET_B(net45),
    .D(_084_),
    .Q(\data[76] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _348_ (.RESET_B(net45),
    .D(_085_),
    .Q(\data[77] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _349_ (.RESET_B(net38),
    .D(_086_),
    .Q(\data[78] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _350_ (.RESET_B(net39),
    .D(_087_),
    .Q(\data[79] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _351_ (.RESET_B(net39),
    .D(_088_),
    .Q(\data[80] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _352_ (.RESET_B(net38),
    .D(_089_),
    .Q(\data[81] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _353_ (.RESET_B(net38),
    .D(_090_),
    .Q(\data[82] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _354_ (.RESET_B(net38),
    .D(_091_),
    .Q(\data[83] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _355_ (.RESET_B(net38),
    .D(_092_),
    .Q(\data[84] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _356_ (.RESET_B(net36),
    .D(_093_),
    .Q(\data[85] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _357_ (.RESET_B(net34),
    .D(_094_),
    .Q(\u_shift_reg.locked ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dlhq_1 _358_ (.D(_000_),
    .GATE(\data[84] ),
    .Q(\u_custom_cells.u_latch0.D ));
 sg13g2_dlhq_1 _359_ (.D(\u_custom_cells.u_latch0.D ),
    .GATE(\data[85] ),
    .Q(\u_custom_cells.u_latch0.Q ));
 sg13g2_tielo heichips25_internal_47 (.L_LO(net47));
 sg13g2_tielo heichips25_internal_48 (.L_LO(net48));
 sg13g2_tielo heichips25_internal_49 (.L_LO(net49));
 sg13g2_tielo heichips25_internal_50 (.L_LO(net50));
 sg13g2_tielo heichips25_internal_51 (.L_LO(net51));
 sg13g2_tielo heichips25_internal_52 (.L_LO(net52));
 sg13g2_tielo heichips25_internal_53 (.L_LO(net53));
 sg13g2_tielo heichips25_internal_54 (.L_LO(net54));
 sg13g2_tielo heichips25_internal_55 (.L_LO(net55));
 sg13g2_tielo heichips25_internal_56 (.L_LO(net56));
 sg13g2_tielo heichips25_internal_57 (.L_LO(net57));
 sg13g2_tielo heichips25_internal_58 (.L_LO(net58));
 sg13g2_tielo heichips25_internal_59 (.L_LO(net59));
 sg13g2_tielo heichips25_internal_60 (.L_LO(net60));
 sg13g2_tielo heichips25_internal_61 (.L_LO(net61));
 sg13g2_buf_16 clkbuf_regs_0_clk (.X(clk_regs),
    .A(clk));
 adc u_adc (.analog_in(analog_adc),
    .clk(clknet_1_1__leaf_clk),
    .ready(adc_ready),
    .start(\data[66] ),
    .data_out({\adc_data[7] ,
    \adc_data[6] ,
    \adc_data[5] ,
    \adc_data[4] ,
    \adc_data[3] ,
    \adc_data[2] ,
    \adc_data[1] ,
    \adc_data[0] }));
 sg13g2_buf_16 \u_clkbuf_analog_pin0.u_buf  (.X(analog_pin0),
    .A(clk0_out));
 sg13g2_buf_16 \u_clkbuf_analog_pin1.u_buf  (.X(analog_pin1),
    .A(clk1_out));
 delay_line u_delay_line (.clk(clknet_1_0__leaf_clk),
    .clk_delayed(clk_delayed),
    .reset(net44),
    .sel({\data[77] ,
    \data[76] ,
    \data[75] }),
    .trim({\data[74] ,
    \data[73] ,
    \data[72] ,
    \data[71] ,
    \data[70] ,
    \data[69] ,
    \data[68] ,
    \data[67] }));
 multimode_dll u_multimode_dll (.bias(\data[38] ),
    .clk0_out(clk0_out),
    .clk1_out(clk1_out),
    .clk2_out(clk2_out),
    .dco(\data[39] ),
    .enable(ena),
    .osc(clknet_1_0__leaf_clk),
    .osc_out(osc_out),
    .resetb(net35),
    .stable(stable),
    .clk0_phase_sel({\data[24] ,
    \data[23] ,
    \data[22] ,
    \data[21] ,
    \data[20] }),
    .clk1_phase_sel({\data[29] ,
    \data[28] ,
    \data[27] ,
    \data[26] ,
    \data[25] }),
    .clk2_phase_sel({\data[34] ,
    \data[33] ,
    \data[32] ,
    \data[31] ,
    \data[30] }),
    .ext_trim({\data[65] ,
    \data[64] ,
    \data[63] ,
    \data[62] ,
    \data[61] ,
    \data[60] ,
    \data[59] ,
    \data[58] ,
    \data[57] ,
    \data[56] ,
    \data[55] ,
    \data[54] ,
    \data[53] ,
    \data[52] ,
    \data[51] ,
    \data[50] ,
    \data[49] ,
    \data[48] ,
    \data[47] ,
    \data[46] ,
    \data[45] ,
    \data[44] ,
    \data[43] ,
    \data[42] ,
    \data[41] ,
    \data[40] }),
    .f_clk0_divider({\data[9] ,
    \data[8] ,
    \data[7] ,
    \data[6] ,
    \data[5] }),
    .f_clk1_divider({\data[14] ,
    \data[13] ,
    \data[12] ,
    \data[11] ,
    \data[10] }),
    .f_clk2_divider({\data[19] ,
    \data[18] ,
    \data[17] ,
    \data[16] ,
    \data[15] }),
    .f_osc_multiply_factor({\data[4] ,
    \data[3] ,
    \data[2] ,
    \data[1] ,
    \data[0] }),
    .mode_xor({\data[37] ,
    \data[36] ,
    \data[35] }));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[7]));
 sg13g2_buf_1 fanout14 (.A(net15),
    .X(net14));
 sg13g2_buf_1 fanout15 (.A(net16),
    .X(net15));
 sg13g2_buf_1 fanout16 (.A(net23),
    .X(net16));
 sg13g2_buf_1 fanout17 (.A(net23),
    .X(net17));
 sg13g2_buf_1 fanout18 (.A(net23),
    .X(net18));
 sg13g2_buf_1 fanout19 (.A(net23),
    .X(net19));
 sg13g2_buf_1 fanout20 (.A(net23),
    .X(net20));
 sg13g2_buf_1 fanout21 (.A(net22),
    .X(net21));
 sg13g2_buf_1 fanout22 (.A(net23),
    .X(net22));
 sg13g2_buf_1 fanout23 (.A(_113_),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(net25),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(net28),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(net27),
    .X(net26));
 sg13g2_buf_1 fanout27 (.A(net28),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(_113_),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(_112_),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(net31),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net41),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(net41),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(net41),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net36),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(net40),
    .X(net36));
 sg13g2_buf_1 fanout37 (.A(net39),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(net39),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(net40),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net1),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net46),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(net46),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net46),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net1),
    .X(net46));
 sg13g2_tielo heichips25_internal (.L_LO(net));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(delaynet_0_clk));
 sg13g2_buf_16 clkbuf_1_0__f_clk (.X(clknet_1_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_1_1__f_clk (.X(clknet_1_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_0_clk_regs (.X(clknet_0_clk_regs),
    .A(clk_regs));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clk_regs));
 sg13g2_buf_16 delaybuf_0_clk (.X(delaynet_0_clk),
    .A(clk));
 sg13g2_antennanp ANTENNA_1 (.A(\adc_data[7] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_4 FILLER_0_266 ();
 sg13g2_fill_1 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_fill_1 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_4 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_4 FILLER_0_351 ();
 sg13g2_fill_1 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_fill_2 FILLER_0_387 ();
 sg13g2_fill_1 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_4 FILLER_0_407 ();
 sg13g2_fill_1 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_439 ();
 sg13g2_decap_8 FILLER_0_446 ();
 sg13g2_fill_1 FILLER_0_480 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_fill_2 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_215 ();
 sg13g2_decap_8 FILLER_1_222 ();
 sg13g2_decap_8 FILLER_1_229 ();
 sg13g2_decap_8 FILLER_1_236 ();
 sg13g2_decap_8 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_decap_4 FILLER_1_267 ();
 sg13g2_fill_2 FILLER_1_271 ();
 sg13g2_fill_2 FILLER_1_300 ();
 sg13g2_fill_1 FILLER_1_356 ();
 sg13g2_fill_2 FILLER_1_384 ();
 sg13g2_decap_4 FILLER_1_413 ();
 sg13g2_fill_2 FILLER_1_417 ();
 sg13g2_decap_8 FILLER_1_456 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_fill_1 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_fill_2 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_4 FILLER_2_200 ();
 sg13g2_fill_1 FILLER_2_204 ();
 sg13g2_decap_4 FILLER_2_232 ();
 sg13g2_fill_2 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_4 FILLER_2_279 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_4 FILLER_2_301 ();
 sg13g2_fill_1 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_316 ();
 sg13g2_decap_4 FILLER_2_323 ();
 sg13g2_fill_2 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_fill_2 FILLER_2_340 ();
 sg13g2_fill_1 FILLER_2_342 ();
 sg13g2_decap_4 FILLER_2_370 ();
 sg13g2_fill_1 FILLER_2_374 ();
 sg13g2_decap_4 FILLER_2_402 ();
 sg13g2_fill_1 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_fill_1 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_fill_2 FILLER_2_487 ();
 sg13g2_fill_1 FILLER_2_489 ();
 sg13g2_decap_8 FILLER_2_500 ();
 sg13g2_decap_8 FILLER_2_507 ();
 sg13g2_decap_8 FILLER_2_514 ();
 sg13g2_decap_8 FILLER_2_521 ();
 sg13g2_decap_8 FILLER_2_528 ();
 sg13g2_decap_8 FILLER_2_535 ();
 sg13g2_decap_8 FILLER_2_542 ();
 sg13g2_decap_8 FILLER_2_549 ();
 sg13g2_decap_8 FILLER_2_556 ();
 sg13g2_decap_8 FILLER_2_563 ();
 sg13g2_decap_8 FILLER_2_570 ();
 sg13g2_decap_8 FILLER_2_577 ();
 sg13g2_decap_8 FILLER_2_584 ();
 sg13g2_decap_8 FILLER_2_591 ();
 sg13g2_decap_8 FILLER_2_598 ();
 sg13g2_decap_8 FILLER_2_605 ();
 sg13g2_decap_8 FILLER_2_612 ();
 sg13g2_decap_8 FILLER_2_619 ();
 sg13g2_decap_8 FILLER_2_626 ();
 sg13g2_decap_8 FILLER_2_633 ();
 sg13g2_decap_8 FILLER_2_640 ();
 sg13g2_decap_8 FILLER_2_647 ();
 sg13g2_decap_8 FILLER_2_654 ();
 sg13g2_decap_8 FILLER_2_661 ();
 sg13g2_decap_8 FILLER_2_668 ();
 sg13g2_decap_8 FILLER_2_675 ();
 sg13g2_decap_8 FILLER_2_682 ();
 sg13g2_decap_8 FILLER_2_689 ();
 sg13g2_decap_8 FILLER_2_696 ();
 sg13g2_decap_8 FILLER_2_703 ();
 sg13g2_decap_8 FILLER_2_710 ();
 sg13g2_decap_8 FILLER_2_717 ();
 sg13g2_decap_8 FILLER_2_724 ();
 sg13g2_decap_8 FILLER_2_731 ();
 sg13g2_decap_8 FILLER_2_738 ();
 sg13g2_decap_8 FILLER_2_745 ();
 sg13g2_decap_8 FILLER_2_752 ();
 sg13g2_decap_8 FILLER_2_759 ();
 sg13g2_decap_8 FILLER_2_766 ();
 sg13g2_decap_8 FILLER_2_773 ();
 sg13g2_decap_8 FILLER_2_780 ();
 sg13g2_decap_8 FILLER_2_787 ();
 sg13g2_decap_8 FILLER_2_794 ();
 sg13g2_decap_8 FILLER_2_801 ();
 sg13g2_decap_8 FILLER_2_808 ();
 sg13g2_decap_8 FILLER_2_815 ();
 sg13g2_decap_8 FILLER_2_822 ();
 sg13g2_decap_4 FILLER_2_829 ();
 sg13g2_fill_2 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_4 FILLER_3_207 ();
 sg13g2_fill_2 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_223 ();
 sg13g2_decap_4 FILLER_3_230 ();
 sg13g2_fill_2 FILLER_3_234 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_4 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_4 FILLER_3_336 ();
 sg13g2_fill_1 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_4 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_fill_1 FILLER_3_404 ();
 sg13g2_decap_8 FILLER_3_442 ();
 sg13g2_decap_4 FILLER_3_486 ();
 sg13g2_fill_2 FILLER_3_490 ();
 sg13g2_fill_2 FILLER_3_502 ();
 sg13g2_decap_4 FILLER_3_514 ();
 sg13g2_decap_8 FILLER_3_528 ();
 sg13g2_decap_8 FILLER_3_535 ();
 sg13g2_decap_8 FILLER_3_569 ();
 sg13g2_decap_8 FILLER_3_576 ();
 sg13g2_decap_8 FILLER_3_583 ();
 sg13g2_decap_8 FILLER_3_590 ();
 sg13g2_decap_8 FILLER_3_597 ();
 sg13g2_decap_8 FILLER_3_604 ();
 sg13g2_decap_8 FILLER_3_611 ();
 sg13g2_decap_8 FILLER_3_618 ();
 sg13g2_decap_8 FILLER_3_625 ();
 sg13g2_decap_8 FILLER_3_632 ();
 sg13g2_decap_8 FILLER_3_639 ();
 sg13g2_decap_8 FILLER_3_646 ();
 sg13g2_decap_8 FILLER_3_653 ();
 sg13g2_decap_8 FILLER_3_660 ();
 sg13g2_decap_8 FILLER_3_667 ();
 sg13g2_decap_8 FILLER_3_674 ();
 sg13g2_decap_8 FILLER_3_681 ();
 sg13g2_decap_8 FILLER_3_688 ();
 sg13g2_decap_8 FILLER_3_695 ();
 sg13g2_decap_8 FILLER_3_702 ();
 sg13g2_decap_8 FILLER_3_709 ();
 sg13g2_decap_8 FILLER_3_716 ();
 sg13g2_decap_8 FILLER_3_723 ();
 sg13g2_decap_8 FILLER_3_730 ();
 sg13g2_decap_8 FILLER_3_737 ();
 sg13g2_decap_8 FILLER_3_744 ();
 sg13g2_decap_8 FILLER_3_751 ();
 sg13g2_decap_8 FILLER_3_758 ();
 sg13g2_decap_8 FILLER_3_765 ();
 sg13g2_decap_8 FILLER_3_772 ();
 sg13g2_decap_8 FILLER_3_779 ();
 sg13g2_decap_8 FILLER_3_786 ();
 sg13g2_decap_8 FILLER_3_793 ();
 sg13g2_decap_8 FILLER_3_800 ();
 sg13g2_decap_8 FILLER_3_807 ();
 sg13g2_decap_8 FILLER_3_814 ();
 sg13g2_decap_8 FILLER_3_821 ();
 sg13g2_decap_8 FILLER_3_828 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_4 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_fill_2 FILLER_4_249 ();
 sg13g2_fill_1 FILLER_4_322 ();
 sg13g2_fill_2 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_4 FILLER_4_350 ();
 sg13g2_decap_4 FILLER_4_359 ();
 sg13g2_fill_1 FILLER_4_363 ();
 sg13g2_fill_2 FILLER_4_373 ();
 sg13g2_fill_1 FILLER_4_375 ();
 sg13g2_fill_2 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_fill_2 FILLER_4_395 ();
 sg13g2_fill_1 FILLER_4_397 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_1 FILLER_4_428 ();
 sg13g2_decap_4 FILLER_4_466 ();
 sg13g2_fill_2 FILLER_4_470 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_fill_2 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_fill_1 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_220 ();
 sg13g2_decap_4 FILLER_5_241 ();
 sg13g2_fill_2 FILLER_5_245 ();
 sg13g2_decap_4 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_269 ();
 sg13g2_decap_8 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_4 FILLER_5_318 ();
 sg13g2_fill_1 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_4 FILLER_5_379 ();
 sg13g2_fill_2 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_fill_2 FILLER_5_398 ();
 sg13g2_fill_1 FILLER_5_400 ();
 sg13g2_decap_8 FILLER_5_425 ();
 sg13g2_fill_1 FILLER_5_432 ();
 sg13g2_fill_2 FILLER_5_437 ();
 sg13g2_decap_4 FILLER_5_468 ();
 sg13g2_fill_1 FILLER_5_472 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_fill_2 FILLER_5_504 ();
 sg13g2_fill_1 FILLER_5_506 ();
 sg13g2_decap_8 FILLER_5_516 ();
 sg13g2_decap_8 FILLER_5_523 ();
 sg13g2_decap_4 FILLER_5_530 ();
 sg13g2_fill_2 FILLER_5_534 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_fill_2 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_fill_2 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_decap_8 FILLER_6_765 ();
 sg13g2_decap_8 FILLER_6_772 ();
 sg13g2_decap_8 FILLER_6_779 ();
 sg13g2_decap_8 FILLER_6_786 ();
 sg13g2_decap_8 FILLER_6_793 ();
 sg13g2_decap_8 FILLER_6_800 ();
 sg13g2_decap_8 FILLER_6_807 ();
 sg13g2_decap_8 FILLER_6_814 ();
 sg13g2_decap_8 FILLER_6_821 ();
 sg13g2_decap_8 FILLER_6_828 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_765 ();
 sg13g2_decap_8 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_779 ();
 sg13g2_decap_8 FILLER_7_786 ();
 sg13g2_decap_8 FILLER_7_793 ();
 sg13g2_decap_8 FILLER_7_800 ();
 sg13g2_fill_2 FILLER_7_807 ();
 sg13g2_fill_1 FILLER_7_809 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_4 FILLER_8_32 ();
 sg13g2_fill_2 FILLER_8_36 ();
 sg13g2_decap_8 FILLER_8_48 ();
 sg13g2_fill_1 FILLER_8_55 ();
 sg13g2_decap_8 FILLER_8_765 ();
 sg13g2_decap_8 FILLER_8_772 ();
 sg13g2_decap_8 FILLER_8_779 ();
 sg13g2_decap_8 FILLER_8_786 ();
 sg13g2_decap_8 FILLER_8_793 ();
 sg13g2_decap_8 FILLER_8_800 ();
 sg13g2_decap_8 FILLER_8_807 ();
 sg13g2_decap_8 FILLER_8_814 ();
 sg13g2_decap_8 FILLER_8_821 ();
 sg13g2_decap_8 FILLER_8_828 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_4 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_765 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_8 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_786 ();
 sg13g2_decap_8 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_55 ();
 sg13g2_decap_8 FILLER_10_765 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_4 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_765 ();
 sg13g2_decap_8 FILLER_11_772 ();
 sg13g2_decap_8 FILLER_11_779 ();
 sg13g2_decap_8 FILLER_11_786 ();
 sg13g2_decap_8 FILLER_11_793 ();
 sg13g2_decap_8 FILLER_11_800 ();
 sg13g2_decap_8 FILLER_11_807 ();
 sg13g2_decap_8 FILLER_11_814 ();
 sg13g2_decap_8 FILLER_11_821 ();
 sg13g2_decap_8 FILLER_11_828 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_4 FILLER_12_11 ();
 sg13g2_fill_2 FILLER_12_15 ();
 sg13g2_decap_8 FILLER_12_27 ();
 sg13g2_decap_8 FILLER_12_44 ();
 sg13g2_decap_4 FILLER_12_51 ();
 sg13g2_fill_1 FILLER_12_55 ();
 sg13g2_decap_8 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_772 ();
 sg13g2_decap_8 FILLER_12_779 ();
 sg13g2_decap_8 FILLER_12_786 ();
 sg13g2_decap_8 FILLER_12_793 ();
 sg13g2_decap_8 FILLER_12_800 ();
 sg13g2_decap_8 FILLER_12_807 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_8 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_828 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_fill_1 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_fill_2 FILLER_13_53 ();
 sg13g2_fill_1 FILLER_13_55 ();
 sg13g2_decap_8 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_772 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_decap_8 FILLER_13_786 ();
 sg13g2_decap_8 FILLER_13_793 ();
 sg13g2_decap_8 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_4 FILLER_15_25 ();
 sg13g2_fill_1 FILLER_15_29 ();
 sg13g2_decap_8 FILLER_15_40 ();
 sg13g2_decap_8 FILLER_15_47 ();
 sg13g2_fill_2 FILLER_15_54 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_8 FILLER_15_772 ();
 sg13g2_decap_8 FILLER_15_779 ();
 sg13g2_decap_8 FILLER_15_786 ();
 sg13g2_decap_8 FILLER_15_793 ();
 sg13g2_decap_8 FILLER_15_800 ();
 sg13g2_decap_8 FILLER_15_807 ();
 sg13g2_decap_8 FILLER_15_814 ();
 sg13g2_decap_8 FILLER_15_821 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_6 ();
 sg13g2_decap_8 FILLER_17_17 ();
 sg13g2_decap_4 FILLER_17_24 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_40 ();
 sg13g2_decap_8 FILLER_17_47 ();
 sg13g2_fill_2 FILLER_17_54 ();
 sg13g2_decap_8 FILLER_17_765 ();
 sg13g2_decap_8 FILLER_17_772 ();
 sg13g2_decap_8 FILLER_17_779 ();
 sg13g2_decap_8 FILLER_17_786 ();
 sg13g2_decap_8 FILLER_17_793 ();
 sg13g2_decap_8 FILLER_17_800 ();
 sg13g2_decap_8 FILLER_17_807 ();
 sg13g2_decap_8 FILLER_17_814 ();
 sg13g2_decap_8 FILLER_17_821 ();
 sg13g2_decap_8 FILLER_17_828 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_fill_1 FILLER_19_8 ();
 sg13g2_decap_8 FILLER_19_19 ();
 sg13g2_decap_8 FILLER_19_26 ();
 sg13g2_decap_4 FILLER_19_33 ();
 sg13g2_decap_8 FILLER_19_47 ();
 sg13g2_fill_2 FILLER_19_54 ();
 sg13g2_decap_8 FILLER_19_765 ();
 sg13g2_decap_8 FILLER_19_772 ();
 sg13g2_decap_8 FILLER_19_779 ();
 sg13g2_decap_8 FILLER_19_786 ();
 sg13g2_decap_8 FILLER_19_793 ();
 sg13g2_decap_8 FILLER_19_800 ();
 sg13g2_decap_8 FILLER_19_807 ();
 sg13g2_decap_8 FILLER_19_814 ();
 sg13g2_decap_8 FILLER_19_821 ();
 sg13g2_decap_8 FILLER_19_828 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_765 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_779 ();
 sg13g2_decap_8 FILLER_20_786 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_8 FILLER_20_817 ();
 sg13g2_decap_8 FILLER_20_824 ();
 sg13g2_decap_4 FILLER_20_831 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_4 FILLER_21_11 ();
 sg13g2_fill_1 FILLER_21_15 ();
 sg13g2_fill_1 FILLER_21_26 ();
 sg13g2_decap_8 FILLER_21_31 ();
 sg13g2_decap_8 FILLER_21_38 ();
 sg13g2_decap_8 FILLER_21_45 ();
 sg13g2_decap_4 FILLER_21_52 ();
 sg13g2_decap_8 FILLER_21_765 ();
 sg13g2_decap_8 FILLER_21_772 ();
 sg13g2_decap_8 FILLER_21_779 ();
 sg13g2_decap_8 FILLER_21_786 ();
 sg13g2_decap_8 FILLER_21_793 ();
 sg13g2_decap_8 FILLER_21_800 ();
 sg13g2_fill_1 FILLER_21_807 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_4 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_15 ();
 sg13g2_decap_8 FILLER_22_48 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_decap_8 FILLER_22_779 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_793 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_4 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_765 ();
 sg13g2_decap_8 FILLER_23_772 ();
 sg13g2_decap_8 FILLER_23_779 ();
 sg13g2_decap_8 FILLER_23_786 ();
 sg13g2_decap_8 FILLER_23_793 ();
 sg13g2_decap_8 FILLER_23_800 ();
 sg13g2_decap_8 FILLER_23_807 ();
 sg13g2_decap_8 FILLER_23_814 ();
 sg13g2_decap_8 FILLER_23_821 ();
 sg13g2_decap_8 FILLER_23_828 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_4 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_22 ();
 sg13g2_decap_8 FILLER_24_41 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_786 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_4 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_8 FILLER_25_856 ();
 sg13g2_decap_8 FILLER_25_863 ();
 sg13g2_decap_8 FILLER_25_870 ();
 sg13g2_decap_8 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_25_884 ();
 sg13g2_decap_8 FILLER_25_891 ();
 sg13g2_decap_8 FILLER_25_898 ();
 sg13g2_decap_8 FILLER_25_905 ();
 sg13g2_decap_8 FILLER_25_912 ();
 sg13g2_decap_8 FILLER_25_919 ();
 sg13g2_decap_8 FILLER_25_926 ();
 sg13g2_decap_8 FILLER_25_933 ();
 sg13g2_decap_8 FILLER_25_940 ();
 sg13g2_decap_8 FILLER_25_947 ();
 sg13g2_decap_8 FILLER_25_954 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_968 ();
 sg13g2_decap_8 FILLER_25_975 ();
 sg13g2_decap_8 FILLER_25_982 ();
 sg13g2_decap_8 FILLER_25_989 ();
 sg13g2_decap_4 FILLER_25_996 ();
 sg13g2_decap_4 FILLER_25_1025 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_4 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_22 ();
 sg13g2_decap_4 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_decap_8 FILLER_26_765 ();
 sg13g2_decap_8 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_779 ();
 sg13g2_decap_8 FILLER_26_786 ();
 sg13g2_decap_8 FILLER_26_793 ();
 sg13g2_decap_8 FILLER_26_800 ();
 sg13g2_decap_8 FILLER_26_807 ();
 sg13g2_decap_8 FILLER_26_814 ();
 sg13g2_decap_8 FILLER_26_821 ();
 sg13g2_decap_8 FILLER_26_828 ();
 sg13g2_fill_2 FILLER_26_835 ();
 sg13g2_fill_1 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_875 ();
 sg13g2_decap_8 FILLER_26_882 ();
 sg13g2_decap_8 FILLER_26_889 ();
 sg13g2_decap_8 FILLER_26_896 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_910 ();
 sg13g2_decap_8 FILLER_26_917 ();
 sg13g2_decap_8 FILLER_26_924 ();
 sg13g2_decap_8 FILLER_26_931 ();
 sg13g2_decap_8 FILLER_26_938 ();
 sg13g2_decap_8 FILLER_26_945 ();
 sg13g2_decap_8 FILLER_26_952 ();
 sg13g2_decap_8 FILLER_26_959 ();
 sg13g2_decap_8 FILLER_26_966 ();
 sg13g2_decap_8 FILLER_26_973 ();
 sg13g2_decap_8 FILLER_26_980 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_decap_8 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_1001 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_decap_8 FILLER_27_772 ();
 sg13g2_decap_8 FILLER_27_779 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_decap_8 FILLER_27_954 ();
 sg13g2_decap_8 FILLER_27_961 ();
 sg13g2_decap_8 FILLER_27_968 ();
 sg13g2_decap_8 FILLER_27_975 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_4 FILLER_27_1024 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_4 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_765 ();
 sg13g2_decap_8 FILLER_28_772 ();
 sg13g2_decap_8 FILLER_28_779 ();
 sg13g2_decap_8 FILLER_28_786 ();
 sg13g2_decap_8 FILLER_28_793 ();
 sg13g2_decap_8 FILLER_28_800 ();
 sg13g2_decap_8 FILLER_28_807 ();
 sg13g2_decap_8 FILLER_28_814 ();
 sg13g2_decap_8 FILLER_28_821 ();
 sg13g2_decap_8 FILLER_28_828 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_decap_8 FILLER_28_842 ();
 sg13g2_decap_8 FILLER_28_849 ();
 sg13g2_decap_4 FILLER_28_856 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_18 ();
 sg13g2_fill_2 FILLER_29_25 ();
 sg13g2_decap_8 FILLER_29_47 ();
 sg13g2_fill_2 FILLER_29_54 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_11 ();
 sg13g2_decap_8 FILLER_30_18 ();
 sg13g2_decap_4 FILLER_30_25 ();
 sg13g2_decap_8 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_772 ();
 sg13g2_decap_8 FILLER_30_779 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_18 ();
 sg13g2_decap_8 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_53 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_765 ();
 sg13g2_decap_8 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_779 ();
 sg13g2_decap_8 FILLER_31_786 ();
 sg13g2_decap_8 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_fill_1 FILLER_31_828 ();
 sg13g2_decap_4 FILLER_31_856 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_4 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_decap_8 FILLER_32_47 ();
 sg13g2_fill_2 FILLER_32_54 ();
 sg13g2_decap_8 FILLER_32_765 ();
 sg13g2_decap_8 FILLER_32_772 ();
 sg13g2_decap_8 FILLER_32_779 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_decap_8 FILLER_32_793 ();
 sg13g2_decap_8 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_814 ();
 sg13g2_decap_8 FILLER_32_821 ();
 sg13g2_fill_1 FILLER_32_828 ();
 sg13g2_decap_8 FILLER_32_849 ();
 sg13g2_decap_4 FILLER_32_856 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_765 ();
 sg13g2_decap_8 FILLER_33_772 ();
 sg13g2_decap_8 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_decap_8 FILLER_33_821 ();
 sg13g2_fill_1 FILLER_33_828 ();
 sg13g2_decap_4 FILLER_33_856 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_765 ();
 sg13g2_decap_8 FILLER_34_772 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_8 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_793 ();
 sg13g2_decap_8 FILLER_34_800 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_decap_8 FILLER_34_814 ();
 sg13g2_decap_4 FILLER_34_821 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_772 ();
 sg13g2_decap_8 FILLER_35_779 ();
 sg13g2_decap_8 FILLER_35_786 ();
 sg13g2_decap_8 FILLER_35_793 ();
 sg13g2_decap_8 FILLER_35_800 ();
 sg13g2_decap_8 FILLER_35_807 ();
 sg13g2_decap_8 FILLER_35_814 ();
 sg13g2_decap_4 FILLER_35_821 ();
 sg13g2_fill_2 FILLER_35_825 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_4 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_4 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_790 ();
 sg13g2_decap_8 FILLER_36_797 ();
 sg13g2_decap_8 FILLER_36_804 ();
 sg13g2_decap_8 FILLER_36_811 ();
 sg13g2_decap_8 FILLER_36_818 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_765 ();
 sg13g2_decap_8 FILLER_37_772 ();
 sg13g2_decap_8 FILLER_37_779 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_807 ();
 sg13g2_decap_4 FILLER_37_814 ();
 sg13g2_fill_2 FILLER_37_818 ();
 sg13g2_decap_4 FILLER_37_830 ();
 sg13g2_fill_1 FILLER_37_834 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_765 ();
 sg13g2_decap_8 FILLER_38_772 ();
 sg13g2_decap_8 FILLER_38_779 ();
 sg13g2_decap_8 FILLER_38_786 ();
 sg13g2_decap_8 FILLER_38_793 ();
 sg13g2_decap_8 FILLER_38_800 ();
 sg13g2_decap_8 FILLER_38_807 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_4 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_fill_2 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_47 ();
 sg13g2_fill_2 FILLER_39_54 ();
 sg13g2_decap_8 FILLER_39_765 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_4 FILLER_39_814 ();
 sg13g2_fill_2 FILLER_39_859 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_fill_1 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_765 ();
 sg13g2_decap_8 FILLER_40_772 ();
 sg13g2_decap_8 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_fill_2 FILLER_40_832 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_4 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_765 ();
 sg13g2_decap_8 FILLER_41_772 ();
 sg13g2_decap_8 FILLER_41_779 ();
 sg13g2_decap_8 FILLER_41_786 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_828 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_53 ();
 sg13g2_fill_1 FILLER_42_55 ();
 sg13g2_decap_8 FILLER_42_765 ();
 sg13g2_decap_8 FILLER_42_772 ();
 sg13g2_decap_8 FILLER_42_779 ();
 sg13g2_decap_8 FILLER_42_786 ();
 sg13g2_decap_8 FILLER_42_793 ();
 sg13g2_decap_8 FILLER_42_800 ();
 sg13g2_decap_8 FILLER_42_807 ();
 sg13g2_decap_8 FILLER_42_814 ();
 sg13g2_decap_8 FILLER_42_821 ();
 sg13g2_decap_4 FILLER_42_842 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_decap_4 FILLER_42_857 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_765 ();
 sg13g2_decap_8 FILLER_43_772 ();
 sg13g2_decap_8 FILLER_43_779 ();
 sg13g2_decap_8 FILLER_43_786 ();
 sg13g2_decap_8 FILLER_43_793 ();
 sg13g2_decap_8 FILLER_43_800 ();
 sg13g2_decap_8 FILLER_43_807 ();
 sg13g2_decap_8 FILLER_43_814 ();
 sg13g2_decap_8 FILLER_43_821 ();
 sg13g2_decap_8 FILLER_43_828 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_78 ();
 sg13g2_decap_8 FILLER_44_85 ();
 sg13g2_decap_4 FILLER_44_92 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_167 ();
 sg13g2_fill_2 FILLER_44_209 ();
 sg13g2_decap_8 FILLER_44_227 ();
 sg13g2_decap_4 FILLER_44_261 ();
 sg13g2_fill_2 FILLER_44_265 ();
 sg13g2_fill_2 FILLER_44_368 ();
 sg13g2_decap_4 FILLER_44_393 ();
 sg13g2_fill_2 FILLER_44_424 ();
 sg13g2_decap_4 FILLER_44_526 ();
 sg13g2_decap_8 FILLER_44_570 ();
 sg13g2_decap_8 FILLER_44_577 ();
 sg13g2_decap_8 FILLER_44_584 ();
 sg13g2_decap_8 FILLER_44_591 ();
 sg13g2_decap_8 FILLER_44_598 ();
 sg13g2_decap_8 FILLER_44_605 ();
 sg13g2_decap_8 FILLER_44_612 ();
 sg13g2_decap_8 FILLER_44_619 ();
 sg13g2_decap_8 FILLER_44_626 ();
 sg13g2_decap_4 FILLER_44_671 ();
 sg13g2_decap_8 FILLER_44_688 ();
 sg13g2_decap_8 FILLER_44_695 ();
 sg13g2_decap_8 FILLER_44_741 ();
 sg13g2_decap_8 FILLER_44_748 ();
 sg13g2_decap_8 FILLER_44_755 ();
 sg13g2_decap_8 FILLER_44_762 ();
 sg13g2_decap_8 FILLER_44_769 ();
 sg13g2_decap_8 FILLER_44_776 ();
 sg13g2_decap_8 FILLER_44_783 ();
 sg13g2_decap_8 FILLER_44_790 ();
 sg13g2_decap_8 FILLER_44_797 ();
 sg13g2_decap_8 FILLER_44_804 ();
 sg13g2_decap_8 FILLER_44_811 ();
 sg13g2_decap_8 FILLER_44_818 ();
 sg13g2_decap_8 FILLER_44_825 ();
 sg13g2_decap_8 FILLER_44_832 ();
 sg13g2_decap_8 FILLER_44_839 ();
 sg13g2_decap_8 FILLER_44_846 ();
 sg13g2_decap_8 FILLER_44_853 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_4 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_106 ();
 sg13g2_decap_8 FILLER_45_113 ();
 sg13g2_decap_8 FILLER_45_120 ();
 sg13g2_fill_1 FILLER_45_127 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_decap_8 FILLER_45_236 ();
 sg13g2_decap_8 FILLER_45_243 ();
 sg13g2_fill_2 FILLER_45_250 ();
 sg13g2_decap_8 FILLER_45_292 ();
 sg13g2_decap_8 FILLER_45_299 ();
 sg13g2_decap_8 FILLER_45_333 ();
 sg13g2_fill_1 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_450 ();
 sg13g2_decap_8 FILLER_45_563 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_decap_8 FILLER_45_577 ();
 sg13g2_decap_8 FILLER_45_584 ();
 sg13g2_decap_8 FILLER_45_591 ();
 sg13g2_decap_8 FILLER_45_598 ();
 sg13g2_decap_8 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_decap_8 FILLER_45_619 ();
 sg13g2_decap_8 FILLER_45_626 ();
 sg13g2_decap_8 FILLER_45_633 ();
 sg13g2_decap_8 FILLER_45_640 ();
 sg13g2_decap_8 FILLER_45_647 ();
 sg13g2_fill_2 FILLER_45_654 ();
 sg13g2_fill_1 FILLER_45_656 ();
 sg13g2_decap_8 FILLER_45_670 ();
 sg13g2_decap_8 FILLER_45_677 ();
 sg13g2_decap_8 FILLER_45_684 ();
 sg13g2_decap_8 FILLER_45_691 ();
 sg13g2_decap_8 FILLER_45_698 ();
 sg13g2_decap_8 FILLER_45_705 ();
 sg13g2_decap_8 FILLER_45_712 ();
 sg13g2_decap_4 FILLER_45_719 ();
 sg13g2_fill_1 FILLER_45_723 ();
 sg13g2_decap_8 FILLER_45_727 ();
 sg13g2_decap_8 FILLER_45_734 ();
 sg13g2_decap_8 FILLER_45_741 ();
 sg13g2_decap_8 FILLER_45_748 ();
 sg13g2_decap_8 FILLER_45_755 ();
 sg13g2_decap_8 FILLER_45_762 ();
 sg13g2_decap_8 FILLER_45_769 ();
 sg13g2_decap_8 FILLER_45_776 ();
 sg13g2_decap_8 FILLER_45_783 ();
 sg13g2_decap_8 FILLER_45_790 ();
 sg13g2_decap_8 FILLER_45_797 ();
 sg13g2_decap_8 FILLER_45_804 ();
 sg13g2_decap_8 FILLER_45_811 ();
 sg13g2_decap_8 FILLER_45_818 ();
 sg13g2_decap_8 FILLER_45_825 ();
 sg13g2_decap_8 FILLER_45_832 ();
 sg13g2_decap_8 FILLER_45_839 ();
 sg13g2_decap_8 FILLER_45_846 ();
 sg13g2_decap_8 FILLER_45_853 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_4 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_142 ();
 sg13g2_decap_8 FILLER_46_149 ();
 sg13g2_decap_4 FILLER_46_156 ();
 sg13g2_fill_1 FILLER_46_160 ();
 sg13g2_decap_8 FILLER_46_171 ();
 sg13g2_decap_8 FILLER_46_178 ();
 sg13g2_fill_2 FILLER_46_195 ();
 sg13g2_fill_2 FILLER_46_234 ();
 sg13g2_fill_2 FILLER_46_263 ();
 sg13g2_fill_2 FILLER_46_278 ();
 sg13g2_decap_8 FILLER_46_285 ();
 sg13g2_decap_8 FILLER_46_292 ();
 sg13g2_decap_8 FILLER_46_299 ();
 sg13g2_decap_8 FILLER_46_306 ();
 sg13g2_decap_8 FILLER_46_313 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_418 ();
 sg13g2_decap_8 FILLER_46_429 ();
 sg13g2_decap_4 FILLER_46_436 ();
 sg13g2_fill_1 FILLER_46_440 ();
 sg13g2_fill_2 FILLER_46_455 ();
 sg13g2_decap_4 FILLER_46_461 ();
 sg13g2_fill_2 FILLER_46_465 ();
 sg13g2_decap_8 FILLER_46_477 ();
 sg13g2_decap_8 FILLER_46_484 ();
 sg13g2_decap_8 FILLER_46_491 ();
 sg13g2_decap_4 FILLER_46_498 ();
 sg13g2_decap_8 FILLER_46_512 ();
 sg13g2_fill_1 FILLER_46_519 ();
 sg13g2_decap_8 FILLER_46_540 ();
 sg13g2_decap_8 FILLER_46_547 ();
 sg13g2_decap_8 FILLER_46_554 ();
 sg13g2_decap_8 FILLER_46_561 ();
 sg13g2_decap_8 FILLER_46_568 ();
 sg13g2_decap_8 FILLER_46_575 ();
 sg13g2_decap_8 FILLER_46_582 ();
 sg13g2_decap_8 FILLER_46_589 ();
 sg13g2_decap_8 FILLER_46_596 ();
 sg13g2_decap_8 FILLER_46_603 ();
 sg13g2_decap_8 FILLER_46_610 ();
 sg13g2_decap_8 FILLER_46_617 ();
 sg13g2_decap_8 FILLER_46_624 ();
 sg13g2_decap_8 FILLER_46_631 ();
 sg13g2_decap_8 FILLER_46_638 ();
 sg13g2_decap_8 FILLER_46_645 ();
 sg13g2_decap_8 FILLER_46_652 ();
 sg13g2_decap_8 FILLER_46_659 ();
 sg13g2_decap_8 FILLER_46_666 ();
 sg13g2_decap_8 FILLER_46_673 ();
 sg13g2_decap_8 FILLER_46_680 ();
 sg13g2_decap_8 FILLER_46_687 ();
 sg13g2_decap_8 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_701 ();
 sg13g2_decap_8 FILLER_46_708 ();
 sg13g2_decap_8 FILLER_46_715 ();
 sg13g2_decap_8 FILLER_46_722 ();
 sg13g2_decap_8 FILLER_46_729 ();
 sg13g2_decap_8 FILLER_46_736 ();
 sg13g2_decap_8 FILLER_46_743 ();
 sg13g2_decap_8 FILLER_46_750 ();
 sg13g2_decap_8 FILLER_46_757 ();
 sg13g2_decap_8 FILLER_46_764 ();
 sg13g2_decap_8 FILLER_46_771 ();
 sg13g2_decap_8 FILLER_46_778 ();
 sg13g2_decap_8 FILLER_46_785 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_8 FILLER_46_799 ();
 sg13g2_decap_8 FILLER_46_806 ();
 sg13g2_decap_8 FILLER_46_813 ();
 sg13g2_decap_8 FILLER_46_820 ();
 sg13g2_decap_8 FILLER_46_827 ();
 sg13g2_decap_8 FILLER_46_834 ();
 sg13g2_decap_8 FILLER_46_841 ();
 sg13g2_decap_8 FILLER_46_848 ();
 sg13g2_decap_8 FILLER_46_855 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_4 FILLER_47_182 ();
 sg13g2_fill_2 FILLER_47_186 ();
 sg13g2_decap_4 FILLER_47_218 ();
 sg13g2_fill_1 FILLER_47_222 ();
 sg13g2_fill_1 FILLER_47_230 ();
 sg13g2_fill_2 FILLER_47_239 ();
 sg13g2_fill_1 FILLER_47_241 ();
 sg13g2_fill_2 FILLER_47_264 ();
 sg13g2_fill_1 FILLER_47_274 ();
 sg13g2_decap_8 FILLER_47_288 ();
 sg13g2_decap_8 FILLER_47_295 ();
 sg13g2_fill_1 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_fill_2 FILLER_47_403 ();
 sg13g2_decap_8 FILLER_47_415 ();
 sg13g2_decap_4 FILLER_47_422 ();
 sg13g2_decap_8 FILLER_47_453 ();
 sg13g2_decap_8 FILLER_47_460 ();
 sg13g2_decap_8 FILLER_47_467 ();
 sg13g2_decap_8 FILLER_47_474 ();
 sg13g2_decap_8 FILLER_47_481 ();
 sg13g2_decap_8 FILLER_47_488 ();
 sg13g2_decap_8 FILLER_47_495 ();
 sg13g2_decap_8 FILLER_47_502 ();
 sg13g2_decap_8 FILLER_47_509 ();
 sg13g2_decap_8 FILLER_47_516 ();
 sg13g2_decap_8 FILLER_47_523 ();
 sg13g2_decap_8 FILLER_47_530 ();
 sg13g2_decap_8 FILLER_47_537 ();
 sg13g2_decap_8 FILLER_47_544 ();
 sg13g2_decap_8 FILLER_47_551 ();
 sg13g2_decap_8 FILLER_47_558 ();
 sg13g2_decap_8 FILLER_47_565 ();
 sg13g2_decap_8 FILLER_47_572 ();
 sg13g2_decap_8 FILLER_47_579 ();
 sg13g2_decap_8 FILLER_47_586 ();
 sg13g2_decap_8 FILLER_47_593 ();
 sg13g2_decap_8 FILLER_47_600 ();
 sg13g2_decap_8 FILLER_47_607 ();
 sg13g2_decap_8 FILLER_47_614 ();
 sg13g2_decap_8 FILLER_47_621 ();
 sg13g2_decap_8 FILLER_47_628 ();
 sg13g2_decap_8 FILLER_47_635 ();
 sg13g2_decap_8 FILLER_47_642 ();
 sg13g2_decap_8 FILLER_47_649 ();
 sg13g2_decap_8 FILLER_47_656 ();
 sg13g2_decap_8 FILLER_47_663 ();
 sg13g2_decap_8 FILLER_47_670 ();
 sg13g2_decap_8 FILLER_47_677 ();
 sg13g2_decap_8 FILLER_47_684 ();
 sg13g2_decap_8 FILLER_47_691 ();
 sg13g2_decap_8 FILLER_47_698 ();
 sg13g2_decap_8 FILLER_47_705 ();
 sg13g2_decap_8 FILLER_47_712 ();
 sg13g2_decap_8 FILLER_47_719 ();
 sg13g2_decap_8 FILLER_47_726 ();
 sg13g2_decap_8 FILLER_47_733 ();
 sg13g2_decap_8 FILLER_47_740 ();
 sg13g2_decap_8 FILLER_47_747 ();
 sg13g2_decap_8 FILLER_47_754 ();
 sg13g2_decap_8 FILLER_47_761 ();
 sg13g2_decap_8 FILLER_47_768 ();
 sg13g2_decap_8 FILLER_47_775 ();
 sg13g2_decap_8 FILLER_47_782 ();
 sg13g2_decap_8 FILLER_47_789 ();
 sg13g2_decap_8 FILLER_47_796 ();
 sg13g2_decap_8 FILLER_47_803 ();
 sg13g2_decap_8 FILLER_47_810 ();
 sg13g2_decap_8 FILLER_47_817 ();
 sg13g2_decap_8 FILLER_47_824 ();
 sg13g2_decap_8 FILLER_47_831 ();
 sg13g2_decap_8 FILLER_47_838 ();
 sg13g2_decap_8 FILLER_47_845 ();
 sg13g2_decap_8 FILLER_47_852 ();
 sg13g2_fill_2 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_fill_1 FILLER_48_196 ();
 sg13g2_decap_4 FILLER_48_201 ();
 sg13g2_fill_1 FILLER_48_205 ();
 sg13g2_fill_1 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_335 ();
 sg13g2_decap_4 FILLER_48_367 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_436 ();
 sg13g2_decap_8 FILLER_48_443 ();
 sg13g2_decap_8 FILLER_48_450 ();
 sg13g2_decap_8 FILLER_48_457 ();
 sg13g2_decap_8 FILLER_48_464 ();
 sg13g2_decap_8 FILLER_48_471 ();
 sg13g2_decap_8 FILLER_48_478 ();
 sg13g2_decap_8 FILLER_48_485 ();
 sg13g2_decap_8 FILLER_48_492 ();
 sg13g2_decap_8 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_506 ();
 sg13g2_decap_8 FILLER_48_513 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_decap_8 FILLER_48_527 ();
 sg13g2_decap_8 FILLER_48_534 ();
 sg13g2_decap_8 FILLER_48_541 ();
 sg13g2_decap_8 FILLER_48_548 ();
 sg13g2_decap_8 FILLER_48_555 ();
 sg13g2_decap_8 FILLER_48_562 ();
 sg13g2_decap_8 FILLER_48_569 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_583 ();
 sg13g2_decap_8 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_597 ();
 sg13g2_decap_8 FILLER_48_604 ();
 sg13g2_decap_8 FILLER_48_611 ();
 sg13g2_decap_8 FILLER_48_618 ();
 sg13g2_decap_8 FILLER_48_625 ();
 sg13g2_decap_8 FILLER_48_632 ();
 sg13g2_decap_8 FILLER_48_639 ();
 sg13g2_decap_8 FILLER_48_646 ();
 sg13g2_decap_8 FILLER_48_653 ();
 sg13g2_decap_8 FILLER_48_660 ();
 sg13g2_decap_8 FILLER_48_667 ();
 sg13g2_decap_8 FILLER_48_674 ();
 sg13g2_decap_8 FILLER_48_681 ();
 sg13g2_decap_8 FILLER_48_688 ();
 sg13g2_decap_8 FILLER_48_695 ();
 sg13g2_decap_8 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_709 ();
 sg13g2_decap_8 FILLER_48_716 ();
 sg13g2_decap_8 FILLER_48_723 ();
 sg13g2_decap_8 FILLER_48_730 ();
 sg13g2_decap_8 FILLER_48_737 ();
 sg13g2_decap_8 FILLER_48_744 ();
 sg13g2_decap_8 FILLER_48_751 ();
 sg13g2_decap_8 FILLER_48_758 ();
 sg13g2_decap_8 FILLER_48_765 ();
 sg13g2_decap_8 FILLER_48_772 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_793 ();
 sg13g2_decap_8 FILLER_48_800 ();
 sg13g2_decap_8 FILLER_48_807 ();
 sg13g2_decap_8 FILLER_48_814 ();
 sg13g2_decap_8 FILLER_48_821 ();
 sg13g2_decap_8 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_835 ();
 sg13g2_decap_8 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_4 FILLER_48_856 ();
 sg13g2_fill_2 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_4 FILLER_49_214 ();
 sg13g2_fill_2 FILLER_49_218 ();
 sg13g2_fill_2 FILLER_49_225 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_232 ();
 sg13g2_fill_1 FILLER_49_239 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_4 FILLER_49_259 ();
 sg13g2_fill_1 FILLER_49_263 ();
 sg13g2_fill_2 FILLER_49_267 ();
 sg13g2_decap_4 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_285 ();
 sg13g2_fill_2 FILLER_49_292 ();
 sg13g2_fill_1 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_307 ();
 sg13g2_decap_8 FILLER_49_314 ();
 sg13g2_decap_8 FILLER_49_321 ();
 sg13g2_decap_8 FILLER_49_328 ();
 sg13g2_decap_4 FILLER_49_335 ();
 sg13g2_decap_8 FILLER_49_349 ();
 sg13g2_decap_8 FILLER_49_356 ();
 sg13g2_decap_8 FILLER_49_363 ();
 sg13g2_decap_8 FILLER_49_370 ();
 sg13g2_fill_2 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_390 ();
 sg13g2_decap_8 FILLER_49_397 ();
 sg13g2_decap_8 FILLER_49_404 ();
 sg13g2_decap_8 FILLER_49_411 ();
 sg13g2_decap_8 FILLER_49_418 ();
 sg13g2_decap_8 FILLER_49_425 ();
 sg13g2_decap_8 FILLER_49_432 ();
 sg13g2_decap_8 FILLER_49_439 ();
 sg13g2_decap_8 FILLER_49_446 ();
 sg13g2_decap_8 FILLER_49_453 ();
 sg13g2_decap_8 FILLER_49_460 ();
 sg13g2_decap_8 FILLER_49_467 ();
 sg13g2_decap_8 FILLER_49_474 ();
 sg13g2_decap_8 FILLER_49_481 ();
 sg13g2_decap_8 FILLER_49_488 ();
 sg13g2_decap_8 FILLER_49_495 ();
 sg13g2_decap_8 FILLER_49_502 ();
 sg13g2_decap_8 FILLER_49_509 ();
 sg13g2_decap_8 FILLER_49_516 ();
 sg13g2_decap_8 FILLER_49_523 ();
 sg13g2_decap_8 FILLER_49_530 ();
 sg13g2_decap_8 FILLER_49_537 ();
 sg13g2_decap_8 FILLER_49_544 ();
 sg13g2_decap_8 FILLER_49_551 ();
 sg13g2_decap_8 FILLER_49_558 ();
 sg13g2_decap_8 FILLER_49_565 ();
 sg13g2_decap_8 FILLER_49_572 ();
 sg13g2_decap_8 FILLER_49_579 ();
 sg13g2_decap_8 FILLER_49_586 ();
 sg13g2_decap_8 FILLER_49_593 ();
 sg13g2_decap_8 FILLER_49_600 ();
 sg13g2_decap_8 FILLER_49_607 ();
 sg13g2_decap_8 FILLER_49_614 ();
 sg13g2_decap_8 FILLER_49_621 ();
 sg13g2_decap_8 FILLER_49_628 ();
 sg13g2_decap_8 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_decap_8 FILLER_49_649 ();
 sg13g2_decap_8 FILLER_49_656 ();
 sg13g2_decap_8 FILLER_49_663 ();
 sg13g2_decap_8 FILLER_49_670 ();
 sg13g2_decap_8 FILLER_49_677 ();
 sg13g2_decap_8 FILLER_49_684 ();
 sg13g2_decap_8 FILLER_49_691 ();
 sg13g2_decap_8 FILLER_49_698 ();
 sg13g2_decap_8 FILLER_49_705 ();
 sg13g2_decap_8 FILLER_49_712 ();
 sg13g2_decap_8 FILLER_49_719 ();
 sg13g2_decap_8 FILLER_49_726 ();
 sg13g2_decap_8 FILLER_49_733 ();
 sg13g2_decap_8 FILLER_49_740 ();
 sg13g2_decap_8 FILLER_49_747 ();
 sg13g2_decap_8 FILLER_49_754 ();
 sg13g2_decap_8 FILLER_49_761 ();
 sg13g2_decap_8 FILLER_49_768 ();
 sg13g2_decap_8 FILLER_49_775 ();
 sg13g2_decap_8 FILLER_49_782 ();
 sg13g2_decap_8 FILLER_49_789 ();
 sg13g2_decap_8 FILLER_49_796 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_810 ();
 sg13g2_decap_8 FILLER_49_817 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_decap_8 FILLER_49_838 ();
 sg13g2_decap_8 FILLER_49_845 ();
 sg13g2_decap_8 FILLER_49_852 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 assign uio_oe[0] = net;
 assign uio_oe[1] = net47;
 assign uio_oe[2] = net48;
 assign uio_oe[3] = net49;
 assign uio_oe[4] = net50;
 assign uio_oe[5] = net51;
 assign uio_oe[6] = net52;
 assign uio_oe[7] = net53;
 assign uo_out[0] = net54;
 assign uo_out[1] = net55;
 assign uo_out[2] = net56;
 assign uo_out[3] = net57;
 assign uo_out[4] = net58;
 assign uo_out[5] = net59;
 assign uo_out[6] = net60;
 assign uo_out[7] = net61;
endmodule
