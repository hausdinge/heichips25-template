VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO delay_line
  CLASS BLOCK ;
  FOREIGN delay_line ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 60.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 15.380 0.000 17.580 60.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 16.280 60.000 18.480 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 46.280 60.000 48.480 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 21.580 0.000 23.780 60.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 22.480 60.000 24.680 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 59.600 34.280 60.000 ;
    END
  END clk
  PIN clk_delayed
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.900 0.400 44.300 ;
    END
  END clk_delayed
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2.200 0.000 2.600 0.400 ;
    END
  END reset
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 29.080 59.600 29.480 60.000 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.980 0.400 33.380 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.820 0.400 34.220 ;
    END
  END sel[2]
  PIN trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.600 36.340 60.000 36.740 ;
    END
  END trim[0]
  PIN trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.600 22.060 60.000 22.460 ;
    END
  END trim[1]
  PIN trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END trim[2]
  PIN trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.420 0.400 25.820 ;
    END
  END trim[3]
  PIN trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 39.640 59.600 40.040 60.000 ;
    END
  END trim[4]
  PIN trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.600 27.100 60.000 27.500 ;
    END
  END trim[5]
  PIN trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END trim[6]
  PIN trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.340 0.400 15.740 ;
    END
  END trim[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 57.120 53.070 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 57.120 53.140 ;
      LAYER Metal2 ;
        RECT 2.775 59.390 28.870 59.600 ;
        RECT 29.690 59.390 33.670 59.600 ;
        RECT 34.490 59.390 39.430 59.600 ;
        RECT 40.250 59.390 59.625 59.600 ;
        RECT 2.775 0.610 59.625 59.390 ;
        RECT 2.810 0.400 19.270 0.610 ;
        RECT 20.090 0.400 30.790 0.610 ;
        RECT 31.610 0.400 59.625 0.610 ;
      LAYER Metal3 ;
        RECT 0.400 44.510 59.665 56.380 ;
        RECT 0.610 43.690 59.665 44.510 ;
        RECT 0.400 36.950 59.665 43.690 ;
        RECT 0.400 36.130 59.390 36.950 ;
        RECT 0.400 34.430 59.665 36.130 ;
        RECT 0.610 33.610 59.665 34.430 ;
        RECT 0.400 33.590 59.665 33.610 ;
        RECT 0.610 32.770 59.665 33.590 ;
        RECT 0.400 27.710 59.665 32.770 ;
        RECT 0.400 26.890 59.390 27.710 ;
        RECT 0.400 26.030 59.665 26.890 ;
        RECT 0.610 25.210 59.665 26.030 ;
        RECT 0.400 22.670 59.665 25.210 ;
        RECT 0.400 21.850 59.390 22.670 ;
        RECT 0.400 15.950 59.665 21.850 ;
        RECT 0.610 15.130 59.665 15.950 ;
        RECT 0.400 1.160 59.665 15.130 ;
      LAYER Metal4 ;
        RECT 20.060 5.315 21.370 40.045 ;
        RECT 23.990 5.315 53.385 40.045 ;
      LAYER Metal5 ;
        RECT 25.775 21.320 53.425 21.520 ;
  END
END delay_line
END LIBRARY

